-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jul 24 2025 23:36:46

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__48096\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48094\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48083\ : std_logic;
signal \N__48076\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48058\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48047\ : std_logic;
signal \N__48040\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48038\ : std_logic;
signal \N__48031\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48022\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48012\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48002\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47984\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47940\ : std_logic;
signal \N__47939\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47936\ : std_logic;
signal \N__47933\ : std_logic;
signal \N__47932\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47926\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47909\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47900\ : std_logic;
signal \N__47899\ : std_logic;
signal \N__47896\ : std_logic;
signal \N__47893\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47845\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47790\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47710\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47646\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47585\ : std_logic;
signal \N__47574\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47571\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47558\ : std_logic;
signal \N__47551\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47535\ : std_logic;
signal \N__47532\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47521\ : std_logic;
signal \N__47518\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47506\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47491\ : std_logic;
signal \N__47488\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47471\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47459\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47441\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47438\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47435\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47420\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47417\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47389\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47386\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47338\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47318\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46989\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46984\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46941\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46894\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46865\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46521\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46511\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46489\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46472\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46437\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46368\ : std_logic;
signal \N__46365\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46357\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46337\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46330\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46260\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46147\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46127\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45969\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45922\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45910\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45846\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45776\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45770\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45738\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45720\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45710\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45675\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45566\ : std_logic;
signal \N__45565\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45521\ : std_logic;
signal \N__45518\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45420\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45413\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45379\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45360\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45331\ : std_logic;
signal \N__45322\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45308\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45275\ : std_logic;
signal \N__45272\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45258\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45204\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45192\ : std_logic;
signal \N__45189\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45179\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45171\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44891\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44881\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44876\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44814\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44797\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44767\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44729\ : std_logic;
signal \N__44726\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44690\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44681\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44608\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44598\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44511\ : std_logic;
signal \N__44508\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44501\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44484\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44447\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44412\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44391\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44384\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44284\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44211\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44064\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43996\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43942\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43925\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43918\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43877\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43867\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43785\ : std_logic;
signal \N__43782\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43689\ : std_logic;
signal \N__43686\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43624\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43541\ : std_logic;
signal \N__43540\ : std_logic;
signal \N__43537\ : std_logic;
signal \N__43534\ : std_logic;
signal \N__43531\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43444\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43422\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43374\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43343\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43301\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43234\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43207\ : std_logic;
signal \N__43204\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43188\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43083\ : std_logic;
signal \N__43080\ : std_logic;
signal \N__43077\ : std_logic;
signal \N__43074\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43026\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43015\ : std_logic;
signal \N__43012\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__43002\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42946\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42922\ : std_logic;
signal \N__42919\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42854\ : std_logic;
signal \N__42851\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42679\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42673\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42662\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42497\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42493\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42273\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42243\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42207\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42178\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42130\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42101\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42059\ : std_logic;
signal \N__42056\ : std_logic;
signal \N__42055\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42008\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41870\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41849\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41839\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41762\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41725\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41553\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41460\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41450\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41404\ : std_logic;
signal \N__41401\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41236\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41149\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41111\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40890\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40823\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40799\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40777\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40662\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40395\ : std_logic;
signal \N__40392\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40295\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40289\ : std_logic;
signal \N__40286\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40137\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40074\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40047\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40042\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39868\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39784\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39734\ : std_logic;
signal \N__39731\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39672\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39644\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39438\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39312\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38818\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38798\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38695\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38234\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38142\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38063\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37684\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37321\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36436\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \current_shift_inst.PI_CTRL.m7_2_cascade_\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_7\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_15\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_16\ : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_5 : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal \N_22_i_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.m14_2\ : std_logic;
signal pwm_duty_input_10 : std_logic;
signal pwm_duty_input_4 : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \current_shift_inst.PI_CTRL.N_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_13_cascade_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_23\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_178\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal un7_start_stop_0_a3 : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\ : std_logic;
signal \bfn_3_8_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_7\ : std_logic;
signal \bfn_3_9_0_\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_8\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_0\ : std_logic;
signal \bfn_3_11_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_8\ : std_logic;
signal \bfn_3_12_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_3_13_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \bfn_4_5_0_\ : std_logic;
signal un5_counter_cry_1 : std_logic;
signal un5_counter_cry_2 : std_logic;
signal un5_counter_cry_3 : std_logic;
signal un5_counter_cry_4 : std_logic;
signal un5_counter_cry_5 : std_logic;
signal un5_counter_cry_6 : std_logic;
signal un5_counter_cry_7 : std_logic;
signal un5_counter_cry_8 : std_logic;
signal \bfn_4_6_0_\ : std_logic;
signal un5_counter_cry_9 : std_logic;
signal un5_counter_cry_10 : std_logic;
signal un5_counter_cry_11 : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\ : std_logic;
signal pwm_duty_input_6 : std_logic;
signal i8_mux : std_logic;
signal \N_28_mux\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \bfn_4_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \counter_RNO_0Z0Z_7\ : std_logic;
signal \counterZ0Z_7\ : std_logic;
signal \counterZ0Z_2\ : std_logic;
signal \counterZ0Z_1\ : std_logic;
signal \un2_counter_5_cascade_\ : std_logic;
signal \counterZ0Z_8\ : std_logic;
signal \counterZ0Z_11\ : std_logic;
signal \counterZ0Z_9\ : std_logic;
signal \counterZ0Z_5\ : std_logic;
signal \counterZ0Z_4\ : std_logic;
signal \counterZ0Z_6\ : std_logic;
signal \counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_6\ : std_logic;
signal \counter_RNO_0Z0Z_12\ : std_logic;
signal \counterZ0Z_12\ : std_logic;
signal \counter_RNO_0Z0Z_10\ : std_logic;
signal \counterZ0Z_10\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_0\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal \counterZ0Z_0\ : std_logic;
signal \clk_10khz_RNIIENAZ0Z2_cascade_\ : std_logic;
signal \clk_10khz_RNIIENAZ0Z2\ : std_logic;
signal un2_counter_8 : std_logic;
signal un2_counter_7 : std_logic;
signal un2_counter_9 : std_logic;
signal clk_10khz_i : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_1\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_21_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_34\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_7\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_15\ : std_logic;
signal \bfn_7_21_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_23\ : std_logic;
signal \bfn_7_22_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_28\ : std_logic;
signal il_min_comp2_c : std_logic;
signal il_max_comp1_c : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_76\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_75\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \N_655_g\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_0\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_1_cry_0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_8\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_13\ : std_logic;
signal \current_shift_inst.control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_14\ : std_logic;
signal \current_shift_inst.control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_15\ : std_logic;
signal \current_shift_inst.control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_16\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_17\ : std_logic;
signal \current_shift_inst.control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_18\ : std_logic;
signal \current_shift_inst.control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_19\ : std_logic;
signal \current_shift_inst.control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_20\ : std_logic;
signal \current_shift_inst.control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_21\ : std_logic;
signal \current_shift_inst.control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_22\ : std_logic;
signal \current_shift_inst.control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_23\ : std_logic;
signal \current_shift_inst.control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_24\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \current_shift_inst.control_input_1_cry_24\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_8\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_16\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_24\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_phase.running_i\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \current_shift_inst.S1_syncZ0Z0\ : std_logic;
signal \current_shift_inst.S1_syncZ0Z1\ : std_logic;
signal \current_shift_inst.S1_sync_prevZ0\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \current_shift_inst.z_i_0_31\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_3_c_invZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_2\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_4\ : std_logic;
signal \current_shift_inst.control_input_1_axb_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_6\ : std_logic;
signal \current_shift_inst.control_input_1_axb_1\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8\ : std_logic;
signal \current_shift_inst.control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9\ : std_logic;
signal \current_shift_inst.control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10\ : std_logic;
signal \current_shift_inst.control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNILORI_11\ : std_logic;
signal \current_shift_inst.control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_11\ : std_logic;
signal \current_shift_inst.control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13\ : std_logic;
signal \current_shift_inst.control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_14\ : std_logic;
signal \current_shift_inst.control_input_1_axb_9\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_15\ : std_logic;
signal \current_shift_inst.control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIH6661_17\ : std_logic;
signal \current_shift_inst.control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIE6961_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18\ : std_logic;
signal \current_shift_inst.control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPC571_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19\ : std_logic;
signal \current_shift_inst.control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIDR081_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20\ : std_logic;
signal \current_shift_inst.control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21\ : std_logic;
signal \current_shift_inst.control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIR32K_22\ : std_logic;
signal \current_shift_inst.control_input_1_axb_17\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_23\ : std_logic;
signal \current_shift_inst.control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_24\ : std_logic;
signal \current_shift_inst.control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26\ : std_logic;
signal \current_shift_inst.control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINKG81_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27\ : std_logic;
signal \current_shift_inst.control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28\ : std_logic;
signal \current_shift_inst.control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\ : std_logic;
signal \current_shift_inst.control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_30\ : std_logic;
signal \current_shift_inst.control_input_1_cry_24_THRU_CO\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_25\ : std_logic;
signal \current_shift_inst.phase_valid_RNISLORZ0Z2\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \current_shift_inst.z_5_cry_1\ : std_logic;
signal \current_shift_inst.z_5_cry_2\ : std_logic;
signal \current_shift_inst.z_5_cry_3\ : std_logic;
signal \current_shift_inst.z_5_cry_4\ : std_logic;
signal \current_shift_inst.z_5_cry_5\ : std_logic;
signal \current_shift_inst.z_5_cry_6\ : std_logic;
signal \current_shift_inst.z_5_cry_7\ : std_logic;
signal \current_shift_inst.z_5_cry_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_9\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_10\ : std_logic;
signal \current_shift_inst.z_5_cry_9\ : std_logic;
signal \current_shift_inst.z_5_cry_10\ : std_logic;
signal \current_shift_inst.z_5_cry_11\ : std_logic;
signal \current_shift_inst.z_5_cry_12\ : std_logic;
signal \current_shift_inst.z_5_cry_13\ : std_logic;
signal \current_shift_inst.z_5_cry_14\ : std_logic;
signal \current_shift_inst.z_5_cry_15\ : std_logic;
signal \current_shift_inst.z_5_cry_16\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_18\ : std_logic;
signal \current_shift_inst.z_5_cry_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_19\ : std_logic;
signal \current_shift_inst.z_5_cry_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_20\ : std_logic;
signal \current_shift_inst.z_5_cry_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_21\ : std_logic;
signal \current_shift_inst.z_5_cry_20\ : std_logic;
signal \current_shift_inst.z_5_cry_21\ : std_logic;
signal \current_shift_inst.z_5_cry_22\ : std_logic;
signal \current_shift_inst.z_5_cry_23\ : std_logic;
signal \current_shift_inst.z_5_cry_24\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \current_shift_inst.z_5_cry_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_27\ : std_logic;
signal \current_shift_inst.z_5_cry_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_28\ : std_logic;
signal \current_shift_inst.z_5_cry_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_29\ : std_logic;
signal \current_shift_inst.z_5_cry_28\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.z_5_cry_29\ : std_logic;
signal \current_shift_inst.z_5_cry_30\ : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_5_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13_cascade_\ : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal measured_delay_hc_22 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30_2_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIER9V_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5M161_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI190J_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIBU361_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.N_1633_i\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_0\ : std_logic;
signal \current_shift_inst.timer_phase.N_188_i_g\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3_cascade_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0\ : std_logic;
signal \G_406\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_1\ : std_logic;
signal \G_405\ : std_logic;
signal \current_shift_inst.z_cry_0\ : std_logic;
signal \current_shift_inst.z_5_2\ : std_logic;
signal \current_shift_inst.z_cry_1\ : std_logic;
signal \current_shift_inst.z_5_3\ : std_logic;
signal \current_shift_inst.z_cry_2\ : std_logic;
signal \current_shift_inst.z_5_4\ : std_logic;
signal \current_shift_inst.z_cry_3\ : std_logic;
signal \current_shift_inst.z_5_5\ : std_logic;
signal \current_shift_inst.z_cry_4\ : std_logic;
signal \current_shift_inst.z_5_6\ : std_logic;
signal \current_shift_inst.z_cry_5\ : std_logic;
signal \current_shift_inst.z_5_7\ : std_logic;
signal \current_shift_inst.z_cry_6\ : std_logic;
signal \current_shift_inst.z_cry_7\ : std_logic;
signal \current_shift_inst.z_5_8\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \current_shift_inst.z_5_9\ : std_logic;
signal \current_shift_inst.z_cry_8\ : std_logic;
signal \current_shift_inst.z_5_10\ : std_logic;
signal \current_shift_inst.z_cry_9\ : std_logic;
signal \current_shift_inst.z_5_11\ : std_logic;
signal \current_shift_inst.z_cry_10\ : std_logic;
signal \current_shift_inst.z_5_12\ : std_logic;
signal \current_shift_inst.z_cry_11\ : std_logic;
signal \current_shift_inst.z_5_13\ : std_logic;
signal \current_shift_inst.z_cry_12\ : std_logic;
signal \current_shift_inst.z_5_14\ : std_logic;
signal \current_shift_inst.z_cry_13\ : std_logic;
signal \current_shift_inst.z_5_15\ : std_logic;
signal \current_shift_inst.z_cry_14\ : std_logic;
signal \current_shift_inst.z_cry_15\ : std_logic;
signal \current_shift_inst.z_5_16\ : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal \current_shift_inst.z_5_17\ : std_logic;
signal \current_shift_inst.z_cry_16\ : std_logic;
signal \current_shift_inst.z_5_18\ : std_logic;
signal \current_shift_inst.z_cry_17\ : std_logic;
signal \current_shift_inst.z_5_19\ : std_logic;
signal \current_shift_inst.z_cry_18\ : std_logic;
signal \current_shift_inst.z_5_20\ : std_logic;
signal \current_shift_inst.z_cry_19\ : std_logic;
signal \current_shift_inst.z_5_21\ : std_logic;
signal \current_shift_inst.z_cry_20\ : std_logic;
signal \current_shift_inst.z_5_22\ : std_logic;
signal \current_shift_inst.z_cry_21\ : std_logic;
signal \current_shift_inst.z_5_23\ : std_logic;
signal \current_shift_inst.z_cry_22\ : std_logic;
signal \current_shift_inst.z_cry_23\ : std_logic;
signal \current_shift_inst.z_5_24\ : std_logic;
signal \bfn_10_20_0_\ : std_logic;
signal \current_shift_inst.z_5_25\ : std_logic;
signal \current_shift_inst.z_cry_24\ : std_logic;
signal \current_shift_inst.z_5_26\ : std_logic;
signal \current_shift_inst.z_cry_25\ : std_logic;
signal \current_shift_inst.z_5_27\ : std_logic;
signal \current_shift_inst.z_cry_26\ : std_logic;
signal \current_shift_inst.z_5_28\ : std_logic;
signal \current_shift_inst.z_cry_27\ : std_logic;
signal \current_shift_inst.z_5_29\ : std_logic;
signal \current_shift_inst.z_cry_28\ : std_logic;
signal \current_shift_inst.z_5_30\ : std_logic;
signal \current_shift_inst.z_cry_29\ : std_logic;
signal \current_shift_inst.z_5_cry_30_THRU_CO\ : std_logic;
signal \current_shift_inst.z_cry_30\ : std_logic;
signal measured_delay_hc_21 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0_cascade_\ : std_logic;
signal measured_delay_hc_20 : std_logic;
signal measured_delay_hc_23 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlt30_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.N_187_i\ : std_logic;
signal \current_shift_inst.phase_validZ0\ : std_logic;
signal measured_delay_hc_27 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_fast_31\ : std_logic;
signal \current_shift_inst.un38_control_input_0\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_24\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5S981_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24\ : std_logic;
signal \current_shift_inst.z_31\ : std_logic;
signal \current_shift_inst.z_i_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_24\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIU73K_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_31\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_axb_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_26\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_22\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPB581_22\ : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto9_cZ0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \bfn_12_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\ : std_logic;
signal \current_shift_inst.S3_sync_prevZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt15\ : std_logic;
signal \current_shift_inst.S3_riseZ0\ : std_logic;
signal \current_shift_inst.S1_riseZ0\ : std_logic;
signal \current_shift_inst.N_199\ : std_logic;
signal \current_shift_inst.meas_stateZ0Z_0\ : std_logic;
signal measured_delay_hc_28 : std_logic;
signal measured_delay_hc_29 : std_logic;
signal measured_delay_hc_30 : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_3\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.N_187_i_g\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_29\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_28\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_20\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_30\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_19\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_19\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_26\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_27\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_27\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_25\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_22\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_12_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_12_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_191_i\ : std_logic;
signal \current_shift_inst.timer_phase.N_188_i\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal measured_delay_hc_25 : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal measured_delay_hc_26 : std_logic;
signal measured_delay_hc_24 : std_logic;
signal s1_phy_c : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \delay_measurement_inst.prev_hc_sigZ0\ : std_logic;
signal \delay_measurement_inst.hc_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.N_221_0\ : std_logic;
signal \current_shift_inst.S3_syncZ0Z1\ : std_logic;
signal \current_shift_inst.S3_syncZ0Z0\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_24\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_15\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_16\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_17\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_21\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_10\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_11\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_11\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_12\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_18\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_13\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_14\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_321_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_320_4\ : std_logic;
signal \delay_measurement_inst.N_305_1_cascade_\ : std_logic;
signal \delay_measurement_inst.N_305_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_299\ : std_logic;
signal \delay_measurement_inst.N_358_cascade_\ : std_logic;
signal \current_shift_inst.stop_timer_phaseZ0\ : std_logic;
signal \current_shift_inst.start_timer_phaseZ0\ : std_logic;
signal \current_shift_inst.timer_phase.runningZ0\ : std_logic;
signal \current_shift_inst.timer_phase.N_192_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_296\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_293_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\ : std_logic;
signal \delay_measurement_inst.N_307\ : std_logic;
signal s2_phy_c : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_335_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_14_5_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\ : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_N_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_1\ : std_logic;
signal delay_hc_d2 : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_3\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal measured_delay_hc_18 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30_2\ : std_logic;
signal red_c_i : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.N_232\ : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_slave.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.N_214\ : std_logic;
signal s4_phy_c : std_logic;
signal \phase_controller_slave.stateZ0Z_2\ : std_logic;
signal \phase_controller_slave.hc_time_passed\ : std_logic;
signal s3_phy_c : std_logic;
signal \phase_controller_slave.N_211_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa_cascade_\ : std_logic;
signal \phase_controller_slave.tr_time_passed\ : std_logic;
signal \phase_controller_slave.stateZ0Z_0\ : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \phase_controller_slave.N_211\ : std_logic;
signal \phase_controller_slave.stateZ0Z_3\ : std_logic;
signal \delay_measurement_inst.tr_stateZ0Z_0\ : std_logic;
signal \delay_measurement_inst.prev_tr_sigZ0\ : std_logic;
signal start_stop_c : std_logic;
signal shift_flag_start : std_logic;
signal \phase_controller_slave.stateZ0Z_4\ : std_logic;
signal \phase_controller_slave.N_213\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_slave.stateZ0Z_1\ : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \phase_controller_slave.start_timer_tr_0_sqmuxa\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6_cascade_\ : std_logic;
signal \delay_measurement_inst.N_358\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_331\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_331_cascade_\ : std_logic;
signal \delay_measurement_inst.N_333_cascade_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.N_333\ : std_logic;
signal \delay_measurement_inst.N_328\ : std_logic;
signal \delay_measurement_inst.N_324\ : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_3\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_11\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_19\ : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_337_i\ : std_logic;
signal delay_tr_input_c : std_logic;
signal delay_tr_d1 : std_logic;
signal delay_tr_d2 : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.N_228\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal measured_delay_hc_11 : std_logic;
signal measured_delay_hc_12 : std_logic;
signal measured_delay_hc_19 : std_logic;
signal measured_delay_hc_17 : std_logic;
signal measured_delay_hc_9 : std_logic;
signal measured_delay_hc_0 : std_logic;
signal measured_delay_hc_6 : std_logic;
signal measured_delay_hc_1 : std_logic;
signal measured_delay_hc_3 : std_logic;
signal measured_delay_hc_4 : std_logic;
signal measured_delay_hc_16 : std_logic;
signal measured_delay_hc_14 : std_logic;
signal measured_delay_hc_10 : std_logic;
signal measured_delay_hc_8 : std_logic;
signal measured_delay_hc_31 : std_logic;
signal measured_delay_hc_5 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt31_0\ : std_logic;
signal measured_delay_hc_13 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal measured_delay_hc_7 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_338_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_5_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt13_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclt31_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lt31_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_16_12_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_16_13_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\ : std_logic;
signal \delay_measurement_inst.N_284_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto15\ : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_tr_0_i\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\ : std_logic;
signal measured_delay_tr_8 : std_logic;
signal measured_delay_tr_2 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\ : std_logic;
signal measured_delay_tr_1 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_20_li\ : std_logic;
signal measured_delay_tr_3 : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_16_18_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_16_20_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal delay_hc_input_c : std_logic;
signal delay_hc_d1 : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto31_0_0\ : std_logic;
signal measured_delay_hc_2 : std_logic;
signal \delay_measurement_inst.un1_elapsed_time_hc\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3\ : std_logic;
signal measured_delay_hc_15 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_3\ : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_11\ : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_19\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_335_i_g\ : std_logic;
signal \phase_controller_slave.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_4\ : std_logic;
signal \phase_controller_inst1.N_231\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal measured_delay_tr_7 : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal measured_delay_tr_14 : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal measured_delay_tr_6 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal measured_delay_tr_11 : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal measured_delay_tr_12 : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal measured_delay_tr_13 : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\ : std_logic;
signal measured_delay_tr_15 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\ : std_logic;
signal measured_delay_tr_10 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_18_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_18_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_18_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_18_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_336_i\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_18_11_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\ : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\ : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_slave.start_timer_trZ0\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal red_c_g : std_logic;
signal measured_delay_tr_18 : std_logic;
signal measured_delay_tr_17 : std_logic;
signal measured_delay_tr_19 : std_logic;
signal measured_delay_tr_16 : std_logic;
signal measured_delay_tr_5 : std_logic;
signal measured_delay_tr_4 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_21\ : std_logic;
signal measured_delay_tr_9 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal reset_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ <= '0'&\N__18556\&\N__18560\&\N__18557\&\N__18561\&\N__18558\&\N__18605\&\N__18584\&\N__18260\&\N__20513\&\N__18242\&\N__18451\&\N__18349\&\N__18399\&\N__18417\&\N__18380\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__27715\&\N__27712\&'0'&'0'&'0'&\N__27710\&\N__27714\&\N__27711\&\N__27713\;
    \pwm_generator_inst.un2_threshold_acc_1_25\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_acc_1_24\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_acc_1_23\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_acc_1_22\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_acc_1_21\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_acc_1_20\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_acc_1_19\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_acc_1_18\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_acc_1_17\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_acc_1_16\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_1_15\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold_acc\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__18533\&\N__18526\&\N__18531\&\N__18525\&\N__18532\&\N__18524\&\N__18534\&\N__18521\&\N__18527\&\N__18520\&\N__18528\&\N__18522\&\N__18529\&\N__18523\&\N__18530\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__27837\&\N__27833\&'0'&'0'&'0'&\N__27831\&\N__27836\&\N__27832\&\N__27835\;
    \pwm_generator_inst.un2_threshold_acc_2_1_16\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_2_1_15\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_acc_2_14\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_acc_2_13\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_acc_2_12\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_acc_2_11\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_acc_2_10\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_acc_2_9\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_acc_2_8\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_acc_2_7\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_acc_2_6\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_acc_2_5\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_acc_2_4\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_acc_2_3\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_acc_2_2\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_acc_2_1\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_acc_2_0\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__32628\,
            RESETB => \N__34797\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__27778\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__27709\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__27834\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__27830\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__48094\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48096\,
            DIN => \N__48095\,
            DOUT => \N__48094\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48096\,
            PADOUT => \N__48095\,
            PADIN => \N__48094\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48085\,
            DIN => \N__48084\,
            DOUT => \N__48083\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48085\,
            PADOUT => \N__48084\,
            PADIN => \N__48083\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48076\,
            DIN => \N__48075\,
            DOUT => \N__48074\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48076\,
            PADOUT => \N__48075\,
            PADIN => \N__48074\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48067\,
            DIN => \N__48066\,
            DOUT => \N__48065\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48067\,
            PADOUT => \N__48066\,
            PADIN => \N__48065\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23682\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48058\,
            DIN => \N__48057\,
            DOUT => \N__48056\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48058\,
            PADOUT => \N__48057\,
            PADIN => \N__48056\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48049\,
            DIN => \N__48048\,
            DOUT => \N__48047\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48049\,
            PADOUT => \N__48048\,
            PADIN => \N__48047\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33861\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48040\,
            DIN => \N__48039\,
            DOUT => \N__48038\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48040\,
            PADOUT => \N__48039\,
            PADIN => \N__48038\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48031\,
            DIN => \N__48030\,
            DOUT => \N__48029\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48031\,
            PADOUT => \N__48030\,
            PADIN => \N__48029\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48022\,
            DIN => \N__48021\,
            DOUT => \N__48020\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48022\,
            PADOUT => \N__48021\,
            PADIN => \N__48020\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48013\,
            DIN => \N__48012\,
            DOUT => \N__48011\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48013\,
            PADOUT => \N__48012\,
            PADIN => \N__48011\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32934\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48004\,
            DIN => \N__48003\,
            DOUT => \N__48002\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48004\,
            PADOUT => \N__48003\,
            PADIN => \N__48002\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34902\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47995\,
            DIN => \N__47994\,
            DOUT => \N__47993\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__47995\,
            PADOUT => \N__47994\,
            PADIN => \N__47993\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__47986\,
            DIN => \N__47985\,
            DOUT => \N__47984\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__47986\,
            PADOUT => \N__47985\,
            PADIN => \N__47984\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34836\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11450\ : InMux
    port map (
            O => \N__47967\,
            I => \N__47964\
        );

    \I__11449\ : LocalMux
    port map (
            O => \N__47964\,
            I => \N__47961\
        );

    \I__11448\ : Odrv4
    port map (
            O => \N__47961\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\
        );

    \I__11447\ : InMux
    port map (
            O => \N__47958\,
            I => \N__47954\
        );

    \I__11446\ : InMux
    port map (
            O => \N__47957\,
            I => \N__47951\
        );

    \I__11445\ : LocalMux
    port map (
            O => \N__47954\,
            I => \N__47948\
        );

    \I__11444\ : LocalMux
    port map (
            O => \N__47951\,
            I => \N__47945\
        );

    \I__11443\ : Odrv12
    port map (
            O => \N__47948\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__11442\ : Odrv4
    port map (
            O => \N__47945\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__11441\ : CascadeMux
    port map (
            O => \N__47940\,
            I => \N__47933\
        );

    \I__11440\ : CascadeMux
    port map (
            O => \N__47939\,
            I => \N__47927\
        );

    \I__11439\ : CascadeMux
    port map (
            O => \N__47938\,
            I => \N__47918\
        );

    \I__11438\ : CascadeMux
    port map (
            O => \N__47937\,
            I => \N__47915\
        );

    \I__11437\ : CascadeMux
    port map (
            O => \N__47936\,
            I => \N__47912\
        );

    \I__11436\ : InMux
    port map (
            O => \N__47933\,
            I => \N__47901\
        );

    \I__11435\ : InMux
    port map (
            O => \N__47932\,
            I => \N__47901\
        );

    \I__11434\ : CascadeMux
    port map (
            O => \N__47931\,
            I => \N__47896\
        );

    \I__11433\ : CascadeMux
    port map (
            O => \N__47930\,
            I => \N__47893\
        );

    \I__11432\ : InMux
    port map (
            O => \N__47927\,
            I => \N__47886\
        );

    \I__11431\ : InMux
    port map (
            O => \N__47926\,
            I => \N__47886\
        );

    \I__11430\ : InMux
    port map (
            O => \N__47925\,
            I => \N__47883\
        );

    \I__11429\ : InMux
    port map (
            O => \N__47924\,
            I => \N__47880\
        );

    \I__11428\ : InMux
    port map (
            O => \N__47923\,
            I => \N__47867\
        );

    \I__11427\ : InMux
    port map (
            O => \N__47922\,
            I => \N__47867\
        );

    \I__11426\ : InMux
    port map (
            O => \N__47921\,
            I => \N__47867\
        );

    \I__11425\ : InMux
    port map (
            O => \N__47918\,
            I => \N__47867\
        );

    \I__11424\ : InMux
    port map (
            O => \N__47915\,
            I => \N__47867\
        );

    \I__11423\ : InMux
    port map (
            O => \N__47912\,
            I => \N__47867\
        );

    \I__11422\ : InMux
    port map (
            O => \N__47911\,
            I => \N__47854\
        );

    \I__11421\ : InMux
    port map (
            O => \N__47910\,
            I => \N__47854\
        );

    \I__11420\ : InMux
    port map (
            O => \N__47909\,
            I => \N__47854\
        );

    \I__11419\ : InMux
    port map (
            O => \N__47908\,
            I => \N__47854\
        );

    \I__11418\ : InMux
    port map (
            O => \N__47907\,
            I => \N__47854\
        );

    \I__11417\ : InMux
    port map (
            O => \N__47906\,
            I => \N__47854\
        );

    \I__11416\ : LocalMux
    port map (
            O => \N__47901\,
            I => \N__47851\
        );

    \I__11415\ : InMux
    port map (
            O => \N__47900\,
            I => \N__47848\
        );

    \I__11414\ : CascadeMux
    port map (
            O => \N__47899\,
            I => \N__47845\
        );

    \I__11413\ : InMux
    port map (
            O => \N__47896\,
            I => \N__47836\
        );

    \I__11412\ : InMux
    port map (
            O => \N__47893\,
            I => \N__47836\
        );

    \I__11411\ : InMux
    port map (
            O => \N__47892\,
            I => \N__47836\
        );

    \I__11410\ : InMux
    port map (
            O => \N__47891\,
            I => \N__47836\
        );

    \I__11409\ : LocalMux
    port map (
            O => \N__47886\,
            I => \N__47833\
        );

    \I__11408\ : LocalMux
    port map (
            O => \N__47883\,
            I => \N__47830\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__47880\,
            I => \N__47823\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__47867\,
            I => \N__47823\
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__47854\,
            I => \N__47823\
        );

    \I__11404\ : Span4Mux_v
    port map (
            O => \N__47851\,
            I => \N__47820\
        );

    \I__11403\ : LocalMux
    port map (
            O => \N__47848\,
            I => \N__47817\
        );

    \I__11402\ : InMux
    port map (
            O => \N__47845\,
            I => \N__47814\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__47836\,
            I => \N__47809\
        );

    \I__11400\ : Span4Mux_v
    port map (
            O => \N__47833\,
            I => \N__47809\
        );

    \I__11399\ : Span4Mux_v
    port map (
            O => \N__47830\,
            I => \N__47804\
        );

    \I__11398\ : Span4Mux_v
    port map (
            O => \N__47823\,
            I => \N__47804\
        );

    \I__11397\ : Span4Mux_h
    port map (
            O => \N__47820\,
            I => \N__47799\
        );

    \I__11396\ : Span4Mux_h
    port map (
            O => \N__47817\,
            I => \N__47799\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__47814\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__11394\ : Odrv4
    port map (
            O => \N__47809\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__11393\ : Odrv4
    port map (
            O => \N__47804\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__11392\ : Odrv4
    port map (
            O => \N__47799\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__11391\ : CascadeMux
    port map (
            O => \N__47790\,
            I => \N__47786\
        );

    \I__11390\ : InMux
    port map (
            O => \N__47789\,
            I => \N__47759\
        );

    \I__11389\ : InMux
    port map (
            O => \N__47786\,
            I => \N__47759\
        );

    \I__11388\ : InMux
    port map (
            O => \N__47785\,
            I => \N__47759\
        );

    \I__11387\ : InMux
    port map (
            O => \N__47784\,
            I => \N__47759\
        );

    \I__11386\ : InMux
    port map (
            O => \N__47783\,
            I => \N__47759\
        );

    \I__11385\ : InMux
    port map (
            O => \N__47782\,
            I => \N__47759\
        );

    \I__11384\ : InMux
    port map (
            O => \N__47781\,
            I => \N__47759\
        );

    \I__11383\ : InMux
    port map (
            O => \N__47780\,
            I => \N__47744\
        );

    \I__11382\ : InMux
    port map (
            O => \N__47779\,
            I => \N__47744\
        );

    \I__11381\ : InMux
    port map (
            O => \N__47778\,
            I => \N__47744\
        );

    \I__11380\ : InMux
    port map (
            O => \N__47777\,
            I => \N__47744\
        );

    \I__11379\ : InMux
    port map (
            O => \N__47776\,
            I => \N__47744\
        );

    \I__11378\ : InMux
    port map (
            O => \N__47775\,
            I => \N__47744\
        );

    \I__11377\ : InMux
    port map (
            O => \N__47774\,
            I => \N__47744\
        );

    \I__11376\ : LocalMux
    port map (
            O => \N__47759\,
            I => \N__47738\
        );

    \I__11375\ : LocalMux
    port map (
            O => \N__47744\,
            I => \N__47735\
        );

    \I__11374\ : CascadeMux
    port map (
            O => \N__47743\,
            I => \N__47731\
        );

    \I__11373\ : InMux
    port map (
            O => \N__47742\,
            I => \N__47726\
        );

    \I__11372\ : CascadeMux
    port map (
            O => \N__47741\,
            I => \N__47722\
        );

    \I__11371\ : Span4Mux_h
    port map (
            O => \N__47738\,
            I => \N__47716\
        );

    \I__11370\ : Span4Mux_v
    port map (
            O => \N__47735\,
            I => \N__47716\
        );

    \I__11369\ : InMux
    port map (
            O => \N__47734\,
            I => \N__47713\
        );

    \I__11368\ : InMux
    port map (
            O => \N__47731\,
            I => \N__47710\
        );

    \I__11367\ : InMux
    port map (
            O => \N__47730\,
            I => \N__47705\
        );

    \I__11366\ : InMux
    port map (
            O => \N__47729\,
            I => \N__47705\
        );

    \I__11365\ : LocalMux
    port map (
            O => \N__47726\,
            I => \N__47702\
        );

    \I__11364\ : InMux
    port map (
            O => \N__47725\,
            I => \N__47699\
        );

    \I__11363\ : InMux
    port map (
            O => \N__47722\,
            I => \N__47696\
        );

    \I__11362\ : InMux
    port map (
            O => \N__47721\,
            I => \N__47693\
        );

    \I__11361\ : Span4Mux_v
    port map (
            O => \N__47716\,
            I => \N__47688\
        );

    \I__11360\ : LocalMux
    port map (
            O => \N__47713\,
            I => \N__47688\
        );

    \I__11359\ : LocalMux
    port map (
            O => \N__47710\,
            I => \N__47681\
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__47705\,
            I => \N__47681\
        );

    \I__11357\ : Span4Mux_h
    port map (
            O => \N__47702\,
            I => \N__47676\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__47699\,
            I => \N__47676\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__47696\,
            I => \N__47669\
        );

    \I__11354\ : LocalMux
    port map (
            O => \N__47693\,
            I => \N__47669\
        );

    \I__11353\ : Span4Mux_h
    port map (
            O => \N__47688\,
            I => \N__47669\
        );

    \I__11352\ : InMux
    port map (
            O => \N__47687\,
            I => \N__47664\
        );

    \I__11351\ : InMux
    port map (
            O => \N__47686\,
            I => \N__47664\
        );

    \I__11350\ : Span12Mux_h
    port map (
            O => \N__47681\,
            I => \N__47661\
        );

    \I__11349\ : Span4Mux_v
    port map (
            O => \N__47676\,
            I => \N__47658\
        );

    \I__11348\ : Span4Mux_v
    port map (
            O => \N__47669\,
            I => \N__47655\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__47664\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__11346\ : Odrv12
    port map (
            O => \N__47661\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__11345\ : Odrv4
    port map (
            O => \N__47658\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__11344\ : Odrv4
    port map (
            O => \N__47655\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__11343\ : CascadeMux
    port map (
            O => \N__47646\,
            I => \N__47643\
        );

    \I__11342\ : InMux
    port map (
            O => \N__47643\,
            I => \N__47640\
        );

    \I__11341\ : LocalMux
    port map (
            O => \N__47640\,
            I => \N__47637\
        );

    \I__11340\ : Span4Mux_h
    port map (
            O => \N__47637\,
            I => \N__47634\
        );

    \I__11339\ : Odrv4
    port map (
            O => \N__47634\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\
        );

    \I__11338\ : CascadeMux
    port map (
            O => \N__47631\,
            I => \N__47617\
        );

    \I__11337\ : CascadeMux
    port map (
            O => \N__47630\,
            I => \N__47612\
        );

    \I__11336\ : CascadeMux
    port map (
            O => \N__47629\,
            I => \N__47609\
        );

    \I__11335\ : CascadeMux
    port map (
            O => \N__47628\,
            I => \N__47606\
        );

    \I__11334\ : InMux
    port map (
            O => \N__47627\,
            I => \N__47590\
        );

    \I__11333\ : InMux
    port map (
            O => \N__47626\,
            I => \N__47590\
        );

    \I__11332\ : InMux
    port map (
            O => \N__47625\,
            I => \N__47590\
        );

    \I__11331\ : InMux
    port map (
            O => \N__47624\,
            I => \N__47590\
        );

    \I__11330\ : InMux
    port map (
            O => \N__47623\,
            I => \N__47590\
        );

    \I__11329\ : InMux
    port map (
            O => \N__47622\,
            I => \N__47590\
        );

    \I__11328\ : InMux
    port map (
            O => \N__47621\,
            I => \N__47590\
        );

    \I__11327\ : InMux
    port map (
            O => \N__47620\,
            I => \N__47585\
        );

    \I__11326\ : InMux
    port map (
            O => \N__47617\,
            I => \N__47585\
        );

    \I__11325\ : InMux
    port map (
            O => \N__47616\,
            I => \N__47574\
        );

    \I__11324\ : InMux
    port map (
            O => \N__47615\,
            I => \N__47574\
        );

    \I__11323\ : InMux
    port map (
            O => \N__47612\,
            I => \N__47574\
        );

    \I__11322\ : InMux
    port map (
            O => \N__47609\,
            I => \N__47574\
        );

    \I__11321\ : InMux
    port map (
            O => \N__47606\,
            I => \N__47574\
        );

    \I__11320\ : InMux
    port map (
            O => \N__47605\,
            I => \N__47566\
        );

    \I__11319\ : LocalMux
    port map (
            O => \N__47590\,
            I => \N__47563\
        );

    \I__11318\ : LocalMux
    port map (
            O => \N__47585\,
            I => \N__47558\
        );

    \I__11317\ : LocalMux
    port map (
            O => \N__47574\,
            I => \N__47558\
        );

    \I__11316\ : InMux
    port map (
            O => \N__47573\,
            I => \N__47551\
        );

    \I__11315\ : InMux
    port map (
            O => \N__47572\,
            I => \N__47551\
        );

    \I__11314\ : InMux
    port map (
            O => \N__47571\,
            I => \N__47551\
        );

    \I__11313\ : InMux
    port map (
            O => \N__47570\,
            I => \N__47546\
        );

    \I__11312\ : InMux
    port map (
            O => \N__47569\,
            I => \N__47546\
        );

    \I__11311\ : LocalMux
    port map (
            O => \N__47566\,
            I => \N__47543\
        );

    \I__11310\ : Span4Mux_h
    port map (
            O => \N__47563\,
            I => \N__47537\
        );

    \I__11309\ : Span4Mux_v
    port map (
            O => \N__47558\,
            I => \N__47537\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__47551\,
            I => \N__47532\
        );

    \I__11307\ : LocalMux
    port map (
            O => \N__47546\,
            I => \N__47527\
        );

    \I__11306\ : Span4Mux_v
    port map (
            O => \N__47543\,
            I => \N__47527\
        );

    \I__11305\ : InMux
    port map (
            O => \N__47542\,
            I => \N__47524\
        );

    \I__11304\ : Span4Mux_v
    port map (
            O => \N__47537\,
            I => \N__47521\
        );

    \I__11303\ : InMux
    port map (
            O => \N__47536\,
            I => \N__47518\
        );

    \I__11302\ : CascadeMux
    port map (
            O => \N__47535\,
            I => \N__47515\
        );

    \I__11301\ : Span4Mux_v
    port map (
            O => \N__47532\,
            I => \N__47511\
        );

    \I__11300\ : Span4Mux_h
    port map (
            O => \N__47527\,
            I => \N__47506\
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__47524\,
            I => \N__47506\
        );

    \I__11298\ : Sp12to4
    port map (
            O => \N__47521\,
            I => \N__47501\
        );

    \I__11297\ : LocalMux
    port map (
            O => \N__47518\,
            I => \N__47501\
        );

    \I__11296\ : InMux
    port map (
            O => \N__47515\,
            I => \N__47496\
        );

    \I__11295\ : InMux
    port map (
            O => \N__47514\,
            I => \N__47496\
        );

    \I__11294\ : Span4Mux_h
    port map (
            O => \N__47511\,
            I => \N__47491\
        );

    \I__11293\ : Span4Mux_v
    port map (
            O => \N__47506\,
            I => \N__47491\
        );

    \I__11292\ : Span12Mux_h
    port map (
            O => \N__47501\,
            I => \N__47488\
        );

    \I__11291\ : LocalMux
    port map (
            O => \N__47496\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__11290\ : Odrv4
    port map (
            O => \N__47491\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__11289\ : Odrv12
    port map (
            O => \N__47488\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__11288\ : InMux
    port map (
            O => \N__47481\,
            I => \N__47477\
        );

    \I__11287\ : InMux
    port map (
            O => \N__47480\,
            I => \N__47474\
        );

    \I__11286\ : LocalMux
    port map (
            O => \N__47477\,
            I => \N__47471\
        );

    \I__11285\ : LocalMux
    port map (
            O => \N__47474\,
            I => \N__47468\
        );

    \I__11284\ : Odrv12
    port map (
            O => \N__47471\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__11283\ : Odrv4
    port map (
            O => \N__47468\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__11282\ : ClkMux
    port map (
            O => \N__47463\,
            I => \N__46992\
        );

    \I__11281\ : ClkMux
    port map (
            O => \N__47462\,
            I => \N__46992\
        );

    \I__11280\ : ClkMux
    port map (
            O => \N__47461\,
            I => \N__46992\
        );

    \I__11279\ : ClkMux
    port map (
            O => \N__47460\,
            I => \N__46992\
        );

    \I__11278\ : ClkMux
    port map (
            O => \N__47459\,
            I => \N__46992\
        );

    \I__11277\ : ClkMux
    port map (
            O => \N__47458\,
            I => \N__46992\
        );

    \I__11276\ : ClkMux
    port map (
            O => \N__47457\,
            I => \N__46992\
        );

    \I__11275\ : ClkMux
    port map (
            O => \N__47456\,
            I => \N__46992\
        );

    \I__11274\ : ClkMux
    port map (
            O => \N__47455\,
            I => \N__46992\
        );

    \I__11273\ : ClkMux
    port map (
            O => \N__47454\,
            I => \N__46992\
        );

    \I__11272\ : ClkMux
    port map (
            O => \N__47453\,
            I => \N__46992\
        );

    \I__11271\ : ClkMux
    port map (
            O => \N__47452\,
            I => \N__46992\
        );

    \I__11270\ : ClkMux
    port map (
            O => \N__47451\,
            I => \N__46992\
        );

    \I__11269\ : ClkMux
    port map (
            O => \N__47450\,
            I => \N__46992\
        );

    \I__11268\ : ClkMux
    port map (
            O => \N__47449\,
            I => \N__46992\
        );

    \I__11267\ : ClkMux
    port map (
            O => \N__47448\,
            I => \N__46992\
        );

    \I__11266\ : ClkMux
    port map (
            O => \N__47447\,
            I => \N__46992\
        );

    \I__11265\ : ClkMux
    port map (
            O => \N__47446\,
            I => \N__46992\
        );

    \I__11264\ : ClkMux
    port map (
            O => \N__47445\,
            I => \N__46992\
        );

    \I__11263\ : ClkMux
    port map (
            O => \N__47444\,
            I => \N__46992\
        );

    \I__11262\ : ClkMux
    port map (
            O => \N__47443\,
            I => \N__46992\
        );

    \I__11261\ : ClkMux
    port map (
            O => \N__47442\,
            I => \N__46992\
        );

    \I__11260\ : ClkMux
    port map (
            O => \N__47441\,
            I => \N__46992\
        );

    \I__11259\ : ClkMux
    port map (
            O => \N__47440\,
            I => \N__46992\
        );

    \I__11258\ : ClkMux
    port map (
            O => \N__47439\,
            I => \N__46992\
        );

    \I__11257\ : ClkMux
    port map (
            O => \N__47438\,
            I => \N__46992\
        );

    \I__11256\ : ClkMux
    port map (
            O => \N__47437\,
            I => \N__46992\
        );

    \I__11255\ : ClkMux
    port map (
            O => \N__47436\,
            I => \N__46992\
        );

    \I__11254\ : ClkMux
    port map (
            O => \N__47435\,
            I => \N__46992\
        );

    \I__11253\ : ClkMux
    port map (
            O => \N__47434\,
            I => \N__46992\
        );

    \I__11252\ : ClkMux
    port map (
            O => \N__47433\,
            I => \N__46992\
        );

    \I__11251\ : ClkMux
    port map (
            O => \N__47432\,
            I => \N__46992\
        );

    \I__11250\ : ClkMux
    port map (
            O => \N__47431\,
            I => \N__46992\
        );

    \I__11249\ : ClkMux
    port map (
            O => \N__47430\,
            I => \N__46992\
        );

    \I__11248\ : ClkMux
    port map (
            O => \N__47429\,
            I => \N__46992\
        );

    \I__11247\ : ClkMux
    port map (
            O => \N__47428\,
            I => \N__46992\
        );

    \I__11246\ : ClkMux
    port map (
            O => \N__47427\,
            I => \N__46992\
        );

    \I__11245\ : ClkMux
    port map (
            O => \N__47426\,
            I => \N__46992\
        );

    \I__11244\ : ClkMux
    port map (
            O => \N__47425\,
            I => \N__46992\
        );

    \I__11243\ : ClkMux
    port map (
            O => \N__47424\,
            I => \N__46992\
        );

    \I__11242\ : ClkMux
    port map (
            O => \N__47423\,
            I => \N__46992\
        );

    \I__11241\ : ClkMux
    port map (
            O => \N__47422\,
            I => \N__46992\
        );

    \I__11240\ : ClkMux
    port map (
            O => \N__47421\,
            I => \N__46992\
        );

    \I__11239\ : ClkMux
    port map (
            O => \N__47420\,
            I => \N__46992\
        );

    \I__11238\ : ClkMux
    port map (
            O => \N__47419\,
            I => \N__46992\
        );

    \I__11237\ : ClkMux
    port map (
            O => \N__47418\,
            I => \N__46992\
        );

    \I__11236\ : ClkMux
    port map (
            O => \N__47417\,
            I => \N__46992\
        );

    \I__11235\ : ClkMux
    port map (
            O => \N__47416\,
            I => \N__46992\
        );

    \I__11234\ : ClkMux
    port map (
            O => \N__47415\,
            I => \N__46992\
        );

    \I__11233\ : ClkMux
    port map (
            O => \N__47414\,
            I => \N__46992\
        );

    \I__11232\ : ClkMux
    port map (
            O => \N__47413\,
            I => \N__46992\
        );

    \I__11231\ : ClkMux
    port map (
            O => \N__47412\,
            I => \N__46992\
        );

    \I__11230\ : ClkMux
    port map (
            O => \N__47411\,
            I => \N__46992\
        );

    \I__11229\ : ClkMux
    port map (
            O => \N__47410\,
            I => \N__46992\
        );

    \I__11228\ : ClkMux
    port map (
            O => \N__47409\,
            I => \N__46992\
        );

    \I__11227\ : ClkMux
    port map (
            O => \N__47408\,
            I => \N__46992\
        );

    \I__11226\ : ClkMux
    port map (
            O => \N__47407\,
            I => \N__46992\
        );

    \I__11225\ : ClkMux
    port map (
            O => \N__47406\,
            I => \N__46992\
        );

    \I__11224\ : ClkMux
    port map (
            O => \N__47405\,
            I => \N__46992\
        );

    \I__11223\ : ClkMux
    port map (
            O => \N__47404\,
            I => \N__46992\
        );

    \I__11222\ : ClkMux
    port map (
            O => \N__47403\,
            I => \N__46992\
        );

    \I__11221\ : ClkMux
    port map (
            O => \N__47402\,
            I => \N__46992\
        );

    \I__11220\ : ClkMux
    port map (
            O => \N__47401\,
            I => \N__46992\
        );

    \I__11219\ : ClkMux
    port map (
            O => \N__47400\,
            I => \N__46992\
        );

    \I__11218\ : ClkMux
    port map (
            O => \N__47399\,
            I => \N__46992\
        );

    \I__11217\ : ClkMux
    port map (
            O => \N__47398\,
            I => \N__46992\
        );

    \I__11216\ : ClkMux
    port map (
            O => \N__47397\,
            I => \N__46992\
        );

    \I__11215\ : ClkMux
    port map (
            O => \N__47396\,
            I => \N__46992\
        );

    \I__11214\ : ClkMux
    port map (
            O => \N__47395\,
            I => \N__46992\
        );

    \I__11213\ : ClkMux
    port map (
            O => \N__47394\,
            I => \N__46992\
        );

    \I__11212\ : ClkMux
    port map (
            O => \N__47393\,
            I => \N__46992\
        );

    \I__11211\ : ClkMux
    port map (
            O => \N__47392\,
            I => \N__46992\
        );

    \I__11210\ : ClkMux
    port map (
            O => \N__47391\,
            I => \N__46992\
        );

    \I__11209\ : ClkMux
    port map (
            O => \N__47390\,
            I => \N__46992\
        );

    \I__11208\ : ClkMux
    port map (
            O => \N__47389\,
            I => \N__46992\
        );

    \I__11207\ : ClkMux
    port map (
            O => \N__47388\,
            I => \N__46992\
        );

    \I__11206\ : ClkMux
    port map (
            O => \N__47387\,
            I => \N__46992\
        );

    \I__11205\ : ClkMux
    port map (
            O => \N__47386\,
            I => \N__46992\
        );

    \I__11204\ : ClkMux
    port map (
            O => \N__47385\,
            I => \N__46992\
        );

    \I__11203\ : ClkMux
    port map (
            O => \N__47384\,
            I => \N__46992\
        );

    \I__11202\ : ClkMux
    port map (
            O => \N__47383\,
            I => \N__46992\
        );

    \I__11201\ : ClkMux
    port map (
            O => \N__47382\,
            I => \N__46992\
        );

    \I__11200\ : ClkMux
    port map (
            O => \N__47381\,
            I => \N__46992\
        );

    \I__11199\ : ClkMux
    port map (
            O => \N__47380\,
            I => \N__46992\
        );

    \I__11198\ : ClkMux
    port map (
            O => \N__47379\,
            I => \N__46992\
        );

    \I__11197\ : ClkMux
    port map (
            O => \N__47378\,
            I => \N__46992\
        );

    \I__11196\ : ClkMux
    port map (
            O => \N__47377\,
            I => \N__46992\
        );

    \I__11195\ : ClkMux
    port map (
            O => \N__47376\,
            I => \N__46992\
        );

    \I__11194\ : ClkMux
    port map (
            O => \N__47375\,
            I => \N__46992\
        );

    \I__11193\ : ClkMux
    port map (
            O => \N__47374\,
            I => \N__46992\
        );

    \I__11192\ : ClkMux
    port map (
            O => \N__47373\,
            I => \N__46992\
        );

    \I__11191\ : ClkMux
    port map (
            O => \N__47372\,
            I => \N__46992\
        );

    \I__11190\ : ClkMux
    port map (
            O => \N__47371\,
            I => \N__46992\
        );

    \I__11189\ : ClkMux
    port map (
            O => \N__47370\,
            I => \N__46992\
        );

    \I__11188\ : ClkMux
    port map (
            O => \N__47369\,
            I => \N__46992\
        );

    \I__11187\ : ClkMux
    port map (
            O => \N__47368\,
            I => \N__46992\
        );

    \I__11186\ : ClkMux
    port map (
            O => \N__47367\,
            I => \N__46992\
        );

    \I__11185\ : ClkMux
    port map (
            O => \N__47366\,
            I => \N__46992\
        );

    \I__11184\ : ClkMux
    port map (
            O => \N__47365\,
            I => \N__46992\
        );

    \I__11183\ : ClkMux
    port map (
            O => \N__47364\,
            I => \N__46992\
        );

    \I__11182\ : ClkMux
    port map (
            O => \N__47363\,
            I => \N__46992\
        );

    \I__11181\ : ClkMux
    port map (
            O => \N__47362\,
            I => \N__46992\
        );

    \I__11180\ : ClkMux
    port map (
            O => \N__47361\,
            I => \N__46992\
        );

    \I__11179\ : ClkMux
    port map (
            O => \N__47360\,
            I => \N__46992\
        );

    \I__11178\ : ClkMux
    port map (
            O => \N__47359\,
            I => \N__46992\
        );

    \I__11177\ : ClkMux
    port map (
            O => \N__47358\,
            I => \N__46992\
        );

    \I__11176\ : ClkMux
    port map (
            O => \N__47357\,
            I => \N__46992\
        );

    \I__11175\ : ClkMux
    port map (
            O => \N__47356\,
            I => \N__46992\
        );

    \I__11174\ : ClkMux
    port map (
            O => \N__47355\,
            I => \N__46992\
        );

    \I__11173\ : ClkMux
    port map (
            O => \N__47354\,
            I => \N__46992\
        );

    \I__11172\ : ClkMux
    port map (
            O => \N__47353\,
            I => \N__46992\
        );

    \I__11171\ : ClkMux
    port map (
            O => \N__47352\,
            I => \N__46992\
        );

    \I__11170\ : ClkMux
    port map (
            O => \N__47351\,
            I => \N__46992\
        );

    \I__11169\ : ClkMux
    port map (
            O => \N__47350\,
            I => \N__46992\
        );

    \I__11168\ : ClkMux
    port map (
            O => \N__47349\,
            I => \N__46992\
        );

    \I__11167\ : ClkMux
    port map (
            O => \N__47348\,
            I => \N__46992\
        );

    \I__11166\ : ClkMux
    port map (
            O => \N__47347\,
            I => \N__46992\
        );

    \I__11165\ : ClkMux
    port map (
            O => \N__47346\,
            I => \N__46992\
        );

    \I__11164\ : ClkMux
    port map (
            O => \N__47345\,
            I => \N__46992\
        );

    \I__11163\ : ClkMux
    port map (
            O => \N__47344\,
            I => \N__46992\
        );

    \I__11162\ : ClkMux
    port map (
            O => \N__47343\,
            I => \N__46992\
        );

    \I__11161\ : ClkMux
    port map (
            O => \N__47342\,
            I => \N__46992\
        );

    \I__11160\ : ClkMux
    port map (
            O => \N__47341\,
            I => \N__46992\
        );

    \I__11159\ : ClkMux
    port map (
            O => \N__47340\,
            I => \N__46992\
        );

    \I__11158\ : ClkMux
    port map (
            O => \N__47339\,
            I => \N__46992\
        );

    \I__11157\ : ClkMux
    port map (
            O => \N__47338\,
            I => \N__46992\
        );

    \I__11156\ : ClkMux
    port map (
            O => \N__47337\,
            I => \N__46992\
        );

    \I__11155\ : ClkMux
    port map (
            O => \N__47336\,
            I => \N__46992\
        );

    \I__11154\ : ClkMux
    port map (
            O => \N__47335\,
            I => \N__46992\
        );

    \I__11153\ : ClkMux
    port map (
            O => \N__47334\,
            I => \N__46992\
        );

    \I__11152\ : ClkMux
    port map (
            O => \N__47333\,
            I => \N__46992\
        );

    \I__11151\ : ClkMux
    port map (
            O => \N__47332\,
            I => \N__46992\
        );

    \I__11150\ : ClkMux
    port map (
            O => \N__47331\,
            I => \N__46992\
        );

    \I__11149\ : ClkMux
    port map (
            O => \N__47330\,
            I => \N__46992\
        );

    \I__11148\ : ClkMux
    port map (
            O => \N__47329\,
            I => \N__46992\
        );

    \I__11147\ : ClkMux
    port map (
            O => \N__47328\,
            I => \N__46992\
        );

    \I__11146\ : ClkMux
    port map (
            O => \N__47327\,
            I => \N__46992\
        );

    \I__11145\ : ClkMux
    port map (
            O => \N__47326\,
            I => \N__46992\
        );

    \I__11144\ : ClkMux
    port map (
            O => \N__47325\,
            I => \N__46992\
        );

    \I__11143\ : ClkMux
    port map (
            O => \N__47324\,
            I => \N__46992\
        );

    \I__11142\ : ClkMux
    port map (
            O => \N__47323\,
            I => \N__46992\
        );

    \I__11141\ : ClkMux
    port map (
            O => \N__47322\,
            I => \N__46992\
        );

    \I__11140\ : ClkMux
    port map (
            O => \N__47321\,
            I => \N__46992\
        );

    \I__11139\ : ClkMux
    port map (
            O => \N__47320\,
            I => \N__46992\
        );

    \I__11138\ : ClkMux
    port map (
            O => \N__47319\,
            I => \N__46992\
        );

    \I__11137\ : ClkMux
    port map (
            O => \N__47318\,
            I => \N__46992\
        );

    \I__11136\ : ClkMux
    port map (
            O => \N__47317\,
            I => \N__46992\
        );

    \I__11135\ : ClkMux
    port map (
            O => \N__47316\,
            I => \N__46992\
        );

    \I__11134\ : ClkMux
    port map (
            O => \N__47315\,
            I => \N__46992\
        );

    \I__11133\ : ClkMux
    port map (
            O => \N__47314\,
            I => \N__46992\
        );

    \I__11132\ : ClkMux
    port map (
            O => \N__47313\,
            I => \N__46992\
        );

    \I__11131\ : ClkMux
    port map (
            O => \N__47312\,
            I => \N__46992\
        );

    \I__11130\ : ClkMux
    port map (
            O => \N__47311\,
            I => \N__46992\
        );

    \I__11129\ : ClkMux
    port map (
            O => \N__47310\,
            I => \N__46992\
        );

    \I__11128\ : ClkMux
    port map (
            O => \N__47309\,
            I => \N__46992\
        );

    \I__11127\ : ClkMux
    port map (
            O => \N__47308\,
            I => \N__46992\
        );

    \I__11126\ : ClkMux
    port map (
            O => \N__47307\,
            I => \N__46992\
        );

    \I__11125\ : GlobalMux
    port map (
            O => \N__46992\,
            I => clk_100mhz_0
        );

    \I__11124\ : CascadeMux
    port map (
            O => \N__46989\,
            I => \N__46981\
        );

    \I__11123\ : CascadeMux
    port map (
            O => \N__46988\,
            I => \N__46978\
        );

    \I__11122\ : InMux
    port map (
            O => \N__46987\,
            I => \N__46974\
        );

    \I__11121\ : InMux
    port map (
            O => \N__46986\,
            I => \N__46971\
        );

    \I__11120\ : InMux
    port map (
            O => \N__46985\,
            I => \N__46968\
        );

    \I__11119\ : InMux
    port map (
            O => \N__46984\,
            I => \N__46965\
        );

    \I__11118\ : InMux
    port map (
            O => \N__46981\,
            I => \N__46962\
        );

    \I__11117\ : InMux
    port map (
            O => \N__46978\,
            I => \N__46959\
        );

    \I__11116\ : InMux
    port map (
            O => \N__46977\,
            I => \N__46956\
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__46974\,
            I => \N__46953\
        );

    \I__11114\ : LocalMux
    port map (
            O => \N__46971\,
            I => \N__46950\
        );

    \I__11113\ : LocalMux
    port map (
            O => \N__46968\,
            I => \N__46947\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__46965\,
            I => \N__46897\
        );

    \I__11111\ : LocalMux
    port map (
            O => \N__46962\,
            I => \N__46878\
        );

    \I__11110\ : LocalMux
    port map (
            O => \N__46959\,
            I => \N__46869\
        );

    \I__11109\ : LocalMux
    port map (
            O => \N__46956\,
            I => \N__46837\
        );

    \I__11108\ : Glb2LocalMux
    port map (
            O => \N__46953\,
            I => \N__46521\
        );

    \I__11107\ : Glb2LocalMux
    port map (
            O => \N__46950\,
            I => \N__46521\
        );

    \I__11106\ : Glb2LocalMux
    port map (
            O => \N__46947\,
            I => \N__46521\
        );

    \I__11105\ : SRMux
    port map (
            O => \N__46946\,
            I => \N__46521\
        );

    \I__11104\ : SRMux
    port map (
            O => \N__46945\,
            I => \N__46521\
        );

    \I__11103\ : SRMux
    port map (
            O => \N__46944\,
            I => \N__46521\
        );

    \I__11102\ : SRMux
    port map (
            O => \N__46943\,
            I => \N__46521\
        );

    \I__11101\ : SRMux
    port map (
            O => \N__46942\,
            I => \N__46521\
        );

    \I__11100\ : SRMux
    port map (
            O => \N__46941\,
            I => \N__46521\
        );

    \I__11099\ : SRMux
    port map (
            O => \N__46940\,
            I => \N__46521\
        );

    \I__11098\ : SRMux
    port map (
            O => \N__46939\,
            I => \N__46521\
        );

    \I__11097\ : SRMux
    port map (
            O => \N__46938\,
            I => \N__46521\
        );

    \I__11096\ : SRMux
    port map (
            O => \N__46937\,
            I => \N__46521\
        );

    \I__11095\ : SRMux
    port map (
            O => \N__46936\,
            I => \N__46521\
        );

    \I__11094\ : SRMux
    port map (
            O => \N__46935\,
            I => \N__46521\
        );

    \I__11093\ : SRMux
    port map (
            O => \N__46934\,
            I => \N__46521\
        );

    \I__11092\ : SRMux
    port map (
            O => \N__46933\,
            I => \N__46521\
        );

    \I__11091\ : SRMux
    port map (
            O => \N__46932\,
            I => \N__46521\
        );

    \I__11090\ : SRMux
    port map (
            O => \N__46931\,
            I => \N__46521\
        );

    \I__11089\ : SRMux
    port map (
            O => \N__46930\,
            I => \N__46521\
        );

    \I__11088\ : SRMux
    port map (
            O => \N__46929\,
            I => \N__46521\
        );

    \I__11087\ : SRMux
    port map (
            O => \N__46928\,
            I => \N__46521\
        );

    \I__11086\ : SRMux
    port map (
            O => \N__46927\,
            I => \N__46521\
        );

    \I__11085\ : SRMux
    port map (
            O => \N__46926\,
            I => \N__46521\
        );

    \I__11084\ : SRMux
    port map (
            O => \N__46925\,
            I => \N__46521\
        );

    \I__11083\ : SRMux
    port map (
            O => \N__46924\,
            I => \N__46521\
        );

    \I__11082\ : SRMux
    port map (
            O => \N__46923\,
            I => \N__46521\
        );

    \I__11081\ : SRMux
    port map (
            O => \N__46922\,
            I => \N__46521\
        );

    \I__11080\ : SRMux
    port map (
            O => \N__46921\,
            I => \N__46521\
        );

    \I__11079\ : SRMux
    port map (
            O => \N__46920\,
            I => \N__46521\
        );

    \I__11078\ : SRMux
    port map (
            O => \N__46919\,
            I => \N__46521\
        );

    \I__11077\ : SRMux
    port map (
            O => \N__46918\,
            I => \N__46521\
        );

    \I__11076\ : SRMux
    port map (
            O => \N__46917\,
            I => \N__46521\
        );

    \I__11075\ : SRMux
    port map (
            O => \N__46916\,
            I => \N__46521\
        );

    \I__11074\ : SRMux
    port map (
            O => \N__46915\,
            I => \N__46521\
        );

    \I__11073\ : SRMux
    port map (
            O => \N__46914\,
            I => \N__46521\
        );

    \I__11072\ : SRMux
    port map (
            O => \N__46913\,
            I => \N__46521\
        );

    \I__11071\ : SRMux
    port map (
            O => \N__46912\,
            I => \N__46521\
        );

    \I__11070\ : SRMux
    port map (
            O => \N__46911\,
            I => \N__46521\
        );

    \I__11069\ : SRMux
    port map (
            O => \N__46910\,
            I => \N__46521\
        );

    \I__11068\ : SRMux
    port map (
            O => \N__46909\,
            I => \N__46521\
        );

    \I__11067\ : SRMux
    port map (
            O => \N__46908\,
            I => \N__46521\
        );

    \I__11066\ : SRMux
    port map (
            O => \N__46907\,
            I => \N__46521\
        );

    \I__11065\ : SRMux
    port map (
            O => \N__46906\,
            I => \N__46521\
        );

    \I__11064\ : SRMux
    port map (
            O => \N__46905\,
            I => \N__46521\
        );

    \I__11063\ : SRMux
    port map (
            O => \N__46904\,
            I => \N__46521\
        );

    \I__11062\ : SRMux
    port map (
            O => \N__46903\,
            I => \N__46521\
        );

    \I__11061\ : SRMux
    port map (
            O => \N__46902\,
            I => \N__46521\
        );

    \I__11060\ : SRMux
    port map (
            O => \N__46901\,
            I => \N__46521\
        );

    \I__11059\ : SRMux
    port map (
            O => \N__46900\,
            I => \N__46521\
        );

    \I__11058\ : Glb2LocalMux
    port map (
            O => \N__46897\,
            I => \N__46521\
        );

    \I__11057\ : SRMux
    port map (
            O => \N__46896\,
            I => \N__46521\
        );

    \I__11056\ : SRMux
    port map (
            O => \N__46895\,
            I => \N__46521\
        );

    \I__11055\ : SRMux
    port map (
            O => \N__46894\,
            I => \N__46521\
        );

    \I__11054\ : SRMux
    port map (
            O => \N__46893\,
            I => \N__46521\
        );

    \I__11053\ : SRMux
    port map (
            O => \N__46892\,
            I => \N__46521\
        );

    \I__11052\ : SRMux
    port map (
            O => \N__46891\,
            I => \N__46521\
        );

    \I__11051\ : SRMux
    port map (
            O => \N__46890\,
            I => \N__46521\
        );

    \I__11050\ : SRMux
    port map (
            O => \N__46889\,
            I => \N__46521\
        );

    \I__11049\ : SRMux
    port map (
            O => \N__46888\,
            I => \N__46521\
        );

    \I__11048\ : SRMux
    port map (
            O => \N__46887\,
            I => \N__46521\
        );

    \I__11047\ : SRMux
    port map (
            O => \N__46886\,
            I => \N__46521\
        );

    \I__11046\ : SRMux
    port map (
            O => \N__46885\,
            I => \N__46521\
        );

    \I__11045\ : SRMux
    port map (
            O => \N__46884\,
            I => \N__46521\
        );

    \I__11044\ : SRMux
    port map (
            O => \N__46883\,
            I => \N__46521\
        );

    \I__11043\ : SRMux
    port map (
            O => \N__46882\,
            I => \N__46521\
        );

    \I__11042\ : SRMux
    port map (
            O => \N__46881\,
            I => \N__46521\
        );

    \I__11041\ : Glb2LocalMux
    port map (
            O => \N__46878\,
            I => \N__46521\
        );

    \I__11040\ : SRMux
    port map (
            O => \N__46877\,
            I => \N__46521\
        );

    \I__11039\ : SRMux
    port map (
            O => \N__46876\,
            I => \N__46521\
        );

    \I__11038\ : SRMux
    port map (
            O => \N__46875\,
            I => \N__46521\
        );

    \I__11037\ : SRMux
    port map (
            O => \N__46874\,
            I => \N__46521\
        );

    \I__11036\ : SRMux
    port map (
            O => \N__46873\,
            I => \N__46521\
        );

    \I__11035\ : SRMux
    port map (
            O => \N__46872\,
            I => \N__46521\
        );

    \I__11034\ : Glb2LocalMux
    port map (
            O => \N__46869\,
            I => \N__46521\
        );

    \I__11033\ : SRMux
    port map (
            O => \N__46868\,
            I => \N__46521\
        );

    \I__11032\ : SRMux
    port map (
            O => \N__46867\,
            I => \N__46521\
        );

    \I__11031\ : SRMux
    port map (
            O => \N__46866\,
            I => \N__46521\
        );

    \I__11030\ : SRMux
    port map (
            O => \N__46865\,
            I => \N__46521\
        );

    \I__11029\ : SRMux
    port map (
            O => \N__46864\,
            I => \N__46521\
        );

    \I__11028\ : SRMux
    port map (
            O => \N__46863\,
            I => \N__46521\
        );

    \I__11027\ : SRMux
    port map (
            O => \N__46862\,
            I => \N__46521\
        );

    \I__11026\ : SRMux
    port map (
            O => \N__46861\,
            I => \N__46521\
        );

    \I__11025\ : SRMux
    port map (
            O => \N__46860\,
            I => \N__46521\
        );

    \I__11024\ : SRMux
    port map (
            O => \N__46859\,
            I => \N__46521\
        );

    \I__11023\ : SRMux
    port map (
            O => \N__46858\,
            I => \N__46521\
        );

    \I__11022\ : SRMux
    port map (
            O => \N__46857\,
            I => \N__46521\
        );

    \I__11021\ : SRMux
    port map (
            O => \N__46856\,
            I => \N__46521\
        );

    \I__11020\ : SRMux
    port map (
            O => \N__46855\,
            I => \N__46521\
        );

    \I__11019\ : SRMux
    port map (
            O => \N__46854\,
            I => \N__46521\
        );

    \I__11018\ : SRMux
    port map (
            O => \N__46853\,
            I => \N__46521\
        );

    \I__11017\ : SRMux
    port map (
            O => \N__46852\,
            I => \N__46521\
        );

    \I__11016\ : SRMux
    port map (
            O => \N__46851\,
            I => \N__46521\
        );

    \I__11015\ : SRMux
    port map (
            O => \N__46850\,
            I => \N__46521\
        );

    \I__11014\ : SRMux
    port map (
            O => \N__46849\,
            I => \N__46521\
        );

    \I__11013\ : SRMux
    port map (
            O => \N__46848\,
            I => \N__46521\
        );

    \I__11012\ : SRMux
    port map (
            O => \N__46847\,
            I => \N__46521\
        );

    \I__11011\ : SRMux
    port map (
            O => \N__46846\,
            I => \N__46521\
        );

    \I__11010\ : SRMux
    port map (
            O => \N__46845\,
            I => \N__46521\
        );

    \I__11009\ : SRMux
    port map (
            O => \N__46844\,
            I => \N__46521\
        );

    \I__11008\ : SRMux
    port map (
            O => \N__46843\,
            I => \N__46521\
        );

    \I__11007\ : SRMux
    port map (
            O => \N__46842\,
            I => \N__46521\
        );

    \I__11006\ : SRMux
    port map (
            O => \N__46841\,
            I => \N__46521\
        );

    \I__11005\ : SRMux
    port map (
            O => \N__46840\,
            I => \N__46521\
        );

    \I__11004\ : Glb2LocalMux
    port map (
            O => \N__46837\,
            I => \N__46521\
        );

    \I__11003\ : SRMux
    port map (
            O => \N__46836\,
            I => \N__46521\
        );

    \I__11002\ : SRMux
    port map (
            O => \N__46835\,
            I => \N__46521\
        );

    \I__11001\ : SRMux
    port map (
            O => \N__46834\,
            I => \N__46521\
        );

    \I__11000\ : SRMux
    port map (
            O => \N__46833\,
            I => \N__46521\
        );

    \I__10999\ : SRMux
    port map (
            O => \N__46832\,
            I => \N__46521\
        );

    \I__10998\ : SRMux
    port map (
            O => \N__46831\,
            I => \N__46521\
        );

    \I__10997\ : SRMux
    port map (
            O => \N__46830\,
            I => \N__46521\
        );

    \I__10996\ : SRMux
    port map (
            O => \N__46829\,
            I => \N__46521\
        );

    \I__10995\ : SRMux
    port map (
            O => \N__46828\,
            I => \N__46521\
        );

    \I__10994\ : SRMux
    port map (
            O => \N__46827\,
            I => \N__46521\
        );

    \I__10993\ : SRMux
    port map (
            O => \N__46826\,
            I => \N__46521\
        );

    \I__10992\ : SRMux
    port map (
            O => \N__46825\,
            I => \N__46521\
        );

    \I__10991\ : SRMux
    port map (
            O => \N__46824\,
            I => \N__46521\
        );

    \I__10990\ : SRMux
    port map (
            O => \N__46823\,
            I => \N__46521\
        );

    \I__10989\ : SRMux
    port map (
            O => \N__46822\,
            I => \N__46521\
        );

    \I__10988\ : SRMux
    port map (
            O => \N__46821\,
            I => \N__46521\
        );

    \I__10987\ : SRMux
    port map (
            O => \N__46820\,
            I => \N__46521\
        );

    \I__10986\ : SRMux
    port map (
            O => \N__46819\,
            I => \N__46521\
        );

    \I__10985\ : SRMux
    port map (
            O => \N__46818\,
            I => \N__46521\
        );

    \I__10984\ : SRMux
    port map (
            O => \N__46817\,
            I => \N__46521\
        );

    \I__10983\ : SRMux
    port map (
            O => \N__46816\,
            I => \N__46521\
        );

    \I__10982\ : SRMux
    port map (
            O => \N__46815\,
            I => \N__46521\
        );

    \I__10981\ : SRMux
    port map (
            O => \N__46814\,
            I => \N__46521\
        );

    \I__10980\ : SRMux
    port map (
            O => \N__46813\,
            I => \N__46521\
        );

    \I__10979\ : SRMux
    port map (
            O => \N__46812\,
            I => \N__46521\
        );

    \I__10978\ : SRMux
    port map (
            O => \N__46811\,
            I => \N__46521\
        );

    \I__10977\ : SRMux
    port map (
            O => \N__46810\,
            I => \N__46521\
        );

    \I__10976\ : SRMux
    port map (
            O => \N__46809\,
            I => \N__46521\
        );

    \I__10975\ : SRMux
    port map (
            O => \N__46808\,
            I => \N__46521\
        );

    \I__10974\ : SRMux
    port map (
            O => \N__46807\,
            I => \N__46521\
        );

    \I__10973\ : SRMux
    port map (
            O => \N__46806\,
            I => \N__46521\
        );

    \I__10972\ : SRMux
    port map (
            O => \N__46805\,
            I => \N__46521\
        );

    \I__10971\ : SRMux
    port map (
            O => \N__46804\,
            I => \N__46521\
        );

    \I__10970\ : SRMux
    port map (
            O => \N__46803\,
            I => \N__46521\
        );

    \I__10969\ : SRMux
    port map (
            O => \N__46802\,
            I => \N__46521\
        );

    \I__10968\ : GlobalMux
    port map (
            O => \N__46521\,
            I => \N__46518\
        );

    \I__10967\ : gio2CtrlBuf
    port map (
            O => \N__46518\,
            I => red_c_g
        );

    \I__10966\ : InMux
    port map (
            O => \N__46515\,
            I => \N__46511\
        );

    \I__10965\ : InMux
    port map (
            O => \N__46514\,
            I => \N__46507\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__46511\,
            I => \N__46503\
        );

    \I__10963\ : InMux
    port map (
            O => \N__46510\,
            I => \N__46500\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__46507\,
            I => \N__46497\
        );

    \I__10961\ : InMux
    port map (
            O => \N__46506\,
            I => \N__46494\
        );

    \I__10960\ : Span4Mux_v
    port map (
            O => \N__46503\,
            I => \N__46489\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__46500\,
            I => \N__46489\
        );

    \I__10958\ : Span4Mux_h
    port map (
            O => \N__46497\,
            I => \N__46484\
        );

    \I__10957\ : LocalMux
    port map (
            O => \N__46494\,
            I => \N__46484\
        );

    \I__10956\ : Span4Mux_h
    port map (
            O => \N__46489\,
            I => \N__46481\
        );

    \I__10955\ : Span4Mux_h
    port map (
            O => \N__46484\,
            I => \N__46478\
        );

    \I__10954\ : Odrv4
    port map (
            O => \N__46481\,
            I => measured_delay_tr_18
        );

    \I__10953\ : Odrv4
    port map (
            O => \N__46478\,
            I => measured_delay_tr_18
        );

    \I__10952\ : InMux
    port map (
            O => \N__46473\,
            I => \N__46467\
        );

    \I__10951\ : InMux
    port map (
            O => \N__46472\,
            I => \N__46464\
        );

    \I__10950\ : InMux
    port map (
            O => \N__46471\,
            I => \N__46461\
        );

    \I__10949\ : InMux
    port map (
            O => \N__46470\,
            I => \N__46458\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__46467\,
            I => \N__46455\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__46464\,
            I => \N__46452\
        );

    \I__10946\ : LocalMux
    port map (
            O => \N__46461\,
            I => \N__46447\
        );

    \I__10945\ : LocalMux
    port map (
            O => \N__46458\,
            I => \N__46447\
        );

    \I__10944\ : Span4Mux_v
    port map (
            O => \N__46455\,
            I => \N__46440\
        );

    \I__10943\ : Span4Mux_v
    port map (
            O => \N__46452\,
            I => \N__46440\
        );

    \I__10942\ : Span4Mux_h
    port map (
            O => \N__46447\,
            I => \N__46440\
        );

    \I__10941\ : Span4Mux_h
    port map (
            O => \N__46440\,
            I => \N__46437\
        );

    \I__10940\ : Odrv4
    port map (
            O => \N__46437\,
            I => measured_delay_tr_17
        );

    \I__10939\ : CascadeMux
    port map (
            O => \N__46434\,
            I => \N__46429\
        );

    \I__10938\ : InMux
    port map (
            O => \N__46433\,
            I => \N__46426\
        );

    \I__10937\ : CascadeMux
    port map (
            O => \N__46432\,
            I => \N__46423\
        );

    \I__10936\ : InMux
    port map (
            O => \N__46429\,
            I => \N__46419\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__46426\,
            I => \N__46416\
        );

    \I__10934\ : InMux
    port map (
            O => \N__46423\,
            I => \N__46413\
        );

    \I__10933\ : InMux
    port map (
            O => \N__46422\,
            I => \N__46410\
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__46419\,
            I => \N__46407\
        );

    \I__10931\ : Span4Mux_v
    port map (
            O => \N__46416\,
            I => \N__46402\
        );

    \I__10930\ : LocalMux
    port map (
            O => \N__46413\,
            I => \N__46402\
        );

    \I__10929\ : LocalMux
    port map (
            O => \N__46410\,
            I => \N__46397\
        );

    \I__10928\ : Span4Mux_v
    port map (
            O => \N__46407\,
            I => \N__46397\
        );

    \I__10927\ : Span4Mux_v
    port map (
            O => \N__46402\,
            I => \N__46394\
        );

    \I__10926\ : Span4Mux_h
    port map (
            O => \N__46397\,
            I => \N__46391\
        );

    \I__10925\ : Span4Mux_h
    port map (
            O => \N__46394\,
            I => \N__46388\
        );

    \I__10924\ : Odrv4
    port map (
            O => \N__46391\,
            I => measured_delay_tr_19
        );

    \I__10923\ : Odrv4
    port map (
            O => \N__46388\,
            I => measured_delay_tr_19
        );

    \I__10922\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46377\
        );

    \I__10921\ : InMux
    port map (
            O => \N__46382\,
            I => \N__46374\
        );

    \I__10920\ : InMux
    port map (
            O => \N__46381\,
            I => \N__46371\
        );

    \I__10919\ : InMux
    port map (
            O => \N__46380\,
            I => \N__46368\
        );

    \I__10918\ : LocalMux
    port map (
            O => \N__46377\,
            I => \N__46365\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__46374\,
            I => \N__46362\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__46371\,
            I => \N__46357\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__46368\,
            I => \N__46357\
        );

    \I__10914\ : Span4Mux_v
    port map (
            O => \N__46365\,
            I => \N__46350\
        );

    \I__10913\ : Span4Mux_v
    port map (
            O => \N__46362\,
            I => \N__46350\
        );

    \I__10912\ : Span4Mux_h
    port map (
            O => \N__46357\,
            I => \N__46350\
        );

    \I__10911\ : Span4Mux_h
    port map (
            O => \N__46350\,
            I => \N__46347\
        );

    \I__10910\ : Odrv4
    port map (
            O => \N__46347\,
            I => measured_delay_tr_16
        );

    \I__10909\ : CascadeMux
    port map (
            O => \N__46344\,
            I => \N__46341\
        );

    \I__10908\ : InMux
    port map (
            O => \N__46341\,
            I => \N__46337\
        );

    \I__10907\ : InMux
    port map (
            O => \N__46340\,
            I => \N__46333\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__46337\,
            I => \N__46330\
        );

    \I__10905\ : CascadeMux
    port map (
            O => \N__46336\,
            I => \N__46327\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__46333\,
            I => \N__46324\
        );

    \I__10903\ : Span4Mux_h
    port map (
            O => \N__46330\,
            I => \N__46321\
        );

    \I__10902\ : InMux
    port map (
            O => \N__46327\,
            I => \N__46318\
        );

    \I__10901\ : Span4Mux_v
    port map (
            O => \N__46324\,
            I => \N__46315\
        );

    \I__10900\ : Odrv4
    port map (
            O => \N__46321\,
            I => measured_delay_tr_5
        );

    \I__10899\ : LocalMux
    port map (
            O => \N__46318\,
            I => measured_delay_tr_5
        );

    \I__10898\ : Odrv4
    port map (
            O => \N__46315\,
            I => measured_delay_tr_5
        );

    \I__10897\ : InMux
    port map (
            O => \N__46308\,
            I => \N__46303\
        );

    \I__10896\ : CascadeMux
    port map (
            O => \N__46307\,
            I => \N__46300\
        );

    \I__10895\ : InMux
    port map (
            O => \N__46306\,
            I => \N__46297\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__46303\,
            I => \N__46294\
        );

    \I__10893\ : InMux
    port map (
            O => \N__46300\,
            I => \N__46291\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__46297\,
            I => \N__46288\
        );

    \I__10891\ : Span4Mux_h
    port map (
            O => \N__46294\,
            I => \N__46285\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__46291\,
            I => \N__46280\
        );

    \I__10889\ : Span4Mux_v
    port map (
            O => \N__46288\,
            I => \N__46280\
        );

    \I__10888\ : Odrv4
    port map (
            O => \N__46285\,
            I => measured_delay_tr_4
        );

    \I__10887\ : Odrv4
    port map (
            O => \N__46280\,
            I => measured_delay_tr_4
        );

    \I__10886\ : CascadeMux
    port map (
            O => \N__46275\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3_cascade_\
        );

    \I__10885\ : InMux
    port map (
            O => \N__46272\,
            I => \N__46268\
        );

    \I__10884\ : InMux
    port map (
            O => \N__46271\,
            I => \N__46265\
        );

    \I__10883\ : LocalMux
    port map (
            O => \N__46268\,
            I => \phase_controller_inst1.stoper_tr.N_21\
        );

    \I__10882\ : LocalMux
    port map (
            O => \N__46265\,
            I => \phase_controller_inst1.stoper_tr.N_21\
        );

    \I__10881\ : CascadeMux
    port map (
            O => \N__46260\,
            I => \N__46257\
        );

    \I__10880\ : InMux
    port map (
            O => \N__46257\,
            I => \N__46252\
        );

    \I__10879\ : InMux
    port map (
            O => \N__46256\,
            I => \N__46249\
        );

    \I__10878\ : InMux
    port map (
            O => \N__46255\,
            I => \N__46245\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__46252\,
            I => \N__46242\
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__46249\,
            I => \N__46239\
        );

    \I__10875\ : InMux
    port map (
            O => \N__46248\,
            I => \N__46236\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__46245\,
            I => \N__46233\
        );

    \I__10873\ : Span4Mux_h
    port map (
            O => \N__46242\,
            I => \N__46230\
        );

    \I__10872\ : Sp12to4
    port map (
            O => \N__46239\,
            I => \N__46225\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__46236\,
            I => \N__46225\
        );

    \I__10870\ : Span4Mux_v
    port map (
            O => \N__46233\,
            I => \N__46222\
        );

    \I__10869\ : Odrv4
    port map (
            O => \N__46230\,
            I => measured_delay_tr_9
        );

    \I__10868\ : Odrv12
    port map (
            O => \N__46225\,
            I => measured_delay_tr_9
        );

    \I__10867\ : Odrv4
    port map (
            O => \N__46222\,
            I => measured_delay_tr_9
        );

    \I__10866\ : InMux
    port map (
            O => \N__46215\,
            I => \N__46211\
        );

    \I__10865\ : InMux
    port map (
            O => \N__46214\,
            I => \N__46208\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__46211\,
            I => \N__46205\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__46208\,
            I => \N__46202\
        );

    \I__10862\ : Odrv12
    port map (
            O => \N__46205\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6\
        );

    \I__10861\ : Odrv4
    port map (
            O => \N__46202\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6\
        );

    \I__10860\ : CascadeMux
    port map (
            O => \N__46197\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3_cascade_\
        );

    \I__10859\ : InMux
    port map (
            O => \N__46194\,
            I => \N__46189\
        );

    \I__10858\ : InMux
    port map (
            O => \N__46193\,
            I => \N__46186\
        );

    \I__10857\ : InMux
    port map (
            O => \N__46192\,
            I => \N__46183\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__46189\,
            I => \N__46180\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__46186\,
            I => \N__46175\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__46183\,
            I => \N__46175\
        );

    \I__10853\ : Span4Mux_h
    port map (
            O => \N__46180\,
            I => \N__46171\
        );

    \I__10852\ : Span4Mux_h
    port map (
            O => \N__46175\,
            I => \N__46168\
        );

    \I__10851\ : InMux
    port map (
            O => \N__46174\,
            I => \N__46165\
        );

    \I__10850\ : Odrv4
    port map (
            O => \N__46171\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6\
        );

    \I__10849\ : Odrv4
    port map (
            O => \N__46168\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__46165\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6\
        );

    \I__10847\ : InMux
    port map (
            O => \N__46158\,
            I => \N__46148\
        );

    \I__10846\ : InMux
    port map (
            O => \N__46157\,
            I => \N__46148\
        );

    \I__10845\ : InMux
    port map (
            O => \N__46156\,
            I => \N__46148\
        );

    \I__10844\ : InMux
    port map (
            O => \N__46155\,
            I => \N__46143\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__46148\,
            I => \N__46140\
        );

    \I__10842\ : InMux
    port map (
            O => \N__46147\,
            I => \N__46135\
        );

    \I__10841\ : InMux
    port map (
            O => \N__46146\,
            I => \N__46135\
        );

    \I__10840\ : LocalMux
    port map (
            O => \N__46143\,
            I => \N__46132\
        );

    \I__10839\ : Span4Mux_v
    port map (
            O => \N__46140\,
            I => \N__46127\
        );

    \I__10838\ : LocalMux
    port map (
            O => \N__46135\,
            I => \N__46127\
        );

    \I__10837\ : Span4Mux_h
    port map (
            O => \N__46132\,
            I => \N__46124\
        );

    \I__10836\ : Span4Mux_h
    port map (
            O => \N__46127\,
            I => \N__46121\
        );

    \I__10835\ : Odrv4
    port map (
            O => \N__46124\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3\
        );

    \I__10834\ : Odrv4
    port map (
            O => \N__46121\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3\
        );

    \I__10833\ : InMux
    port map (
            O => \N__46116\,
            I => \N__46113\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__46113\,
            I => \N__46110\
        );

    \I__10831\ : Odrv4
    port map (
            O => \N__46110\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__10830\ : InMux
    port map (
            O => \N__46107\,
            I => \N__46104\
        );

    \I__10829\ : LocalMux
    port map (
            O => \N__46104\,
            I => \N__46101\
        );

    \I__10828\ : Odrv4
    port map (
            O => \N__46101\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__10827\ : InMux
    port map (
            O => \N__46098\,
            I => \N__46092\
        );

    \I__10826\ : InMux
    port map (
            O => \N__46097\,
            I => \N__46092\
        );

    \I__10825\ : LocalMux
    port map (
            O => \N__46092\,
            I => \N__46089\
        );

    \I__10824\ : Odrv12
    port map (
            O => \N__46089\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2\
        );

    \I__10823\ : CascadeMux
    port map (
            O => \N__46086\,
            I => \N__46083\
        );

    \I__10822\ : InMux
    port map (
            O => \N__46083\,
            I => \N__46080\
        );

    \I__10821\ : LocalMux
    port map (
            O => \N__46080\,
            I => \N__46077\
        );

    \I__10820\ : Odrv12
    port map (
            O => \N__46077\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\
        );

    \I__10819\ : InMux
    port map (
            O => \N__46074\,
            I => \N__46071\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__46071\,
            I => \N__46067\
        );

    \I__10817\ : InMux
    port map (
            O => \N__46070\,
            I => \N__46064\
        );

    \I__10816\ : Span4Mux_h
    port map (
            O => \N__46067\,
            I => \N__46059\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__46064\,
            I => \N__46059\
        );

    \I__10814\ : Odrv4
    port map (
            O => \N__46059\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__10813\ : InMux
    port map (
            O => \N__46056\,
            I => \N__46053\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__46053\,
            I => \N__46050\
        );

    \I__10811\ : Span4Mux_h
    port map (
            O => \N__46050\,
            I => \N__46047\
        );

    \I__10810\ : Odrv4
    port map (
            O => \N__46047\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\
        );

    \I__10809\ : InMux
    port map (
            O => \N__46044\,
            I => \N__46040\
        );

    \I__10808\ : InMux
    port map (
            O => \N__46043\,
            I => \N__46037\
        );

    \I__10807\ : LocalMux
    port map (
            O => \N__46040\,
            I => \N__46034\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__46037\,
            I => \N__46031\
        );

    \I__10805\ : Odrv12
    port map (
            O => \N__46034\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__10804\ : Odrv4
    port map (
            O => \N__46031\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__10803\ : InMux
    port map (
            O => \N__46026\,
            I => \N__46023\
        );

    \I__10802\ : LocalMux
    port map (
            O => \N__46023\,
            I => \N__46020\
        );

    \I__10801\ : Span4Mux_v
    port map (
            O => \N__46020\,
            I => \N__46017\
        );

    \I__10800\ : Odrv4
    port map (
            O => \N__46017\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\
        );

    \I__10799\ : InMux
    port map (
            O => \N__46014\,
            I => \N__46010\
        );

    \I__10798\ : InMux
    port map (
            O => \N__46013\,
            I => \N__46007\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__46010\,
            I => \N__46002\
        );

    \I__10796\ : LocalMux
    port map (
            O => \N__46007\,
            I => \N__46002\
        );

    \I__10795\ : Odrv4
    port map (
            O => \N__46002\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__10794\ : InMux
    port map (
            O => \N__45999\,
            I => \N__45996\
        );

    \I__10793\ : LocalMux
    port map (
            O => \N__45996\,
            I => \N__45991\
        );

    \I__10792\ : InMux
    port map (
            O => \N__45995\,
            I => \N__45988\
        );

    \I__10791\ : InMux
    port map (
            O => \N__45994\,
            I => \N__45984\
        );

    \I__10790\ : Span4Mux_v
    port map (
            O => \N__45991\,
            I => \N__45979\
        );

    \I__10789\ : LocalMux
    port map (
            O => \N__45988\,
            I => \N__45979\
        );

    \I__10788\ : InMux
    port map (
            O => \N__45987\,
            I => \N__45976\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__45984\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__10786\ : Odrv4
    port map (
            O => \N__45979\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__10785\ : LocalMux
    port map (
            O => \N__45976\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__10784\ : InMux
    port map (
            O => \N__45969\,
            I => \N__45963\
        );

    \I__10783\ : InMux
    port map (
            O => \N__45968\,
            I => \N__45963\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__45963\,
            I => \N__45960\
        );

    \I__10781\ : Span4Mux_h
    port map (
            O => \N__45960\,
            I => \N__45953\
        );

    \I__10780\ : InMux
    port map (
            O => \N__45959\,
            I => \N__45948\
        );

    \I__10779\ : InMux
    port map (
            O => \N__45958\,
            I => \N__45948\
        );

    \I__10778\ : InMux
    port map (
            O => \N__45957\,
            I => \N__45945\
        );

    \I__10777\ : InMux
    port map (
            O => \N__45956\,
            I => \N__45942\
        );

    \I__10776\ : Span4Mux_v
    port map (
            O => \N__45953\,
            I => \N__45937\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__45948\,
            I => \N__45937\
        );

    \I__10774\ : LocalMux
    port map (
            O => \N__45945\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10773\ : LocalMux
    port map (
            O => \N__45942\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10772\ : Odrv4
    port map (
            O => \N__45937\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10771\ : CascadeMux
    port map (
            O => \N__45930\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__10770\ : CascadeMux
    port map (
            O => \N__45927\,
            I => \N__45924\
        );

    \I__10769\ : InMux
    port map (
            O => \N__45924\,
            I => \N__45919\
        );

    \I__10768\ : InMux
    port map (
            O => \N__45923\,
            I => \N__45916\
        );

    \I__10767\ : InMux
    port map (
            O => \N__45922\,
            I => \N__45913\
        );

    \I__10766\ : LocalMux
    port map (
            O => \N__45919\,
            I => \N__45910\
        );

    \I__10765\ : LocalMux
    port map (
            O => \N__45916\,
            I => \N__45907\
        );

    \I__10764\ : LocalMux
    port map (
            O => \N__45913\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10763\ : Odrv12
    port map (
            O => \N__45910\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10762\ : Odrv4
    port map (
            O => \N__45907\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10761\ : InMux
    port map (
            O => \N__45900\,
            I => \N__45897\
        );

    \I__10760\ : LocalMux
    port map (
            O => \N__45897\,
            I => \N__45894\
        );

    \I__10759\ : Odrv4
    port map (
            O => \N__45894\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\
        );

    \I__10758\ : InMux
    port map (
            O => \N__45891\,
            I => \N__45887\
        );

    \I__10757\ : InMux
    port map (
            O => \N__45890\,
            I => \N__45884\
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__45887\,
            I => \N__45881\
        );

    \I__10755\ : LocalMux
    port map (
            O => \N__45884\,
            I => \N__45878\
        );

    \I__10754\ : Odrv4
    port map (
            O => \N__45881\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__10753\ : Odrv4
    port map (
            O => \N__45878\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__10752\ : InMux
    port map (
            O => \N__45873\,
            I => \N__45870\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__45870\,
            I => \N__45867\
        );

    \I__10750\ : Odrv4
    port map (
            O => \N__45867\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\
        );

    \I__10749\ : InMux
    port map (
            O => \N__45864\,
            I => \N__45860\
        );

    \I__10748\ : InMux
    port map (
            O => \N__45863\,
            I => \N__45857\
        );

    \I__10747\ : LocalMux
    port map (
            O => \N__45860\,
            I => \N__45854\
        );

    \I__10746\ : LocalMux
    port map (
            O => \N__45857\,
            I => \N__45851\
        );

    \I__10745\ : Odrv12
    port map (
            O => \N__45854\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__10744\ : Odrv4
    port map (
            O => \N__45851\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__10743\ : CascadeMux
    port map (
            O => \N__45846\,
            I => \N__45843\
        );

    \I__10742\ : InMux
    port map (
            O => \N__45843\,
            I => \N__45840\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__45840\,
            I => \N__45837\
        );

    \I__10740\ : Odrv4
    port map (
            O => \N__45837\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\
        );

    \I__10739\ : InMux
    port map (
            O => \N__45834\,
            I => \N__45830\
        );

    \I__10738\ : InMux
    port map (
            O => \N__45833\,
            I => \N__45827\
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__45830\,
            I => \N__45822\
        );

    \I__10736\ : LocalMux
    port map (
            O => \N__45827\,
            I => \N__45822\
        );

    \I__10735\ : Odrv4
    port map (
            O => \N__45822\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__10734\ : InMux
    port map (
            O => \N__45819\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__10733\ : InMux
    port map (
            O => \N__45816\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__10732\ : InMux
    port map (
            O => \N__45813\,
            I => \N__45810\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__45810\,
            I => \N__45807\
        );

    \I__10730\ : Odrv4
    port map (
            O => \N__45807\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\
        );

    \I__10729\ : CascadeMux
    port map (
            O => \N__45804\,
            I => \N__45801\
        );

    \I__10728\ : InMux
    port map (
            O => \N__45801\,
            I => \N__45798\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__45798\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\
        );

    \I__10726\ : InMux
    port map (
            O => \N__45795\,
            I => \N__45791\
        );

    \I__10725\ : InMux
    port map (
            O => \N__45794\,
            I => \N__45788\
        );

    \I__10724\ : LocalMux
    port map (
            O => \N__45791\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__45788\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__10722\ : InMux
    port map (
            O => \N__45783\,
            I => \N__45780\
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__45780\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\
        );

    \I__10720\ : InMux
    port map (
            O => \N__45777\,
            I => \N__45773\
        );

    \I__10719\ : InMux
    port map (
            O => \N__45776\,
            I => \N__45770\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__45773\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__45770\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__10716\ : InMux
    port map (
            O => \N__45765\,
            I => \N__45762\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__45762\,
            I => \N__45759\
        );

    \I__10714\ : Span4Mux_v
    port map (
            O => \N__45759\,
            I => \N__45756\
        );

    \I__10713\ : Odrv4
    port map (
            O => \N__45756\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\
        );

    \I__10712\ : CascadeMux
    port map (
            O => \N__45753\,
            I => \N__45745\
        );

    \I__10711\ : CascadeMux
    port map (
            O => \N__45752\,
            I => \N__45742\
        );

    \I__10710\ : CascadeMux
    port map (
            O => \N__45751\,
            I => \N__45735\
        );

    \I__10709\ : CascadeMux
    port map (
            O => \N__45750\,
            I => \N__45727\
        );

    \I__10708\ : CascadeMux
    port map (
            O => \N__45749\,
            I => \N__45720\
        );

    \I__10707\ : CascadeMux
    port map (
            O => \N__45748\,
            I => \N__45717\
        );

    \I__10706\ : InMux
    port map (
            O => \N__45745\,
            I => \N__45710\
        );

    \I__10705\ : InMux
    port map (
            O => \N__45742\,
            I => \N__45710\
        );

    \I__10704\ : InMux
    port map (
            O => \N__45741\,
            I => \N__45701\
        );

    \I__10703\ : InMux
    port map (
            O => \N__45740\,
            I => \N__45701\
        );

    \I__10702\ : InMux
    port map (
            O => \N__45739\,
            I => \N__45701\
        );

    \I__10701\ : InMux
    port map (
            O => \N__45738\,
            I => \N__45701\
        );

    \I__10700\ : InMux
    port map (
            O => \N__45735\,
            I => \N__45698\
        );

    \I__10699\ : InMux
    port map (
            O => \N__45734\,
            I => \N__45691\
        );

    \I__10698\ : InMux
    port map (
            O => \N__45733\,
            I => \N__45691\
        );

    \I__10697\ : InMux
    port map (
            O => \N__45732\,
            I => \N__45691\
        );

    \I__10696\ : InMux
    port map (
            O => \N__45731\,
            I => \N__45688\
        );

    \I__10695\ : InMux
    port map (
            O => \N__45730\,
            I => \N__45685\
        );

    \I__10694\ : InMux
    port map (
            O => \N__45727\,
            I => \N__45682\
        );

    \I__10693\ : InMux
    port map (
            O => \N__45726\,
            I => \N__45675\
        );

    \I__10692\ : InMux
    port map (
            O => \N__45725\,
            I => \N__45675\
        );

    \I__10691\ : InMux
    port map (
            O => \N__45724\,
            I => \N__45675\
        );

    \I__10690\ : InMux
    port map (
            O => \N__45723\,
            I => \N__45670\
        );

    \I__10689\ : InMux
    port map (
            O => \N__45720\,
            I => \N__45661\
        );

    \I__10688\ : InMux
    port map (
            O => \N__45717\,
            I => \N__45661\
        );

    \I__10687\ : InMux
    port map (
            O => \N__45716\,
            I => \N__45661\
        );

    \I__10686\ : InMux
    port map (
            O => \N__45715\,
            I => \N__45661\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__45710\,
            I => \N__45651\
        );

    \I__10684\ : LocalMux
    port map (
            O => \N__45701\,
            I => \N__45651\
        );

    \I__10683\ : LocalMux
    port map (
            O => \N__45698\,
            I => \N__45651\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__45691\,
            I => \N__45651\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__45688\,
            I => \N__45648\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__45685\,
            I => \N__45641\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__45682\,
            I => \N__45641\
        );

    \I__10678\ : LocalMux
    port map (
            O => \N__45675\,
            I => \N__45641\
        );

    \I__10677\ : InMux
    port map (
            O => \N__45674\,
            I => \N__45636\
        );

    \I__10676\ : InMux
    port map (
            O => \N__45673\,
            I => \N__45636\
        );

    \I__10675\ : LocalMux
    port map (
            O => \N__45670\,
            I => \N__45633\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__45661\,
            I => \N__45630\
        );

    \I__10673\ : InMux
    port map (
            O => \N__45660\,
            I => \N__45627\
        );

    \I__10672\ : Span4Mux_v
    port map (
            O => \N__45651\,
            I => \N__45624\
        );

    \I__10671\ : Span12Mux_v
    port map (
            O => \N__45648\,
            I => \N__45621\
        );

    \I__10670\ : Span12Mux_h
    port map (
            O => \N__45641\,
            I => \N__45618\
        );

    \I__10669\ : LocalMux
    port map (
            O => \N__45636\,
            I => \N__45609\
        );

    \I__10668\ : Span4Mux_v
    port map (
            O => \N__45633\,
            I => \N__45609\
        );

    \I__10667\ : Span4Mux_h
    port map (
            O => \N__45630\,
            I => \N__45609\
        );

    \I__10666\ : LocalMux
    port map (
            O => \N__45627\,
            I => \N__45609\
        );

    \I__10665\ : Odrv4
    port map (
            O => \N__45624\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__10664\ : Odrv12
    port map (
            O => \N__45621\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__10663\ : Odrv12
    port map (
            O => \N__45618\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__10662\ : Odrv4
    port map (
            O => \N__45609\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__10661\ : CascadeMux
    port map (
            O => \N__45600\,
            I => \N__45593\
        );

    \I__10660\ : CascadeMux
    port map (
            O => \N__45599\,
            I => \N__45587\
        );

    \I__10659\ : CascadeMux
    port map (
            O => \N__45598\,
            I => \N__45584\
        );

    \I__10658\ : CascadeMux
    port map (
            O => \N__45597\,
            I => \N__45580\
        );

    \I__10657\ : CascadeMux
    port map (
            O => \N__45596\,
            I => \N__45577\
        );

    \I__10656\ : InMux
    port map (
            O => \N__45593\,
            I => \N__45570\
        );

    \I__10655\ : CascadeMux
    port map (
            O => \N__45592\,
            I => \N__45566\
        );

    \I__10654\ : CascadeMux
    port map (
            O => \N__45591\,
            I => \N__45562\
        );

    \I__10653\ : InMux
    port map (
            O => \N__45590\,
            I => \N__45553\
        );

    \I__10652\ : InMux
    port map (
            O => \N__45587\,
            I => \N__45553\
        );

    \I__10651\ : InMux
    port map (
            O => \N__45584\,
            I => \N__45544\
        );

    \I__10650\ : InMux
    port map (
            O => \N__45583\,
            I => \N__45544\
        );

    \I__10649\ : InMux
    port map (
            O => \N__45580\,
            I => \N__45544\
        );

    \I__10648\ : InMux
    port map (
            O => \N__45577\,
            I => \N__45544\
        );

    \I__10647\ : InMux
    port map (
            O => \N__45576\,
            I => \N__45535\
        );

    \I__10646\ : InMux
    port map (
            O => \N__45575\,
            I => \N__45535\
        );

    \I__10645\ : InMux
    port map (
            O => \N__45574\,
            I => \N__45535\
        );

    \I__10644\ : InMux
    port map (
            O => \N__45573\,
            I => \N__45535\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__45570\,
            I => \N__45530\
        );

    \I__10642\ : InMux
    port map (
            O => \N__45569\,
            I => \N__45521\
        );

    \I__10641\ : InMux
    port map (
            O => \N__45566\,
            I => \N__45521\
        );

    \I__10640\ : InMux
    port map (
            O => \N__45565\,
            I => \N__45521\
        );

    \I__10639\ : InMux
    port map (
            O => \N__45562\,
            I => \N__45521\
        );

    \I__10638\ : CascadeMux
    port map (
            O => \N__45561\,
            I => \N__45518\
        );

    \I__10637\ : CascadeMux
    port map (
            O => \N__45560\,
            I => \N__45514\
        );

    \I__10636\ : CascadeMux
    port map (
            O => \N__45559\,
            I => \N__45510\
        );

    \I__10635\ : CascadeMux
    port map (
            O => \N__45558\,
            I => \N__45507\
        );

    \I__10634\ : LocalMux
    port map (
            O => \N__45553\,
            I => \N__45504\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__45544\,
            I => \N__45499\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__45535\,
            I => \N__45499\
        );

    \I__10631\ : CascadeMux
    port map (
            O => \N__45534\,
            I => \N__45496\
        );

    \I__10630\ : InMux
    port map (
            O => \N__45533\,
            I => \N__45492\
        );

    \I__10629\ : Span4Mux_v
    port map (
            O => \N__45530\,
            I => \N__45489\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__45521\,
            I => \N__45486\
        );

    \I__10627\ : InMux
    port map (
            O => \N__45518\,
            I => \N__45473\
        );

    \I__10626\ : InMux
    port map (
            O => \N__45517\,
            I => \N__45473\
        );

    \I__10625\ : InMux
    port map (
            O => \N__45514\,
            I => \N__45473\
        );

    \I__10624\ : InMux
    port map (
            O => \N__45513\,
            I => \N__45473\
        );

    \I__10623\ : InMux
    port map (
            O => \N__45510\,
            I => \N__45473\
        );

    \I__10622\ : InMux
    port map (
            O => \N__45507\,
            I => \N__45473\
        );

    \I__10621\ : Span4Mux_v
    port map (
            O => \N__45504\,
            I => \N__45468\
        );

    \I__10620\ : Span4Mux_v
    port map (
            O => \N__45499\,
            I => \N__45468\
        );

    \I__10619\ : InMux
    port map (
            O => \N__45496\,
            I => \N__45463\
        );

    \I__10618\ : InMux
    port map (
            O => \N__45495\,
            I => \N__45463\
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__45492\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__10616\ : Odrv4
    port map (
            O => \N__45489\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__10615\ : Odrv4
    port map (
            O => \N__45486\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__45473\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__10613\ : Odrv4
    port map (
            O => \N__45468\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__45463\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__10611\ : InMux
    port map (
            O => \N__45450\,
            I => \N__45438\
        );

    \I__10610\ : InMux
    port map (
            O => \N__45449\,
            I => \N__45429\
        );

    \I__10609\ : InMux
    port map (
            O => \N__45448\,
            I => \N__45429\
        );

    \I__10608\ : InMux
    port map (
            O => \N__45447\,
            I => \N__45429\
        );

    \I__10607\ : InMux
    port map (
            O => \N__45446\,
            I => \N__45429\
        );

    \I__10606\ : InMux
    port map (
            O => \N__45445\,
            I => \N__45420\
        );

    \I__10605\ : InMux
    port map (
            O => \N__45444\,
            I => \N__45420\
        );

    \I__10604\ : InMux
    port map (
            O => \N__45443\,
            I => \N__45420\
        );

    \I__10603\ : InMux
    port map (
            O => \N__45442\,
            I => \N__45420\
        );

    \I__10602\ : CascadeMux
    port map (
            O => \N__45441\,
            I => \N__45408\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__45438\,
            I => \N__45402\
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__45429\,
            I => \N__45399\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__45420\,
            I => \N__45396\
        );

    \I__10598\ : InMux
    port map (
            O => \N__45419\,
            I => \N__45383\
        );

    \I__10597\ : InMux
    port map (
            O => \N__45418\,
            I => \N__45383\
        );

    \I__10596\ : InMux
    port map (
            O => \N__45417\,
            I => \N__45383\
        );

    \I__10595\ : InMux
    port map (
            O => \N__45416\,
            I => \N__45383\
        );

    \I__10594\ : InMux
    port map (
            O => \N__45415\,
            I => \N__45383\
        );

    \I__10593\ : InMux
    port map (
            O => \N__45414\,
            I => \N__45383\
        );

    \I__10592\ : CascadeMux
    port map (
            O => \N__45413\,
            I => \N__45380\
        );

    \I__10591\ : InMux
    port map (
            O => \N__45412\,
            I => \N__45374\
        );

    \I__10590\ : InMux
    port map (
            O => \N__45411\,
            I => \N__45374\
        );

    \I__10589\ : InMux
    port map (
            O => \N__45408\,
            I => \N__45371\
        );

    \I__10588\ : InMux
    port map (
            O => \N__45407\,
            I => \N__45364\
        );

    \I__10587\ : InMux
    port map (
            O => \N__45406\,
            I => \N__45364\
        );

    \I__10586\ : InMux
    port map (
            O => \N__45405\,
            I => \N__45364\
        );

    \I__10585\ : Span4Mux_v
    port map (
            O => \N__45402\,
            I => \N__45360\
        );

    \I__10584\ : Span4Mux_v
    port map (
            O => \N__45399\,
            I => \N__45353\
        );

    \I__10583\ : Span4Mux_v
    port map (
            O => \N__45396\,
            I => \N__45353\
        );

    \I__10582\ : LocalMux
    port map (
            O => \N__45383\,
            I => \N__45353\
        );

    \I__10581\ : InMux
    port map (
            O => \N__45380\,
            I => \N__45348\
        );

    \I__10580\ : InMux
    port map (
            O => \N__45379\,
            I => \N__45348\
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__45374\,
            I => \N__45345\
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__45371\,
            I => \N__45340\
        );

    \I__10577\ : LocalMux
    port map (
            O => \N__45364\,
            I => \N__45340\
        );

    \I__10576\ : InMux
    port map (
            O => \N__45363\,
            I => \N__45337\
        );

    \I__10575\ : Span4Mux_h
    port map (
            O => \N__45360\,
            I => \N__45334\
        );

    \I__10574\ : Span4Mux_h
    port map (
            O => \N__45353\,
            I => \N__45331\
        );

    \I__10573\ : LocalMux
    port map (
            O => \N__45348\,
            I => \N__45322\
        );

    \I__10572\ : Span4Mux_v
    port map (
            O => \N__45345\,
            I => \N__45322\
        );

    \I__10571\ : Span4Mux_h
    port map (
            O => \N__45340\,
            I => \N__45322\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__45337\,
            I => \N__45322\
        );

    \I__10569\ : Odrv4
    port map (
            O => \N__45334\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__10568\ : Odrv4
    port map (
            O => \N__45331\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__10567\ : Odrv4
    port map (
            O => \N__45322\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__10566\ : InMux
    port map (
            O => \N__45315\,
            I => \N__45311\
        );

    \I__10565\ : InMux
    port map (
            O => \N__45314\,
            I => \N__45308\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__45311\,
            I => \N__45305\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__45308\,
            I => \N__45302\
        );

    \I__10562\ : Span4Mux_h
    port map (
            O => \N__45305\,
            I => \N__45299\
        );

    \I__10561\ : Span4Mux_h
    port map (
            O => \N__45302\,
            I => \N__45296\
        );

    \I__10560\ : Odrv4
    port map (
            O => \N__45299\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__10559\ : Odrv4
    port map (
            O => \N__45296\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__10558\ : InMux
    port map (
            O => \N__45291\,
            I => \N__45288\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__45288\,
            I => \N__45285\
        );

    \I__10556\ : Odrv4
    port map (
            O => \N__45285\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\
        );

    \I__10555\ : CascadeMux
    port map (
            O => \N__45282\,
            I => \N__45279\
        );

    \I__10554\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45275\
        );

    \I__10553\ : InMux
    port map (
            O => \N__45278\,
            I => \N__45272\
        );

    \I__10552\ : LocalMux
    port map (
            O => \N__45275\,
            I => \N__45269\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__45272\,
            I => \N__45266\
        );

    \I__10550\ : Odrv12
    port map (
            O => \N__45269\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__10549\ : Odrv4
    port map (
            O => \N__45266\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__10548\ : CascadeMux
    port map (
            O => \N__45261\,
            I => \N__45258\
        );

    \I__10547\ : InMux
    port map (
            O => \N__45258\,
            I => \N__45255\
        );

    \I__10546\ : LocalMux
    port map (
            O => \N__45255\,
            I => \N__45252\
        );

    \I__10545\ : Odrv12
    port map (
            O => \N__45252\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\
        );

    \I__10544\ : InMux
    port map (
            O => \N__45249\,
            I => \N__45245\
        );

    \I__10543\ : InMux
    port map (
            O => \N__45248\,
            I => \N__45242\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__45245\,
            I => \N__45239\
        );

    \I__10541\ : LocalMux
    port map (
            O => \N__45242\,
            I => \N__45236\
        );

    \I__10540\ : Odrv12
    port map (
            O => \N__45239\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__10539\ : Odrv4
    port map (
            O => \N__45236\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__10538\ : InMux
    port map (
            O => \N__45231\,
            I => \N__45228\
        );

    \I__10537\ : LocalMux
    port map (
            O => \N__45228\,
            I => \N__45225\
        );

    \I__10536\ : Odrv4
    port map (
            O => \N__45225\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\
        );

    \I__10535\ : InMux
    port map (
            O => \N__45222\,
            I => \N__45218\
        );

    \I__10534\ : InMux
    port map (
            O => \N__45221\,
            I => \N__45215\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__45218\,
            I => \N__45210\
        );

    \I__10532\ : LocalMux
    port map (
            O => \N__45215\,
            I => \N__45210\
        );

    \I__10531\ : Odrv4
    port map (
            O => \N__45210\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__10530\ : InMux
    port map (
            O => \N__45207\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__10529\ : InMux
    port map (
            O => \N__45204\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__10528\ : InMux
    port map (
            O => \N__45201\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__10527\ : InMux
    port map (
            O => \N__45198\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__10526\ : InMux
    port map (
            O => \N__45195\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__10525\ : InMux
    port map (
            O => \N__45192\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__10524\ : InMux
    port map (
            O => \N__45189\,
            I => \N__45185\
        );

    \I__10523\ : InMux
    port map (
            O => \N__45188\,
            I => \N__45182\
        );

    \I__10522\ : LocalMux
    port map (
            O => \N__45185\,
            I => \N__45179\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__45182\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__10520\ : Odrv4
    port map (
            O => \N__45179\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__10519\ : InMux
    port map (
            O => \N__45174\,
            I => \N__45171\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__45171\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\
        );

    \I__10517\ : InMux
    port map (
            O => \N__45168\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__10516\ : InMux
    port map (
            O => \N__45165\,
            I => \N__45162\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__45162\,
            I => \N__45158\
        );

    \I__10514\ : InMux
    port map (
            O => \N__45161\,
            I => \N__45155\
        );

    \I__10513\ : Span4Mux_h
    port map (
            O => \N__45158\,
            I => \N__45152\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__45155\,
            I => \N__45149\
        );

    \I__10511\ : Odrv4
    port map (
            O => \N__45152\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__10510\ : Odrv4
    port map (
            O => \N__45149\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__10509\ : InMux
    port map (
            O => \N__45144\,
            I => \N__45141\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__45141\,
            I => \N__45138\
        );

    \I__10507\ : Odrv4
    port map (
            O => \N__45138\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\
        );

    \I__10506\ : InMux
    port map (
            O => \N__45135\,
            I => \bfn_18_16_0_\
        );

    \I__10505\ : InMux
    port map (
            O => \N__45132\,
            I => \N__45129\
        );

    \I__10504\ : LocalMux
    port map (
            O => \N__45129\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\
        );

    \I__10503\ : InMux
    port map (
            O => \N__45126\,
            I => \N__45123\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__45123\,
            I => \N__45120\
        );

    \I__10501\ : Span4Mux_h
    port map (
            O => \N__45120\,
            I => \N__45116\
        );

    \I__10500\ : InMux
    port map (
            O => \N__45119\,
            I => \N__45113\
        );

    \I__10499\ : Odrv4
    port map (
            O => \N__45116\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__10498\ : LocalMux
    port map (
            O => \N__45113\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__10497\ : InMux
    port map (
            O => \N__45108\,
            I => \N__45105\
        );

    \I__10496\ : LocalMux
    port map (
            O => \N__45105\,
            I => \N__45102\
        );

    \I__10495\ : Span4Mux_h
    port map (
            O => \N__45102\,
            I => \N__45099\
        );

    \I__10494\ : Odrv4
    port map (
            O => \N__45099\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\
        );

    \I__10493\ : InMux
    port map (
            O => \N__45096\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__10492\ : InMux
    port map (
            O => \N__45093\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__10491\ : InMux
    port map (
            O => \N__45090\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__10490\ : InMux
    port map (
            O => \N__45087\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__10489\ : InMux
    port map (
            O => \N__45084\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__10488\ : InMux
    port map (
            O => \N__45081\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__10487\ : InMux
    port map (
            O => \N__45078\,
            I => \N__45074\
        );

    \I__10486\ : InMux
    port map (
            O => \N__45077\,
            I => \N__45071\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__45074\,
            I => \N__45066\
        );

    \I__10484\ : LocalMux
    port map (
            O => \N__45071\,
            I => \N__45066\
        );

    \I__10483\ : Span4Mux_v
    port map (
            O => \N__45066\,
            I => \N__45063\
        );

    \I__10482\ : Odrv4
    port map (
            O => \N__45063\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__10481\ : InMux
    port map (
            O => \N__45060\,
            I => \N__45057\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__45057\,
            I => \N__45054\
        );

    \I__10479\ : Span4Mux_h
    port map (
            O => \N__45054\,
            I => \N__45051\
        );

    \I__10478\ : Odrv4
    port map (
            O => \N__45051\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\
        );

    \I__10477\ : InMux
    port map (
            O => \N__45048\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__10476\ : InMux
    port map (
            O => \N__45045\,
            I => \N__45041\
        );

    \I__10475\ : InMux
    port map (
            O => \N__45044\,
            I => \N__45038\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__45041\,
            I => \N__45035\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__45038\,
            I => \N__45032\
        );

    \I__10472\ : Span4Mux_v
    port map (
            O => \N__45035\,
            I => \N__45029\
        );

    \I__10471\ : Span4Mux_v
    port map (
            O => \N__45032\,
            I => \N__45026\
        );

    \I__10470\ : Odrv4
    port map (
            O => \N__45029\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__10469\ : Odrv4
    port map (
            O => \N__45026\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__10468\ : InMux
    port map (
            O => \N__45021\,
            I => \N__45018\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__45018\,
            I => \N__45015\
        );

    \I__10466\ : Span4Mux_h
    port map (
            O => \N__45015\,
            I => \N__45012\
        );

    \I__10465\ : Odrv4
    port map (
            O => \N__45012\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\
        );

    \I__10464\ : InMux
    port map (
            O => \N__45009\,
            I => \bfn_18_15_0_\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45006\,
            I => \N__45002\
        );

    \I__10462\ : InMux
    port map (
            O => \N__45005\,
            I => \N__44999\
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__45002\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__44999\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__10459\ : CascadeMux
    port map (
            O => \N__44994\,
            I => \N__44991\
        );

    \I__10458\ : InMux
    port map (
            O => \N__44991\,
            I => \N__44988\
        );

    \I__10457\ : LocalMux
    port map (
            O => \N__44988\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\
        );

    \I__10456\ : InMux
    port map (
            O => \N__44985\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__10455\ : InMux
    port map (
            O => \N__44982\,
            I => \N__44978\
        );

    \I__10454\ : InMux
    port map (
            O => \N__44981\,
            I => \N__44975\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__44978\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__44975\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10451\ : InMux
    port map (
            O => \N__44970\,
            I => \N__44967\
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__44967\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\
        );

    \I__10449\ : InMux
    port map (
            O => \N__44964\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__10448\ : InMux
    port map (
            O => \N__44961\,
            I => \N__44957\
        );

    \I__10447\ : InMux
    port map (
            O => \N__44960\,
            I => \N__44954\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__44957\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__44954\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10444\ : CascadeMux
    port map (
            O => \N__44949\,
            I => \N__44946\
        );

    \I__10443\ : InMux
    port map (
            O => \N__44946\,
            I => \N__44943\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__44943\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\
        );

    \I__10441\ : InMux
    port map (
            O => \N__44940\,
            I => \bfn_18_13_0_\
        );

    \I__10440\ : InMux
    port map (
            O => \N__44937\,
            I => \N__44933\
        );

    \I__10439\ : InMux
    port map (
            O => \N__44936\,
            I => \N__44930\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__44933\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__10437\ : LocalMux
    port map (
            O => \N__44930\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__10436\ : InMux
    port map (
            O => \N__44925\,
            I => \N__44922\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__44922\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\
        );

    \I__10434\ : InMux
    port map (
            O => \N__44919\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__10433\ : InMux
    port map (
            O => \N__44916\,
            I => \N__44912\
        );

    \I__10432\ : InMux
    port map (
            O => \N__44915\,
            I => \N__44909\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__44912\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__44909\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__10429\ : InMux
    port map (
            O => \N__44904\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__10428\ : CascadeMux
    port map (
            O => \N__44901\,
            I => \N__44898\
        );

    \I__10427\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44895\
        );

    \I__10426\ : LocalMux
    port map (
            O => \N__44895\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\
        );

    \I__10425\ : InMux
    port map (
            O => \N__44892\,
            I => \N__44868\
        );

    \I__10424\ : InMux
    port map (
            O => \N__44891\,
            I => \N__44868\
        );

    \I__10423\ : InMux
    port map (
            O => \N__44890\,
            I => \N__44851\
        );

    \I__10422\ : InMux
    port map (
            O => \N__44889\,
            I => \N__44851\
        );

    \I__10421\ : InMux
    port map (
            O => \N__44888\,
            I => \N__44851\
        );

    \I__10420\ : InMux
    port map (
            O => \N__44887\,
            I => \N__44851\
        );

    \I__10419\ : InMux
    port map (
            O => \N__44886\,
            I => \N__44851\
        );

    \I__10418\ : InMux
    port map (
            O => \N__44885\,
            I => \N__44851\
        );

    \I__10417\ : InMux
    port map (
            O => \N__44884\,
            I => \N__44851\
        );

    \I__10416\ : InMux
    port map (
            O => \N__44883\,
            I => \N__44851\
        );

    \I__10415\ : InMux
    port map (
            O => \N__44882\,
            I => \N__44834\
        );

    \I__10414\ : InMux
    port map (
            O => \N__44881\,
            I => \N__44834\
        );

    \I__10413\ : InMux
    port map (
            O => \N__44880\,
            I => \N__44834\
        );

    \I__10412\ : InMux
    port map (
            O => \N__44879\,
            I => \N__44834\
        );

    \I__10411\ : InMux
    port map (
            O => \N__44878\,
            I => \N__44834\
        );

    \I__10410\ : InMux
    port map (
            O => \N__44877\,
            I => \N__44834\
        );

    \I__10409\ : InMux
    port map (
            O => \N__44876\,
            I => \N__44834\
        );

    \I__10408\ : InMux
    port map (
            O => \N__44875\,
            I => \N__44834\
        );

    \I__10407\ : InMux
    port map (
            O => \N__44874\,
            I => \N__44831\
        );

    \I__10406\ : InMux
    port map (
            O => \N__44873\,
            I => \N__44828\
        );

    \I__10405\ : LocalMux
    port map (
            O => \N__44868\,
            I => \N__44823\
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__44851\,
            I => \N__44823\
        );

    \I__10403\ : LocalMux
    port map (
            O => \N__44834\,
            I => \N__44814\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__44831\,
            I => \N__44814\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__44828\,
            I => \N__44811\
        );

    \I__10400\ : Span4Mux_h
    port map (
            O => \N__44823\,
            I => \N__44808\
        );

    \I__10399\ : InMux
    port map (
            O => \N__44822\,
            I => \N__44805\
        );

    \I__10398\ : InMux
    port map (
            O => \N__44821\,
            I => \N__44802\
        );

    \I__10397\ : InMux
    port map (
            O => \N__44820\,
            I => \N__44797\
        );

    \I__10396\ : InMux
    port map (
            O => \N__44819\,
            I => \N__44797\
        );

    \I__10395\ : Span4Mux_h
    port map (
            O => \N__44814\,
            I => \N__44794\
        );

    \I__10394\ : Span4Mux_v
    port map (
            O => \N__44811\,
            I => \N__44787\
        );

    \I__10393\ : Span4Mux_h
    port map (
            O => \N__44808\,
            I => \N__44787\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__44805\,
            I => \N__44787\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__44802\,
            I => \N__44784\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__44797\,
            I => \N__44779\
        );

    \I__10389\ : Span4Mux_v
    port map (
            O => \N__44794\,
            I => \N__44779\
        );

    \I__10388\ : Odrv4
    port map (
            O => \N__44787\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__10387\ : Odrv12
    port map (
            O => \N__44784\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__10386\ : Odrv4
    port map (
            O => \N__44779\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__10385\ : CascadeMux
    port map (
            O => \N__44772\,
            I => \N__44760\
        );

    \I__10384\ : InMux
    port map (
            O => \N__44771\,
            I => \N__44733\
        );

    \I__10383\ : InMux
    port map (
            O => \N__44770\,
            I => \N__44733\
        );

    \I__10382\ : InMux
    port map (
            O => \N__44769\,
            I => \N__44733\
        );

    \I__10381\ : InMux
    port map (
            O => \N__44768\,
            I => \N__44733\
        );

    \I__10380\ : InMux
    port map (
            O => \N__44767\,
            I => \N__44733\
        );

    \I__10379\ : InMux
    port map (
            O => \N__44766\,
            I => \N__44733\
        );

    \I__10378\ : InMux
    port map (
            O => \N__44765\,
            I => \N__44733\
        );

    \I__10377\ : InMux
    port map (
            O => \N__44764\,
            I => \N__44733\
        );

    \I__10376\ : InMux
    port map (
            O => \N__44763\,
            I => \N__44730\
        );

    \I__10375\ : InMux
    port map (
            O => \N__44760\,
            I => \N__44726\
        );

    \I__10374\ : InMux
    port map (
            O => \N__44759\,
            I => \N__44709\
        );

    \I__10373\ : InMux
    port map (
            O => \N__44758\,
            I => \N__44709\
        );

    \I__10372\ : InMux
    port map (
            O => \N__44757\,
            I => \N__44709\
        );

    \I__10371\ : InMux
    port map (
            O => \N__44756\,
            I => \N__44709\
        );

    \I__10370\ : InMux
    port map (
            O => \N__44755\,
            I => \N__44709\
        );

    \I__10369\ : InMux
    port map (
            O => \N__44754\,
            I => \N__44709\
        );

    \I__10368\ : InMux
    port map (
            O => \N__44753\,
            I => \N__44709\
        );

    \I__10367\ : InMux
    port map (
            O => \N__44752\,
            I => \N__44709\
        );

    \I__10366\ : InMux
    port map (
            O => \N__44751\,
            I => \N__44702\
        );

    \I__10365\ : InMux
    port map (
            O => \N__44750\,
            I => \N__44702\
        );

    \I__10364\ : LocalMux
    port map (
            O => \N__44733\,
            I => \N__44697\
        );

    \I__10363\ : LocalMux
    port map (
            O => \N__44730\,
            I => \N__44697\
        );

    \I__10362\ : CascadeMux
    port map (
            O => \N__44729\,
            I => \N__44693\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__44726\,
            I => \N__44690\
        );

    \I__10360\ : LocalMux
    port map (
            O => \N__44709\,
            I => \N__44687\
        );

    \I__10359\ : InMux
    port map (
            O => \N__44708\,
            I => \N__44684\
        );

    \I__10358\ : InMux
    port map (
            O => \N__44707\,
            I => \N__44681\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__44702\,
            I => \N__44676\
        );

    \I__10356\ : Span4Mux_h
    port map (
            O => \N__44697\,
            I => \N__44676\
        );

    \I__10355\ : InMux
    port map (
            O => \N__44696\,
            I => \N__44671\
        );

    \I__10354\ : InMux
    port map (
            O => \N__44693\,
            I => \N__44671\
        );

    \I__10353\ : Span4Mux_v
    port map (
            O => \N__44690\,
            I => \N__44664\
        );

    \I__10352\ : Span4Mux_h
    port map (
            O => \N__44687\,
            I => \N__44664\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__44684\,
            I => \N__44664\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__44681\,
            I => \N__44661\
        );

    \I__10349\ : Span4Mux_v
    port map (
            O => \N__44676\,
            I => \N__44658\
        );

    \I__10348\ : LocalMux
    port map (
            O => \N__44671\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10347\ : Odrv4
    port map (
            O => \N__44664\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10346\ : Odrv12
    port map (
            O => \N__44661\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10345\ : Odrv4
    port map (
            O => \N__44658\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10344\ : InMux
    port map (
            O => \N__44649\,
            I => \N__44644\
        );

    \I__10343\ : InMux
    port map (
            O => \N__44648\,
            I => \N__44638\
        );

    \I__10342\ : InMux
    port map (
            O => \N__44647\,
            I => \N__44638\
        );

    \I__10341\ : LocalMux
    port map (
            O => \N__44644\,
            I => \N__44635\
        );

    \I__10340\ : InMux
    port map (
            O => \N__44643\,
            I => \N__44632\
        );

    \I__10339\ : LocalMux
    port map (
            O => \N__44638\,
            I => \N__44629\
        );

    \I__10338\ : Odrv12
    port map (
            O => \N__44635\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__44632\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__10336\ : Odrv4
    port map (
            O => \N__44629\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__10335\ : InMux
    port map (
            O => \N__44622\,
            I => \N__44615\
        );

    \I__10334\ : InMux
    port map (
            O => \N__44621\,
            I => \N__44615\
        );

    \I__10333\ : InMux
    port map (
            O => \N__44620\,
            I => \N__44612\
        );

    \I__10332\ : LocalMux
    port map (
            O => \N__44615\,
            I => \N__44608\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__44612\,
            I => \N__44604\
        );

    \I__10330\ : InMux
    port map (
            O => \N__44611\,
            I => \N__44601\
        );

    \I__10329\ : Span4Mux_h
    port map (
            O => \N__44608\,
            I => \N__44598\
        );

    \I__10328\ : InMux
    port map (
            O => \N__44607\,
            I => \N__44595\
        );

    \I__10327\ : Span4Mux_h
    port map (
            O => \N__44604\,
            I => \N__44590\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__44601\,
            I => \N__44590\
        );

    \I__10325\ : Odrv4
    port map (
            O => \N__44598\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__44595\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10323\ : Odrv4
    port map (
            O => \N__44590\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10322\ : InMux
    port map (
            O => \N__44583\,
            I => \N__44580\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__44580\,
            I => \N__44577\
        );

    \I__10320\ : Odrv4
    port map (
            O => \N__44577\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\
        );

    \I__10319\ : InMux
    port map (
            O => \N__44574\,
            I => \N__44570\
        );

    \I__10318\ : InMux
    port map (
            O => \N__44573\,
            I => \N__44567\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__44570\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__44567\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__10315\ : CascadeMux
    port map (
            O => \N__44562\,
            I => \N__44559\
        );

    \I__10314\ : InMux
    port map (
            O => \N__44559\,
            I => \N__44556\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__44556\,
            I => \N__44553\
        );

    \I__10312\ : Odrv4
    port map (
            O => \N__44553\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\
        );

    \I__10311\ : InMux
    port map (
            O => \N__44550\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__10310\ : InMux
    port map (
            O => \N__44547\,
            I => \N__44543\
        );

    \I__10309\ : InMux
    port map (
            O => \N__44546\,
            I => \N__44540\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__44543\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__44540\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__10306\ : InMux
    port map (
            O => \N__44535\,
            I => \N__44532\
        );

    \I__10305\ : LocalMux
    port map (
            O => \N__44532\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\
        );

    \I__10304\ : InMux
    port map (
            O => \N__44529\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__10303\ : InMux
    port map (
            O => \N__44526\,
            I => \N__44522\
        );

    \I__10302\ : InMux
    port map (
            O => \N__44525\,
            I => \N__44519\
        );

    \I__10301\ : LocalMux
    port map (
            O => \N__44522\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__44519\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__10299\ : InMux
    port map (
            O => \N__44514\,
            I => \N__44511\
        );

    \I__10298\ : LocalMux
    port map (
            O => \N__44511\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\
        );

    \I__10297\ : InMux
    port map (
            O => \N__44508\,
            I => \bfn_18_12_0_\
        );

    \I__10296\ : InMux
    port map (
            O => \N__44505\,
            I => \N__44501\
        );

    \I__10295\ : InMux
    port map (
            O => \N__44504\,
            I => \N__44498\
        );

    \I__10294\ : LocalMux
    port map (
            O => \N__44501\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__44498\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__10292\ : InMux
    port map (
            O => \N__44493\,
            I => \N__44490\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__44490\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\
        );

    \I__10290\ : InMux
    port map (
            O => \N__44487\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__10289\ : InMux
    port map (
            O => \N__44484\,
            I => \N__44481\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__44481\,
            I => \N__44477\
        );

    \I__10287\ : InMux
    port map (
            O => \N__44480\,
            I => \N__44474\
        );

    \I__10286\ : Odrv12
    port map (
            O => \N__44477\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__44474\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__10284\ : CascadeMux
    port map (
            O => \N__44469\,
            I => \N__44466\
        );

    \I__10283\ : InMux
    port map (
            O => \N__44466\,
            I => \N__44463\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__44463\,
            I => \N__44460\
        );

    \I__10281\ : Odrv4
    port map (
            O => \N__44460\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\
        );

    \I__10280\ : InMux
    port map (
            O => \N__44457\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__10279\ : InMux
    port map (
            O => \N__44454\,
            I => \N__44450\
        );

    \I__10278\ : InMux
    port map (
            O => \N__44453\,
            I => \N__44447\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__44450\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__44447\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__10275\ : CascadeMux
    port map (
            O => \N__44442\,
            I => \N__44439\
        );

    \I__10274\ : InMux
    port map (
            O => \N__44439\,
            I => \N__44436\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__44436\,
            I => \N__44433\
        );

    \I__10272\ : Odrv4
    port map (
            O => \N__44433\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\
        );

    \I__10271\ : InMux
    port map (
            O => \N__44430\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__10270\ : InMux
    port map (
            O => \N__44427\,
            I => \N__44424\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__44424\,
            I => \N__44420\
        );

    \I__10268\ : InMux
    port map (
            O => \N__44423\,
            I => \N__44417\
        );

    \I__10267\ : Span4Mux_h
    port map (
            O => \N__44420\,
            I => \N__44412\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__44417\,
            I => \N__44412\
        );

    \I__10265\ : Span4Mux_h
    port map (
            O => \N__44412\,
            I => \N__44409\
        );

    \I__10264\ : Odrv4
    port map (
            O => \N__44409\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__10263\ : InMux
    port map (
            O => \N__44406\,
            I => \N__44403\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__44403\,
            I => \N__44400\
        );

    \I__10261\ : Span4Mux_v
    port map (
            O => \N__44400\,
            I => \N__44397\
        );

    \I__10260\ : Odrv4
    port map (
            O => \N__44397\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\
        );

    \I__10259\ : InMux
    port map (
            O => \N__44394\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__10258\ : InMux
    port map (
            O => \N__44391\,
            I => \N__44387\
        );

    \I__10257\ : InMux
    port map (
            O => \N__44390\,
            I => \N__44384\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__44387\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__10255\ : LocalMux
    port map (
            O => \N__44384\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__10254\ : CascadeMux
    port map (
            O => \N__44379\,
            I => \N__44376\
        );

    \I__10253\ : InMux
    port map (
            O => \N__44376\,
            I => \N__44373\
        );

    \I__10252\ : LocalMux
    port map (
            O => \N__44373\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\
        );

    \I__10251\ : InMux
    port map (
            O => \N__44370\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__10250\ : CascadeMux
    port map (
            O => \N__44367\,
            I => \N__44363\
        );

    \I__10249\ : InMux
    port map (
            O => \N__44366\,
            I => \N__44360\
        );

    \I__10248\ : InMux
    port map (
            O => \N__44363\,
            I => \N__44357\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__44360\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__44357\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__10245\ : InMux
    port map (
            O => \N__44352\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__10244\ : InMux
    port map (
            O => \N__44349\,
            I => \N__44311\
        );

    \I__10243\ : InMux
    port map (
            O => \N__44348\,
            I => \N__44311\
        );

    \I__10242\ : InMux
    port map (
            O => \N__44347\,
            I => \N__44311\
        );

    \I__10241\ : InMux
    port map (
            O => \N__44346\,
            I => \N__44311\
        );

    \I__10240\ : InMux
    port map (
            O => \N__44345\,
            I => \N__44302\
        );

    \I__10239\ : InMux
    port map (
            O => \N__44344\,
            I => \N__44302\
        );

    \I__10238\ : InMux
    port map (
            O => \N__44343\,
            I => \N__44302\
        );

    \I__10237\ : InMux
    port map (
            O => \N__44342\,
            I => \N__44302\
        );

    \I__10236\ : InMux
    port map (
            O => \N__44341\,
            I => \N__44293\
        );

    \I__10235\ : InMux
    port map (
            O => \N__44340\,
            I => \N__44293\
        );

    \I__10234\ : InMux
    port map (
            O => \N__44339\,
            I => \N__44293\
        );

    \I__10233\ : InMux
    port map (
            O => \N__44338\,
            I => \N__44293\
        );

    \I__10232\ : InMux
    port map (
            O => \N__44337\,
            I => \N__44284\
        );

    \I__10231\ : InMux
    port map (
            O => \N__44336\,
            I => \N__44284\
        );

    \I__10230\ : InMux
    port map (
            O => \N__44335\,
            I => \N__44284\
        );

    \I__10229\ : InMux
    port map (
            O => \N__44334\,
            I => \N__44284\
        );

    \I__10228\ : InMux
    port map (
            O => \N__44333\,
            I => \N__44275\
        );

    \I__10227\ : InMux
    port map (
            O => \N__44332\,
            I => \N__44275\
        );

    \I__10226\ : InMux
    port map (
            O => \N__44331\,
            I => \N__44275\
        );

    \I__10225\ : InMux
    port map (
            O => \N__44330\,
            I => \N__44275\
        );

    \I__10224\ : InMux
    port map (
            O => \N__44329\,
            I => \N__44270\
        );

    \I__10223\ : InMux
    port map (
            O => \N__44328\,
            I => \N__44270\
        );

    \I__10222\ : InMux
    port map (
            O => \N__44327\,
            I => \N__44261\
        );

    \I__10221\ : InMux
    port map (
            O => \N__44326\,
            I => \N__44261\
        );

    \I__10220\ : InMux
    port map (
            O => \N__44325\,
            I => \N__44261\
        );

    \I__10219\ : InMux
    port map (
            O => \N__44324\,
            I => \N__44261\
        );

    \I__10218\ : InMux
    port map (
            O => \N__44323\,
            I => \N__44252\
        );

    \I__10217\ : InMux
    port map (
            O => \N__44322\,
            I => \N__44252\
        );

    \I__10216\ : InMux
    port map (
            O => \N__44321\,
            I => \N__44252\
        );

    \I__10215\ : InMux
    port map (
            O => \N__44320\,
            I => \N__44252\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__44311\,
            I => \N__44243\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__44302\,
            I => \N__44243\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__44293\,
            I => \N__44243\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__44284\,
            I => \N__44243\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__44275\,
            I => \N__44236\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__44270\,
            I => \N__44236\
        );

    \I__10208\ : LocalMux
    port map (
            O => \N__44261\,
            I => \N__44236\
        );

    \I__10207\ : LocalMux
    port map (
            O => \N__44252\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__10206\ : Odrv4
    port map (
            O => \N__44243\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__10205\ : Odrv12
    port map (
            O => \N__44236\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__10204\ : InMux
    port map (
            O => \N__44229\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__10203\ : CascadeMux
    port map (
            O => \N__44226\,
            I => \N__44222\
        );

    \I__10202\ : InMux
    port map (
            O => \N__44225\,
            I => \N__44219\
        );

    \I__10201\ : InMux
    port map (
            O => \N__44222\,
            I => \N__44216\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__44219\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__10199\ : LocalMux
    port map (
            O => \N__44216\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__10198\ : CEMux
    port map (
            O => \N__44211\,
            I => \N__44208\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__44208\,
            I => \N__44202\
        );

    \I__10196\ : CEMux
    port map (
            O => \N__44207\,
            I => \N__44199\
        );

    \I__10195\ : CEMux
    port map (
            O => \N__44206\,
            I => \N__44196\
        );

    \I__10194\ : CEMux
    port map (
            O => \N__44205\,
            I => \N__44193\
        );

    \I__10193\ : Span4Mux_v
    port map (
            O => \N__44202\,
            I => \N__44188\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__44199\,
            I => \N__44188\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__44196\,
            I => \N__44183\
        );

    \I__10190\ : LocalMux
    port map (
            O => \N__44193\,
            I => \N__44183\
        );

    \I__10189\ : Span4Mux_v
    port map (
            O => \N__44188\,
            I => \N__44178\
        );

    \I__10188\ : Span4Mux_v
    port map (
            O => \N__44183\,
            I => \N__44178\
        );

    \I__10187\ : Odrv4
    port map (
            O => \N__44178\,
            I => \delay_measurement_inst.delay_hc_timer.N_336_i\
        );

    \I__10186\ : InMux
    port map (
            O => \N__44175\,
            I => \N__44172\
        );

    \I__10185\ : LocalMux
    port map (
            O => \N__44172\,
            I => \N__44169\
        );

    \I__10184\ : Span4Mux_h
    port map (
            O => \N__44169\,
            I => \N__44166\
        );

    \I__10183\ : Odrv4
    port map (
            O => \N__44166\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\
        );

    \I__10182\ : CascadeMux
    port map (
            O => \N__44163\,
            I => \N__44160\
        );

    \I__10181\ : InMux
    port map (
            O => \N__44160\,
            I => \N__44157\
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__44157\,
            I => \N__44153\
        );

    \I__10179\ : InMux
    port map (
            O => \N__44156\,
            I => \N__44149\
        );

    \I__10178\ : Span4Mux_h
    port map (
            O => \N__44153\,
            I => \N__44146\
        );

    \I__10177\ : InMux
    port map (
            O => \N__44152\,
            I => \N__44143\
        );

    \I__10176\ : LocalMux
    port map (
            O => \N__44149\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__10175\ : Odrv4
    port map (
            O => \N__44146\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__10174\ : LocalMux
    port map (
            O => \N__44143\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__10173\ : InMux
    port map (
            O => \N__44136\,
            I => \N__44132\
        );

    \I__10172\ : InMux
    port map (
            O => \N__44135\,
            I => \N__44129\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__44132\,
            I => \N__44126\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__44129\,
            I => \N__44123\
        );

    \I__10169\ : Odrv4
    port map (
            O => \N__44126\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__10168\ : Odrv4
    port map (
            O => \N__44123\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__10167\ : InMux
    port map (
            O => \N__44118\,
            I => \N__44115\
        );

    \I__10166\ : LocalMux
    port map (
            O => \N__44115\,
            I => \N__44112\
        );

    \I__10165\ : Span4Mux_h
    port map (
            O => \N__44112\,
            I => \N__44109\
        );

    \I__10164\ : Odrv4
    port map (
            O => \N__44109\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\
        );

    \I__10163\ : InMux
    port map (
            O => \N__44106\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__10162\ : CascadeMux
    port map (
            O => \N__44103\,
            I => \N__44100\
        );

    \I__10161\ : InMux
    port map (
            O => \N__44100\,
            I => \N__44096\
        );

    \I__10160\ : InMux
    port map (
            O => \N__44099\,
            I => \N__44093\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__44096\,
            I => \N__44090\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__44093\,
            I => \N__44087\
        );

    \I__10157\ : Odrv4
    port map (
            O => \N__44090\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__10156\ : Odrv4
    port map (
            O => \N__44087\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__10155\ : CascadeMux
    port map (
            O => \N__44082\,
            I => \N__44079\
        );

    \I__10154\ : InMux
    port map (
            O => \N__44079\,
            I => \N__44076\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__44076\,
            I => \N__44073\
        );

    \I__10152\ : Span4Mux_v
    port map (
            O => \N__44073\,
            I => \N__44070\
        );

    \I__10151\ : Odrv4
    port map (
            O => \N__44070\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\
        );

    \I__10150\ : InMux
    port map (
            O => \N__44067\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__10149\ : InMux
    port map (
            O => \N__44064\,
            I => \N__44060\
        );

    \I__10148\ : InMux
    port map (
            O => \N__44063\,
            I => \N__44057\
        );

    \I__10147\ : LocalMux
    port map (
            O => \N__44060\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__10146\ : LocalMux
    port map (
            O => \N__44057\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__10145\ : InMux
    port map (
            O => \N__44052\,
            I => \N__44049\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__44049\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\
        );

    \I__10143\ : InMux
    port map (
            O => \N__44046\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__10142\ : InMux
    port map (
            O => \N__44043\,
            I => \N__44039\
        );

    \I__10141\ : InMux
    port map (
            O => \N__44042\,
            I => \N__44036\
        );

    \I__10140\ : LocalMux
    port map (
            O => \N__44039\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__44036\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__10138\ : CascadeMux
    port map (
            O => \N__44031\,
            I => \N__44028\
        );

    \I__10137\ : InMux
    port map (
            O => \N__44028\,
            I => \N__44025\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__44025\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\
        );

    \I__10135\ : InMux
    port map (
            O => \N__44022\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__10134\ : InMux
    port map (
            O => \N__44019\,
            I => \N__44015\
        );

    \I__10133\ : InMux
    port map (
            O => \N__44018\,
            I => \N__44012\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__44015\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__44012\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__10130\ : InMux
    port map (
            O => \N__44007\,
            I => \N__44004\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__44004\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\
        );

    \I__10128\ : InMux
    port map (
            O => \N__44001\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__10127\ : CascadeMux
    port map (
            O => \N__43998\,
            I => \N__43993\
        );

    \I__10126\ : InMux
    port map (
            O => \N__43997\,
            I => \N__43990\
        );

    \I__10125\ : InMux
    port map (
            O => \N__43996\,
            I => \N__43987\
        );

    \I__10124\ : InMux
    port map (
            O => \N__43993\,
            I => \N__43984\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__43990\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__43987\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__43984\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__10120\ : InMux
    port map (
            O => \N__43977\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__10119\ : CascadeMux
    port map (
            O => \N__43974\,
            I => \N__43969\
        );

    \I__10118\ : InMux
    port map (
            O => \N__43973\,
            I => \N__43966\
        );

    \I__10117\ : InMux
    port map (
            O => \N__43972\,
            I => \N__43963\
        );

    \I__10116\ : InMux
    port map (
            O => \N__43969\,
            I => \N__43960\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__43966\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__10114\ : LocalMux
    port map (
            O => \N__43963\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__43960\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__10112\ : InMux
    port map (
            O => \N__43953\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__10111\ : CascadeMux
    port map (
            O => \N__43950\,
            I => \N__43945\
        );

    \I__10110\ : InMux
    port map (
            O => \N__43949\,
            I => \N__43942\
        );

    \I__10109\ : InMux
    port map (
            O => \N__43948\,
            I => \N__43939\
        );

    \I__10108\ : InMux
    port map (
            O => \N__43945\,
            I => \N__43936\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__43942\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__43939\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__10105\ : LocalMux
    port map (
            O => \N__43936\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__10104\ : InMux
    port map (
            O => \N__43929\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__10103\ : CascadeMux
    port map (
            O => \N__43926\,
            I => \N__43921\
        );

    \I__10102\ : InMux
    port map (
            O => \N__43925\,
            I => \N__43918\
        );

    \I__10101\ : InMux
    port map (
            O => \N__43924\,
            I => \N__43915\
        );

    \I__10100\ : InMux
    port map (
            O => \N__43921\,
            I => \N__43912\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__43918\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__43915\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__43912\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__10096\ : InMux
    port map (
            O => \N__43905\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__10095\ : CascadeMux
    port map (
            O => \N__43902\,
            I => \N__43897\
        );

    \I__10094\ : InMux
    port map (
            O => \N__43901\,
            I => \N__43894\
        );

    \I__10093\ : InMux
    port map (
            O => \N__43900\,
            I => \N__43891\
        );

    \I__10092\ : InMux
    port map (
            O => \N__43897\,
            I => \N__43888\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__43894\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__43891\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__43888\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__10088\ : InMux
    port map (
            O => \N__43881\,
            I => \bfn_18_10_0_\
        );

    \I__10087\ : CascadeMux
    port map (
            O => \N__43878\,
            I => \N__43873\
        );

    \I__10086\ : InMux
    port map (
            O => \N__43877\,
            I => \N__43870\
        );

    \I__10085\ : InMux
    port map (
            O => \N__43876\,
            I => \N__43867\
        );

    \I__10084\ : InMux
    port map (
            O => \N__43873\,
            I => \N__43864\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__43870\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__10082\ : LocalMux
    port map (
            O => \N__43867\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__43864\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__10080\ : InMux
    port map (
            O => \N__43857\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__10079\ : CascadeMux
    port map (
            O => \N__43854\,
            I => \N__43849\
        );

    \I__10078\ : InMux
    port map (
            O => \N__43853\,
            I => \N__43846\
        );

    \I__10077\ : InMux
    port map (
            O => \N__43852\,
            I => \N__43843\
        );

    \I__10076\ : InMux
    port map (
            O => \N__43849\,
            I => \N__43840\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__43846\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__43843\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__10073\ : LocalMux
    port map (
            O => \N__43840\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__10072\ : InMux
    port map (
            O => \N__43833\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__10071\ : CascadeMux
    port map (
            O => \N__43830\,
            I => \N__43825\
        );

    \I__10070\ : InMux
    port map (
            O => \N__43829\,
            I => \N__43822\
        );

    \I__10069\ : InMux
    port map (
            O => \N__43828\,
            I => \N__43819\
        );

    \I__10068\ : InMux
    port map (
            O => \N__43825\,
            I => \N__43816\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__43822\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__10066\ : LocalMux
    port map (
            O => \N__43819\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__43816\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__10064\ : InMux
    port map (
            O => \N__43809\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__10063\ : CascadeMux
    port map (
            O => \N__43806\,
            I => \N__43801\
        );

    \I__10062\ : InMux
    port map (
            O => \N__43805\,
            I => \N__43798\
        );

    \I__10061\ : InMux
    port map (
            O => \N__43804\,
            I => \N__43795\
        );

    \I__10060\ : InMux
    port map (
            O => \N__43801\,
            I => \N__43792\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__43798\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__43795\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__43792\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__10056\ : InMux
    port map (
            O => \N__43785\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__10055\ : CascadeMux
    port map (
            O => \N__43782\,
            I => \N__43777\
        );

    \I__10054\ : InMux
    port map (
            O => \N__43781\,
            I => \N__43774\
        );

    \I__10053\ : InMux
    port map (
            O => \N__43780\,
            I => \N__43771\
        );

    \I__10052\ : InMux
    port map (
            O => \N__43777\,
            I => \N__43768\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__43774\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__43771\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__43768\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__10048\ : InMux
    port map (
            O => \N__43761\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__10047\ : CascadeMux
    port map (
            O => \N__43758\,
            I => \N__43753\
        );

    \I__10046\ : InMux
    port map (
            O => \N__43757\,
            I => \N__43750\
        );

    \I__10045\ : InMux
    port map (
            O => \N__43756\,
            I => \N__43747\
        );

    \I__10044\ : InMux
    port map (
            O => \N__43753\,
            I => \N__43744\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__43750\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__10042\ : LocalMux
    port map (
            O => \N__43747\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__43744\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__10040\ : InMux
    port map (
            O => \N__43737\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__10039\ : CascadeMux
    port map (
            O => \N__43734\,
            I => \N__43729\
        );

    \I__10038\ : InMux
    port map (
            O => \N__43733\,
            I => \N__43726\
        );

    \I__10037\ : InMux
    port map (
            O => \N__43732\,
            I => \N__43723\
        );

    \I__10036\ : InMux
    port map (
            O => \N__43729\,
            I => \N__43720\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__43726\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__10034\ : LocalMux
    port map (
            O => \N__43723\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__43720\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__10032\ : InMux
    port map (
            O => \N__43713\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__10031\ : CascadeMux
    port map (
            O => \N__43710\,
            I => \N__43705\
        );

    \I__10030\ : InMux
    port map (
            O => \N__43709\,
            I => \N__43702\
        );

    \I__10029\ : InMux
    port map (
            O => \N__43708\,
            I => \N__43699\
        );

    \I__10028\ : InMux
    port map (
            O => \N__43705\,
            I => \N__43696\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__43702\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__43699\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__43696\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__10024\ : InMux
    port map (
            O => \N__43689\,
            I => \bfn_18_9_0_\
        );

    \I__10023\ : CascadeMux
    port map (
            O => \N__43686\,
            I => \N__43681\
        );

    \I__10022\ : InMux
    port map (
            O => \N__43685\,
            I => \N__43678\
        );

    \I__10021\ : InMux
    port map (
            O => \N__43684\,
            I => \N__43675\
        );

    \I__10020\ : InMux
    port map (
            O => \N__43681\,
            I => \N__43672\
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__43678\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__10018\ : LocalMux
    port map (
            O => \N__43675\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__43672\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__10016\ : InMux
    port map (
            O => \N__43665\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__10015\ : CascadeMux
    port map (
            O => \N__43662\,
            I => \N__43657\
        );

    \I__10014\ : InMux
    port map (
            O => \N__43661\,
            I => \N__43654\
        );

    \I__10013\ : InMux
    port map (
            O => \N__43660\,
            I => \N__43651\
        );

    \I__10012\ : InMux
    port map (
            O => \N__43657\,
            I => \N__43648\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__43654\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__43651\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__43648\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__10008\ : InMux
    port map (
            O => \N__43641\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__10007\ : CascadeMux
    port map (
            O => \N__43638\,
            I => \N__43633\
        );

    \I__10006\ : InMux
    port map (
            O => \N__43637\,
            I => \N__43630\
        );

    \I__10005\ : InMux
    port map (
            O => \N__43636\,
            I => \N__43627\
        );

    \I__10004\ : InMux
    port map (
            O => \N__43633\,
            I => \N__43624\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__43630\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__43627\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__10001\ : LocalMux
    port map (
            O => \N__43624\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__10000\ : InMux
    port map (
            O => \N__43617\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__9999\ : CascadeMux
    port map (
            O => \N__43614\,
            I => \N__43609\
        );

    \I__9998\ : InMux
    port map (
            O => \N__43613\,
            I => \N__43606\
        );

    \I__9997\ : InMux
    port map (
            O => \N__43612\,
            I => \N__43603\
        );

    \I__9996\ : InMux
    port map (
            O => \N__43609\,
            I => \N__43600\
        );

    \I__9995\ : LocalMux
    port map (
            O => \N__43606\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__43603\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__43600\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9992\ : InMux
    port map (
            O => \N__43593\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__9991\ : CascadeMux
    port map (
            O => \N__43590\,
            I => \N__43585\
        );

    \I__9990\ : InMux
    port map (
            O => \N__43589\,
            I => \N__43582\
        );

    \I__9989\ : InMux
    port map (
            O => \N__43588\,
            I => \N__43579\
        );

    \I__9988\ : InMux
    port map (
            O => \N__43585\,
            I => \N__43576\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__43582\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__43579\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9985\ : LocalMux
    port map (
            O => \N__43576\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9984\ : InMux
    port map (
            O => \N__43569\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__9983\ : CascadeMux
    port map (
            O => \N__43566\,
            I => \N__43561\
        );

    \I__9982\ : InMux
    port map (
            O => \N__43565\,
            I => \N__43558\
        );

    \I__9981\ : InMux
    port map (
            O => \N__43564\,
            I => \N__43555\
        );

    \I__9980\ : InMux
    port map (
            O => \N__43561\,
            I => \N__43552\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__43558\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__43555\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__43552\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9976\ : InMux
    port map (
            O => \N__43545\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__9975\ : CascadeMux
    port map (
            O => \N__43542\,
            I => \N__43537\
        );

    \I__9974\ : InMux
    port map (
            O => \N__43541\,
            I => \N__43534\
        );

    \I__9973\ : InMux
    port map (
            O => \N__43540\,
            I => \N__43531\
        );

    \I__9972\ : InMux
    port map (
            O => \N__43537\,
            I => \N__43528\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__43534\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__43531\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__43528\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9968\ : InMux
    port map (
            O => \N__43521\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__9967\ : CascadeMux
    port map (
            O => \N__43518\,
            I => \N__43513\
        );

    \I__9966\ : InMux
    port map (
            O => \N__43517\,
            I => \N__43510\
        );

    \I__9965\ : InMux
    port map (
            O => \N__43516\,
            I => \N__43507\
        );

    \I__9964\ : InMux
    port map (
            O => \N__43513\,
            I => \N__43504\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__43510\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__43507\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__9961\ : LocalMux
    port map (
            O => \N__43504\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__9960\ : InMux
    port map (
            O => \N__43497\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__9959\ : CascadeMux
    port map (
            O => \N__43494\,
            I => \N__43489\
        );

    \I__9958\ : InMux
    port map (
            O => \N__43493\,
            I => \N__43486\
        );

    \I__9957\ : InMux
    port map (
            O => \N__43492\,
            I => \N__43483\
        );

    \I__9956\ : InMux
    port map (
            O => \N__43489\,
            I => \N__43480\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__43486\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__43483\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__43480\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9952\ : InMux
    port map (
            O => \N__43473\,
            I => \bfn_18_8_0_\
        );

    \I__9951\ : CascadeMux
    port map (
            O => \N__43470\,
            I => \N__43465\
        );

    \I__9950\ : InMux
    port map (
            O => \N__43469\,
            I => \N__43462\
        );

    \I__9949\ : InMux
    port map (
            O => \N__43468\,
            I => \N__43459\
        );

    \I__9948\ : InMux
    port map (
            O => \N__43465\,
            I => \N__43456\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__43462\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__9946\ : LocalMux
    port map (
            O => \N__43459\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__9945\ : LocalMux
    port map (
            O => \N__43456\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__9944\ : InMux
    port map (
            O => \N__43449\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__9943\ : CascadeMux
    port map (
            O => \N__43446\,
            I => \N__43441\
        );

    \I__9942\ : InMux
    port map (
            O => \N__43445\,
            I => \N__43438\
        );

    \I__9941\ : InMux
    port map (
            O => \N__43444\,
            I => \N__43435\
        );

    \I__9940\ : InMux
    port map (
            O => \N__43441\,
            I => \N__43432\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__43438\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__43435\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__43432\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__9936\ : InMux
    port map (
            O => \N__43425\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__9935\ : CascadeMux
    port map (
            O => \N__43422\,
            I => \N__43417\
        );

    \I__9934\ : InMux
    port map (
            O => \N__43421\,
            I => \N__43414\
        );

    \I__9933\ : InMux
    port map (
            O => \N__43420\,
            I => \N__43411\
        );

    \I__9932\ : InMux
    port map (
            O => \N__43417\,
            I => \N__43408\
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__43414\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__43411\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__43408\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__9928\ : InMux
    port map (
            O => \N__43401\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__9927\ : CascadeMux
    port map (
            O => \N__43398\,
            I => \N__43395\
        );

    \I__9926\ : InMux
    port map (
            O => \N__43395\,
            I => \N__43392\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__43392\,
            I => \N__43389\
        );

    \I__9924\ : Odrv4
    port map (
            O => \N__43389\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\
        );

    \I__9923\ : CEMux
    port map (
            O => \N__43386\,
            I => \N__43381\
        );

    \I__9922\ : CEMux
    port map (
            O => \N__43385\,
            I => \N__43377\
        );

    \I__9921\ : CEMux
    port map (
            O => \N__43384\,
            I => \N__43374\
        );

    \I__9920\ : LocalMux
    port map (
            O => \N__43381\,
            I => \N__43371\
        );

    \I__9919\ : CEMux
    port map (
            O => \N__43380\,
            I => \N__43368\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__43377\,
            I => \N__43365\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__43374\,
            I => \N__43362\
        );

    \I__9916\ : Span4Mux_v
    port map (
            O => \N__43371\,
            I => \N__43357\
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__43368\,
            I => \N__43357\
        );

    \I__9914\ : Span4Mux_v
    port map (
            O => \N__43365\,
            I => \N__43352\
        );

    \I__9913\ : Span4Mux_v
    port map (
            O => \N__43362\,
            I => \N__43352\
        );

    \I__9912\ : Span4Mux_v
    port map (
            O => \N__43357\,
            I => \N__43349\
        );

    \I__9911\ : Odrv4
    port map (
            O => \N__43352\,
            I => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9910\ : Odrv4
    port map (
            O => \N__43349\,
            I => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9909\ : CascadeMux
    port map (
            O => \N__43344\,
            I => \N__43336\
        );

    \I__9908\ : CascadeMux
    port map (
            O => \N__43343\,
            I => \N__43333\
        );

    \I__9907\ : InMux
    port map (
            O => \N__43342\,
            I => \N__43319\
        );

    \I__9906\ : InMux
    port map (
            O => \N__43341\,
            I => \N__43319\
        );

    \I__9905\ : InMux
    port map (
            O => \N__43340\,
            I => \N__43319\
        );

    \I__9904\ : InMux
    port map (
            O => \N__43339\,
            I => \N__43319\
        );

    \I__9903\ : InMux
    port map (
            O => \N__43336\,
            I => \N__43306\
        );

    \I__9902\ : InMux
    port map (
            O => \N__43333\,
            I => \N__43306\
        );

    \I__9901\ : InMux
    port map (
            O => \N__43332\,
            I => \N__43306\
        );

    \I__9900\ : InMux
    port map (
            O => \N__43331\,
            I => \N__43306\
        );

    \I__9899\ : InMux
    port map (
            O => \N__43330\,
            I => \N__43306\
        );

    \I__9898\ : InMux
    port map (
            O => \N__43329\,
            I => \N__43306\
        );

    \I__9897\ : InMux
    port map (
            O => \N__43328\,
            I => \N__43303\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__43319\,
            I => \N__43296\
        );

    \I__9895\ : LocalMux
    port map (
            O => \N__43306\,
            I => \N__43293\
        );

    \I__9894\ : LocalMux
    port map (
            O => \N__43303\,
            I => \N__43290\
        );

    \I__9893\ : InMux
    port map (
            O => \N__43302\,
            I => \N__43287\
        );

    \I__9892\ : InMux
    port map (
            O => \N__43301\,
            I => \N__43282\
        );

    \I__9891\ : InMux
    port map (
            O => \N__43300\,
            I => \N__43282\
        );

    \I__9890\ : InMux
    port map (
            O => \N__43299\,
            I => \N__43279\
        );

    \I__9889\ : Span4Mux_v
    port map (
            O => \N__43296\,
            I => \N__43276\
        );

    \I__9888\ : Span4Mux_v
    port map (
            O => \N__43293\,
            I => \N__43271\
        );

    \I__9887\ : Span4Mux_h
    port map (
            O => \N__43290\,
            I => \N__43271\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__43287\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__43282\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__43279\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__9883\ : Odrv4
    port map (
            O => \N__43276\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__9882\ : Odrv4
    port map (
            O => \N__43271\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__9881\ : CascadeMux
    port map (
            O => \N__43260\,
            I => \N__43254\
        );

    \I__9880\ : InMux
    port map (
            O => \N__43259\,
            I => \N__43246\
        );

    \I__9879\ : InMux
    port map (
            O => \N__43258\,
            I => \N__43246\
        );

    \I__9878\ : InMux
    port map (
            O => \N__43257\,
            I => \N__43243\
        );

    \I__9877\ : InMux
    port map (
            O => \N__43254\,
            I => \N__43240\
        );

    \I__9876\ : CascadeMux
    port map (
            O => \N__43253\,
            I => \N__43236\
        );

    \I__9875\ : InMux
    port map (
            O => \N__43252\,
            I => \N__43229\
        );

    \I__9874\ : InMux
    port map (
            O => \N__43251\,
            I => \N__43229\
        );

    \I__9873\ : LocalMux
    port map (
            O => \N__43246\,
            I => \N__43226\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__43243\,
            I => \N__43221\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__43240\,
            I => \N__43221\
        );

    \I__9870\ : InMux
    port map (
            O => \N__43239\,
            I => \N__43218\
        );

    \I__9869\ : InMux
    port map (
            O => \N__43236\,
            I => \N__43215\
        );

    \I__9868\ : InMux
    port map (
            O => \N__43235\,
            I => \N__43210\
        );

    \I__9867\ : InMux
    port map (
            O => \N__43234\,
            I => \N__43210\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__43229\,
            I => \N__43207\
        );

    \I__9865\ : Span4Mux_h
    port map (
            O => \N__43226\,
            I => \N__43204\
        );

    \I__9864\ : Span4Mux_v
    port map (
            O => \N__43221\,
            I => \N__43199\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__43218\,
            I => \N__43199\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__43215\,
            I => measured_delay_tr_15
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__43210\,
            I => measured_delay_tr_15
        );

    \I__9860\ : Odrv4
    port map (
            O => \N__43207\,
            I => measured_delay_tr_15
        );

    \I__9859\ : Odrv4
    port map (
            O => \N__43204\,
            I => measured_delay_tr_15
        );

    \I__9858\ : Odrv4
    port map (
            O => \N__43199\,
            I => measured_delay_tr_15
        );

    \I__9857\ : CascadeMux
    port map (
            O => \N__43188\,
            I => \N__43185\
        );

    \I__9856\ : InMux
    port map (
            O => \N__43185\,
            I => \N__43182\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__43182\,
            I => \N__43179\
        );

    \I__9854\ : Span4Mux_h
    port map (
            O => \N__43179\,
            I => \N__43176\
        );

    \I__9853\ : Odrv4
    port map (
            O => \N__43176\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__9852\ : CascadeMux
    port map (
            O => \N__43173\,
            I => \N__43170\
        );

    \I__9851\ : InMux
    port map (
            O => \N__43170\,
            I => \N__43167\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__43167\,
            I => \N__43164\
        );

    \I__9849\ : Span4Mux_h
    port map (
            O => \N__43164\,
            I => \N__43161\
        );

    \I__9848\ : Odrv4
    port map (
            O => \N__43161\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__9847\ : InMux
    port map (
            O => \N__43158\,
            I => \N__43149\
        );

    \I__9846\ : InMux
    port map (
            O => \N__43157\,
            I => \N__43149\
        );

    \I__9845\ : InMux
    port map (
            O => \N__43156\,
            I => \N__43149\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__43149\,
            I => \N__43145\
        );

    \I__9843\ : InMux
    port map (
            O => \N__43148\,
            I => \N__43142\
        );

    \I__9842\ : Span4Mux_h
    port map (
            O => \N__43145\,
            I => \N__43134\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__43142\,
            I => \N__43131\
        );

    \I__9840\ : InMux
    port map (
            O => \N__43141\,
            I => \N__43128\
        );

    \I__9839\ : InMux
    port map (
            O => \N__43140\,
            I => \N__43119\
        );

    \I__9838\ : InMux
    port map (
            O => \N__43139\,
            I => \N__43119\
        );

    \I__9837\ : InMux
    port map (
            O => \N__43138\,
            I => \N__43119\
        );

    \I__9836\ : InMux
    port map (
            O => \N__43137\,
            I => \N__43119\
        );

    \I__9835\ : Odrv4
    port map (
            O => \N__43134\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\
        );

    \I__9834\ : Odrv4
    port map (
            O => \N__43131\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__43128\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\
        );

    \I__9832\ : LocalMux
    port map (
            O => \N__43119\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\
        );

    \I__9831\ : InMux
    port map (
            O => \N__43110\,
            I => \N__43106\
        );

    \I__9830\ : InMux
    port map (
            O => \N__43109\,
            I => \N__43102\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__43106\,
            I => \N__43099\
        );

    \I__9828\ : InMux
    port map (
            O => \N__43105\,
            I => \N__43096\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__43102\,
            I => \N__43093\
        );

    \I__9826\ : Span4Mux_h
    port map (
            O => \N__43099\,
            I => \N__43088\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__43096\,
            I => \N__43088\
        );

    \I__9824\ : Odrv12
    port map (
            O => \N__43093\,
            I => measured_delay_tr_10
        );

    \I__9823\ : Odrv4
    port map (
            O => \N__43088\,
            I => measured_delay_tr_10
        );

    \I__9822\ : CascadeMux
    port map (
            O => \N__43083\,
            I => \N__43080\
        );

    \I__9821\ : InMux
    port map (
            O => \N__43080\,
            I => \N__43077\
        );

    \I__9820\ : LocalMux
    port map (
            O => \N__43077\,
            I => \N__43074\
        );

    \I__9819\ : Span4Mux_v
    port map (
            O => \N__43074\,
            I => \N__43071\
        );

    \I__9818\ : Odrv4
    port map (
            O => \N__43071\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__9817\ : CEMux
    port map (
            O => \N__43068\,
            I => \N__43064\
        );

    \I__9816\ : CEMux
    port map (
            O => \N__43067\,
            I => \N__43059\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__43064\,
            I => \N__43056\
        );

    \I__9814\ : CEMux
    port map (
            O => \N__43063\,
            I => \N__43053\
        );

    \I__9813\ : CEMux
    port map (
            O => \N__43062\,
            I => \N__43050\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__43059\,
            I => \N__43047\
        );

    \I__9811\ : Span4Mux_v
    port map (
            O => \N__43056\,
            I => \N__43041\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__43053\,
            I => \N__43041\
        );

    \I__9809\ : LocalMux
    port map (
            O => \N__43050\,
            I => \N__43038\
        );

    \I__9808\ : Span4Mux_h
    port map (
            O => \N__43047\,
            I => \N__43035\
        );

    \I__9807\ : CEMux
    port map (
            O => \N__43046\,
            I => \N__43032\
        );

    \I__9806\ : Span4Mux_v
    port map (
            O => \N__43041\,
            I => \N__43029\
        );

    \I__9805\ : Span4Mux_v
    port map (
            O => \N__43038\,
            I => \N__43026\
        );

    \I__9804\ : Span4Mux_v
    port map (
            O => \N__43035\,
            I => \N__43021\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__43032\,
            I => \N__43021\
        );

    \I__9802\ : Span4Mux_h
    port map (
            O => \N__43029\,
            I => \N__43018\
        );

    \I__9801\ : Span4Mux_h
    port map (
            O => \N__43026\,
            I => \N__43015\
        );

    \I__9800\ : Span4Mux_h
    port map (
            O => \N__43021\,
            I => \N__43012\
        );

    \I__9799\ : Odrv4
    port map (
            O => \N__43018\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9798\ : Odrv4
    port map (
            O => \N__43015\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9797\ : Odrv4
    port map (
            O => \N__43012\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9796\ : InMux
    port map (
            O => \N__43005\,
            I => \N__43002\
        );

    \I__9795\ : LocalMux
    port map (
            O => \N__43002\,
            I => \N__42996\
        );

    \I__9794\ : InMux
    port map (
            O => \N__43001\,
            I => \N__42993\
        );

    \I__9793\ : InMux
    port map (
            O => \N__43000\,
            I => \N__42990\
        );

    \I__9792\ : InMux
    port map (
            O => \N__42999\,
            I => \N__42987\
        );

    \I__9791\ : Span4Mux_h
    port map (
            O => \N__42996\,
            I => \N__42984\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__42993\,
            I => \N__42981\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__42990\,
            I => \N__42978\
        );

    \I__9788\ : LocalMux
    port map (
            O => \N__42987\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__9787\ : Odrv4
    port map (
            O => \N__42984\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__9786\ : Odrv12
    port map (
            O => \N__42981\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__9785\ : Odrv4
    port map (
            O => \N__42978\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__9784\ : InMux
    port map (
            O => \N__42969\,
            I => \N__42964\
        );

    \I__9783\ : InMux
    port map (
            O => \N__42968\,
            I => \N__42961\
        );

    \I__9782\ : InMux
    port map (
            O => \N__42967\,
            I => \N__42958\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__42964\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__42961\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__42958\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9778\ : InMux
    port map (
            O => \N__42951\,
            I => \bfn_18_7_0_\
        );

    \I__9777\ : InMux
    port map (
            O => \N__42948\,
            I => \N__42943\
        );

    \I__9776\ : InMux
    port map (
            O => \N__42947\,
            I => \N__42940\
        );

    \I__9775\ : InMux
    port map (
            O => \N__42946\,
            I => \N__42937\
        );

    \I__9774\ : LocalMux
    port map (
            O => \N__42943\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__42940\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__9772\ : LocalMux
    port map (
            O => \N__42937\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__9771\ : InMux
    port map (
            O => \N__42930\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__9770\ : CascadeMux
    port map (
            O => \N__42927\,
            I => \N__42922\
        );

    \I__9769\ : InMux
    port map (
            O => \N__42926\,
            I => \N__42919\
        );

    \I__9768\ : InMux
    port map (
            O => \N__42925\,
            I => \N__42916\
        );

    \I__9767\ : InMux
    port map (
            O => \N__42922\,
            I => \N__42913\
        );

    \I__9766\ : LocalMux
    port map (
            O => \N__42919\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__42916\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__42913\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9763\ : InMux
    port map (
            O => \N__42906\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__9762\ : InMux
    port map (
            O => \N__42903\,
            I => \N__42898\
        );

    \I__9761\ : CascadeMux
    port map (
            O => \N__42902\,
            I => \N__42895\
        );

    \I__9760\ : InMux
    port map (
            O => \N__42901\,
            I => \N__42890\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__42898\,
            I => \N__42887\
        );

    \I__9758\ : InMux
    port map (
            O => \N__42895\,
            I => \N__42884\
        );

    \I__9757\ : InMux
    port map (
            O => \N__42894\,
            I => \N__42881\
        );

    \I__9756\ : InMux
    port map (
            O => \N__42893\,
            I => \N__42878\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__42890\,
            I => \N__42873\
        );

    \I__9754\ : Span4Mux_h
    port map (
            O => \N__42887\,
            I => \N__42873\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__42884\,
            I => measured_delay_tr_14
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__42881\,
            I => measured_delay_tr_14
        );

    \I__9751\ : LocalMux
    port map (
            O => \N__42878\,
            I => measured_delay_tr_14
        );

    \I__9750\ : Odrv4
    port map (
            O => \N__42873\,
            I => measured_delay_tr_14
        );

    \I__9749\ : InMux
    port map (
            O => \N__42864\,
            I => \N__42861\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__42861\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\
        );

    \I__9747\ : InMux
    port map (
            O => \N__42858\,
            I => \N__42854\
        );

    \I__9746\ : InMux
    port map (
            O => \N__42857\,
            I => \N__42851\
        );

    \I__9745\ : LocalMux
    port map (
            O => \N__42854\,
            I => \N__42848\
        );

    \I__9744\ : LocalMux
    port map (
            O => \N__42851\,
            I => \N__42845\
        );

    \I__9743\ : Span12Mux_v
    port map (
            O => \N__42848\,
            I => \N__42841\
        );

    \I__9742\ : Span4Mux_h
    port map (
            O => \N__42845\,
            I => \N__42838\
        );

    \I__9741\ : InMux
    port map (
            O => \N__42844\,
            I => \N__42835\
        );

    \I__9740\ : Odrv12
    port map (
            O => \N__42841\,
            I => measured_delay_tr_6
        );

    \I__9739\ : Odrv4
    port map (
            O => \N__42838\,
            I => measured_delay_tr_6
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__42835\,
            I => measured_delay_tr_6
        );

    \I__9737\ : CascadeMux
    port map (
            O => \N__42828\,
            I => \N__42825\
        );

    \I__9736\ : InMux
    port map (
            O => \N__42825\,
            I => \N__42818\
        );

    \I__9735\ : InMux
    port map (
            O => \N__42824\,
            I => \N__42815\
        );

    \I__9734\ : InMux
    port map (
            O => \N__42823\,
            I => \N__42808\
        );

    \I__9733\ : InMux
    port map (
            O => \N__42822\,
            I => \N__42808\
        );

    \I__9732\ : InMux
    port map (
            O => \N__42821\,
            I => \N__42808\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__42818\,
            I => \N__42803\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__42815\,
            I => \N__42803\
        );

    \I__9729\ : LocalMux
    port map (
            O => \N__42808\,
            I => \N__42800\
        );

    \I__9728\ : Span4Mux_v
    port map (
            O => \N__42803\,
            I => \N__42796\
        );

    \I__9727\ : Span4Mux_v
    port map (
            O => \N__42800\,
            I => \N__42793\
        );

    \I__9726\ : InMux
    port map (
            O => \N__42799\,
            I => \N__42790\
        );

    \I__9725\ : Odrv4
    port map (
            O => \N__42796\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\
        );

    \I__9724\ : Odrv4
    port map (
            O => \N__42793\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__42790\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\
        );

    \I__9722\ : CascadeMux
    port map (
            O => \N__42783\,
            I => \N__42778\
        );

    \I__9721\ : InMux
    port map (
            O => \N__42782\,
            I => \N__42768\
        );

    \I__9720\ : InMux
    port map (
            O => \N__42781\,
            I => \N__42768\
        );

    \I__9719\ : InMux
    port map (
            O => \N__42778\,
            I => \N__42761\
        );

    \I__9718\ : InMux
    port map (
            O => \N__42777\,
            I => \N__42761\
        );

    \I__9717\ : InMux
    port map (
            O => \N__42776\,
            I => \N__42761\
        );

    \I__9716\ : InMux
    port map (
            O => \N__42775\,
            I => \N__42758\
        );

    \I__9715\ : InMux
    port map (
            O => \N__42774\,
            I => \N__42753\
        );

    \I__9714\ : InMux
    port map (
            O => \N__42773\,
            I => \N__42753\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__42768\,
            I => \N__42746\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__42761\,
            I => \N__42746\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__42758\,
            I => \N__42743\
        );

    \I__9710\ : LocalMux
    port map (
            O => \N__42753\,
            I => \N__42740\
        );

    \I__9709\ : InMux
    port map (
            O => \N__42752\,
            I => \N__42736\
        );

    \I__9708\ : InMux
    port map (
            O => \N__42751\,
            I => \N__42733\
        );

    \I__9707\ : Span4Mux_h
    port map (
            O => \N__42746\,
            I => \N__42730\
        );

    \I__9706\ : Span4Mux_v
    port map (
            O => \N__42743\,
            I => \N__42725\
        );

    \I__9705\ : Span4Mux_v
    port map (
            O => \N__42740\,
            I => \N__42725\
        );

    \I__9704\ : InMux
    port map (
            O => \N__42739\,
            I => \N__42722\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__42736\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__42733\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\
        );

    \I__9701\ : Odrv4
    port map (
            O => \N__42730\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\
        );

    \I__9700\ : Odrv4
    port map (
            O => \N__42725\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\
        );

    \I__9699\ : LocalMux
    port map (
            O => \N__42722\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\
        );

    \I__9698\ : CascadeMux
    port map (
            O => \N__42711\,
            I => \N__42708\
        );

    \I__9697\ : InMux
    port map (
            O => \N__42708\,
            I => \N__42705\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__42705\,
            I => \N__42702\
        );

    \I__9695\ : Odrv4
    port map (
            O => \N__42702\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_6\
        );

    \I__9694\ : CascadeMux
    port map (
            O => \N__42699\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15_cascade_\
        );

    \I__9693\ : CascadeMux
    port map (
            O => \N__42696\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13_cascade_\
        );

    \I__9692\ : CascadeMux
    port map (
            O => \N__42693\,
            I => \N__42690\
        );

    \I__9691\ : InMux
    port map (
            O => \N__42690\,
            I => \N__42687\
        );

    \I__9690\ : LocalMux
    port map (
            O => \N__42687\,
            I => \N__42684\
        );

    \I__9689\ : Odrv4
    port map (
            O => \N__42684\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\
        );

    \I__9688\ : InMux
    port map (
            O => \N__42681\,
            I => \N__42676\
        );

    \I__9687\ : InMux
    port map (
            O => \N__42680\,
            I => \N__42673\
        );

    \I__9686\ : InMux
    port map (
            O => \N__42679\,
            I => \N__42670\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__42676\,
            I => \N__42667\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__42673\,
            I => \N__42662\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__42670\,
            I => \N__42662\
        );

    \I__9682\ : Odrv12
    port map (
            O => \N__42667\,
            I => measured_delay_tr_11
        );

    \I__9681\ : Odrv4
    port map (
            O => \N__42662\,
            I => measured_delay_tr_11
        );

    \I__9680\ : CascadeMux
    port map (
            O => \N__42657\,
            I => \N__42654\
        );

    \I__9679\ : InMux
    port map (
            O => \N__42654\,
            I => \N__42651\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__42651\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\
        );

    \I__9677\ : InMux
    port map (
            O => \N__42648\,
            I => \N__42643\
        );

    \I__9676\ : InMux
    port map (
            O => \N__42647\,
            I => \N__42640\
        );

    \I__9675\ : InMux
    port map (
            O => \N__42646\,
            I => \N__42637\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__42643\,
            I => \N__42634\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__42640\,
            I => \N__42629\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__42637\,
            I => \N__42629\
        );

    \I__9671\ : Odrv12
    port map (
            O => \N__42634\,
            I => measured_delay_tr_12
        );

    \I__9670\ : Odrv4
    port map (
            O => \N__42629\,
            I => measured_delay_tr_12
        );

    \I__9669\ : CascadeMux
    port map (
            O => \N__42624\,
            I => \N__42621\
        );

    \I__9668\ : InMux
    port map (
            O => \N__42621\,
            I => \N__42618\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__42618\,
            I => \N__42615\
        );

    \I__9666\ : Odrv12
    port map (
            O => \N__42615\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\
        );

    \I__9665\ : CascadeMux
    port map (
            O => \N__42612\,
            I => \N__42608\
        );

    \I__9664\ : InMux
    port map (
            O => \N__42611\,
            I => \N__42604\
        );

    \I__9663\ : InMux
    port map (
            O => \N__42608\,
            I => \N__42601\
        );

    \I__9662\ : InMux
    port map (
            O => \N__42607\,
            I => \N__42598\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__42604\,
            I => \N__42595\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__42601\,
            I => \N__42592\
        );

    \I__9659\ : LocalMux
    port map (
            O => \N__42598\,
            I => \N__42589\
        );

    \I__9658\ : Span4Mux_v
    port map (
            O => \N__42595\,
            I => \N__42584\
        );

    \I__9657\ : Span4Mux_h
    port map (
            O => \N__42592\,
            I => \N__42584\
        );

    \I__9656\ : Odrv12
    port map (
            O => \N__42589\,
            I => measured_delay_tr_13
        );

    \I__9655\ : Odrv4
    port map (
            O => \N__42584\,
            I => measured_delay_tr_13
        );

    \I__9654\ : CascadeMux
    port map (
            O => \N__42579\,
            I => \N__42576\
        );

    \I__9653\ : InMux
    port map (
            O => \N__42576\,
            I => \N__42573\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__42573\,
            I => \N__42570\
        );

    \I__9651\ : Odrv4
    port map (
            O => \N__42570\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\
        );

    \I__9650\ : InMux
    port map (
            O => \N__42567\,
            I => \N__42564\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__42564\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\
        );

    \I__9648\ : InMux
    port map (
            O => \N__42561\,
            I => \N__42558\
        );

    \I__9647\ : LocalMux
    port map (
            O => \N__42558\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\
        );

    \I__9646\ : InMux
    port map (
            O => \N__42555\,
            I => \N__42552\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__42552\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\
        );

    \I__9644\ : InMux
    port map (
            O => \N__42549\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__9643\ : CascadeMux
    port map (
            O => \N__42546\,
            I => \N__42543\
        );

    \I__9642\ : InMux
    port map (
            O => \N__42543\,
            I => \N__42540\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__42540\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__9640\ : CascadeMux
    port map (
            O => \N__42537\,
            I => \N__42534\
        );

    \I__9639\ : InMux
    port map (
            O => \N__42534\,
            I => \N__42531\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__42531\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__9637\ : CascadeMux
    port map (
            O => \N__42528\,
            I => \N__42525\
        );

    \I__9636\ : InMux
    port map (
            O => \N__42525\,
            I => \N__42522\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__42522\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__9634\ : CascadeMux
    port map (
            O => \N__42519\,
            I => \N__42516\
        );

    \I__9633\ : InMux
    port map (
            O => \N__42516\,
            I => \N__42513\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__42513\,
            I => \N__42510\
        );

    \I__9631\ : Odrv4
    port map (
            O => \N__42510\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\
        );

    \I__9630\ : InMux
    port map (
            O => \N__42507\,
            I => \N__42503\
        );

    \I__9629\ : InMux
    port map (
            O => \N__42506\,
            I => \N__42500\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__42503\,
            I => \N__42497\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__42500\,
            I => \N__42494\
        );

    \I__9626\ : Span4Mux_h
    port map (
            O => \N__42497\,
            I => \N__42490\
        );

    \I__9625\ : Span4Mux_h
    port map (
            O => \N__42494\,
            I => \N__42487\
        );

    \I__9624\ : InMux
    port map (
            O => \N__42493\,
            I => \N__42484\
        );

    \I__9623\ : Odrv4
    port map (
            O => \N__42490\,
            I => measured_delay_tr_7
        );

    \I__9622\ : Odrv4
    port map (
            O => \N__42487\,
            I => measured_delay_tr_7
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__42484\,
            I => measured_delay_tr_7
        );

    \I__9620\ : CascadeMux
    port map (
            O => \N__42477\,
            I => \N__42474\
        );

    \I__9619\ : InMux
    port map (
            O => \N__42474\,
            I => \N__42471\
        );

    \I__9618\ : LocalMux
    port map (
            O => \N__42471\,
            I => \N__42468\
        );

    \I__9617\ : Odrv4
    port map (
            O => \N__42468\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\
        );

    \I__9616\ : CascadeMux
    port map (
            O => \N__42465\,
            I => \N__42462\
        );

    \I__9615\ : InMux
    port map (
            O => \N__42462\,
            I => \N__42459\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__42459\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__9613\ : InMux
    port map (
            O => \N__42456\,
            I => \N__42453\
        );

    \I__9612\ : LocalMux
    port map (
            O => \N__42453\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__9611\ : InMux
    port map (
            O => \N__42450\,
            I => \N__42447\
        );

    \I__9610\ : LocalMux
    port map (
            O => \N__42447\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__9609\ : CascadeMux
    port map (
            O => \N__42444\,
            I => \N__42441\
        );

    \I__9608\ : InMux
    port map (
            O => \N__42441\,
            I => \N__42438\
        );

    \I__9607\ : LocalMux
    port map (
            O => \N__42438\,
            I => \N__42435\
        );

    \I__9606\ : Odrv12
    port map (
            O => \N__42435\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__9605\ : InMux
    port map (
            O => \N__42432\,
            I => \N__42429\
        );

    \I__9604\ : LocalMux
    port map (
            O => \N__42429\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__9603\ : CascadeMux
    port map (
            O => \N__42426\,
            I => \N__42423\
        );

    \I__9602\ : InMux
    port map (
            O => \N__42423\,
            I => \N__42420\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__42420\,
            I => \N__42417\
        );

    \I__9600\ : Odrv12
    port map (
            O => \N__42417\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__9599\ : InMux
    port map (
            O => \N__42414\,
            I => \N__42411\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__42411\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__9597\ : CascadeMux
    port map (
            O => \N__42408\,
            I => \N__42405\
        );

    \I__9596\ : InMux
    port map (
            O => \N__42405\,
            I => \N__42402\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__42402\,
            I => \N__42399\
        );

    \I__9594\ : Span4Mux_h
    port map (
            O => \N__42399\,
            I => \N__42396\
        );

    \I__9593\ : Odrv4
    port map (
            O => \N__42396\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__9592\ : InMux
    port map (
            O => \N__42393\,
            I => \N__42390\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__42390\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__9590\ : CascadeMux
    port map (
            O => \N__42387\,
            I => \N__42384\
        );

    \I__9589\ : InMux
    port map (
            O => \N__42384\,
            I => \N__42381\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__42381\,
            I => \N__42378\
        );

    \I__9587\ : Odrv4
    port map (
            O => \N__42378\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__9586\ : InMux
    port map (
            O => \N__42375\,
            I => \N__42372\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__42372\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__9584\ : InMux
    port map (
            O => \N__42369\,
            I => \N__42366\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__42366\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__9582\ : InMux
    port map (
            O => \N__42363\,
            I => \N__42360\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__42360\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\
        );

    \I__9580\ : CascadeMux
    port map (
            O => \N__42357\,
            I => \N__42354\
        );

    \I__9579\ : InMux
    port map (
            O => \N__42354\,
            I => \N__42351\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__42351\,
            I => \N__42348\
        );

    \I__9577\ : Odrv4
    port map (
            O => \N__42348\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__9576\ : InMux
    port map (
            O => \N__42345\,
            I => \N__42342\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__42342\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__9574\ : CascadeMux
    port map (
            O => \N__42339\,
            I => \N__42336\
        );

    \I__9573\ : InMux
    port map (
            O => \N__42336\,
            I => \N__42333\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__42333\,
            I => \N__42330\
        );

    \I__9571\ : Span4Mux_v
    port map (
            O => \N__42330\,
            I => \N__42327\
        );

    \I__9570\ : Odrv4
    port map (
            O => \N__42327\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__9569\ : InMux
    port map (
            O => \N__42324\,
            I => \N__42321\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__42321\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__9567\ : CascadeMux
    port map (
            O => \N__42318\,
            I => \N__42315\
        );

    \I__9566\ : InMux
    port map (
            O => \N__42315\,
            I => \N__42312\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__42312\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__9564\ : InMux
    port map (
            O => \N__42309\,
            I => \N__42306\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__42306\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__9562\ : CascadeMux
    port map (
            O => \N__42303\,
            I => \N__42300\
        );

    \I__9561\ : InMux
    port map (
            O => \N__42300\,
            I => \N__42297\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__42297\,
            I => \N__42294\
        );

    \I__9559\ : Odrv4
    port map (
            O => \N__42294\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__9558\ : InMux
    port map (
            O => \N__42291\,
            I => \N__42288\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__42288\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__9556\ : CascadeMux
    port map (
            O => \N__42285\,
            I => \N__42282\
        );

    \I__9555\ : InMux
    port map (
            O => \N__42282\,
            I => \N__42279\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__42279\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__9553\ : InMux
    port map (
            O => \N__42276\,
            I => \N__42273\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__42273\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__9551\ : CascadeMux
    port map (
            O => \N__42270\,
            I => \N__42267\
        );

    \I__9550\ : InMux
    port map (
            O => \N__42267\,
            I => \N__42264\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__42264\,
            I => \N__42261\
        );

    \I__9548\ : Odrv4
    port map (
            O => \N__42261\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__9547\ : InMux
    port map (
            O => \N__42258\,
            I => \N__42255\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__42255\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__9545\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42249\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__42249\,
            I => \N__42246\
        );

    \I__9543\ : Span4Mux_h
    port map (
            O => \N__42246\,
            I => \N__42243\
        );

    \I__9542\ : Odrv4
    port map (
            O => \N__42243\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__9541\ : CascadeMux
    port map (
            O => \N__42240\,
            I => \N__42237\
        );

    \I__9540\ : InMux
    port map (
            O => \N__42237\,
            I => \N__42234\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__42234\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__9538\ : CascadeMux
    port map (
            O => \N__42231\,
            I => \N__42227\
        );

    \I__9537\ : CascadeMux
    port map (
            O => \N__42230\,
            I => \N__42214\
        );

    \I__9536\ : InMux
    port map (
            O => \N__42227\,
            I => \N__42209\
        );

    \I__9535\ : InMux
    port map (
            O => \N__42226\,
            I => \N__42209\
        );

    \I__9534\ : CascadeMux
    port map (
            O => \N__42225\,
            I => \N__42202\
        );

    \I__9533\ : CascadeMux
    port map (
            O => \N__42224\,
            I => \N__42199\
        );

    \I__9532\ : CascadeMux
    port map (
            O => \N__42223\,
            I => \N__42196\
        );

    \I__9531\ : CascadeMux
    port map (
            O => \N__42222\,
            I => \N__42193\
        );

    \I__9530\ : CascadeMux
    port map (
            O => \N__42221\,
            I => \N__42189\
        );

    \I__9529\ : CascadeMux
    port map (
            O => \N__42220\,
            I => \N__42186\
        );

    \I__9528\ : CascadeMux
    port map (
            O => \N__42219\,
            I => \N__42183\
        );

    \I__9527\ : CascadeMux
    port map (
            O => \N__42218\,
            I => \N__42180\
        );

    \I__9526\ : InMux
    port map (
            O => \N__42217\,
            I => \N__42171\
        );

    \I__9525\ : InMux
    port map (
            O => \N__42214\,
            I => \N__42171\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__42209\,
            I => \N__42168\
        );

    \I__9523\ : InMux
    port map (
            O => \N__42208\,
            I => \N__42151\
        );

    \I__9522\ : InMux
    port map (
            O => \N__42207\,
            I => \N__42151\
        );

    \I__9521\ : InMux
    port map (
            O => \N__42206\,
            I => \N__42151\
        );

    \I__9520\ : InMux
    port map (
            O => \N__42205\,
            I => \N__42151\
        );

    \I__9519\ : InMux
    port map (
            O => \N__42202\,
            I => \N__42151\
        );

    \I__9518\ : InMux
    port map (
            O => \N__42199\,
            I => \N__42151\
        );

    \I__9517\ : InMux
    port map (
            O => \N__42196\,
            I => \N__42151\
        );

    \I__9516\ : InMux
    port map (
            O => \N__42193\,
            I => \N__42151\
        );

    \I__9515\ : CascadeMux
    port map (
            O => \N__42192\,
            I => \N__42148\
        );

    \I__9514\ : InMux
    port map (
            O => \N__42189\,
            I => \N__42131\
        );

    \I__9513\ : InMux
    port map (
            O => \N__42186\,
            I => \N__42131\
        );

    \I__9512\ : InMux
    port map (
            O => \N__42183\,
            I => \N__42131\
        );

    \I__9511\ : InMux
    port map (
            O => \N__42180\,
            I => \N__42131\
        );

    \I__9510\ : InMux
    port map (
            O => \N__42179\,
            I => \N__42131\
        );

    \I__9509\ : InMux
    port map (
            O => \N__42178\,
            I => \N__42131\
        );

    \I__9508\ : InMux
    port map (
            O => \N__42177\,
            I => \N__42131\
        );

    \I__9507\ : InMux
    port map (
            O => \N__42176\,
            I => \N__42131\
        );

    \I__9506\ : LocalMux
    port map (
            O => \N__42171\,
            I => \N__42122\
        );

    \I__9505\ : Span4Mux_v
    port map (
            O => \N__42168\,
            I => \N__42122\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__42151\,
            I => \N__42122\
        );

    \I__9503\ : InMux
    port map (
            O => \N__42148\,
            I => \N__42119\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__42131\,
            I => \N__42116\
        );

    \I__9501\ : InMux
    port map (
            O => \N__42130\,
            I => \N__42112\
        );

    \I__9500\ : InMux
    port map (
            O => \N__42129\,
            I => \N__42109\
        );

    \I__9499\ : Span4Mux_h
    port map (
            O => \N__42122\,
            I => \N__42106\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__42119\,
            I => \N__42101\
        );

    \I__9497\ : Span4Mux_v
    port map (
            O => \N__42116\,
            I => \N__42101\
        );

    \I__9496\ : InMux
    port map (
            O => \N__42115\,
            I => \N__42098\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__42112\,
            I => \N__42095\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__42109\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9493\ : Odrv4
    port map (
            O => \N__42106\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9492\ : Odrv4
    port map (
            O => \N__42101\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__42098\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9490\ : Odrv12
    port map (
            O => \N__42095\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9489\ : InMux
    port map (
            O => \N__42084\,
            I => \N__42081\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__42081\,
            I => \N__42078\
        );

    \I__9487\ : Span4Mux_h
    port map (
            O => \N__42078\,
            I => \N__42075\
        );

    \I__9486\ : Odrv4
    port map (
            O => \N__42075\,
            I => \phase_controller_inst1.start_timer_tr_0_sqmuxa\
        );

    \I__9485\ : InMux
    port map (
            O => \N__42072\,
            I => \N__42068\
        );

    \I__9484\ : InMux
    port map (
            O => \N__42071\,
            I => \N__42065\
        );

    \I__9483\ : LocalMux
    port map (
            O => \N__42068\,
            I => \N__42062\
        );

    \I__9482\ : LocalMux
    port map (
            O => \N__42065\,
            I => \N__42059\
        );

    \I__9481\ : Span4Mux_h
    port map (
            O => \N__42062\,
            I => \N__42056\
        );

    \I__9480\ : Span4Mux_v
    port map (
            O => \N__42059\,
            I => \N__42051\
        );

    \I__9479\ : Span4Mux_v
    port map (
            O => \N__42056\,
            I => \N__42048\
        );

    \I__9478\ : InMux
    port map (
            O => \N__42055\,
            I => \N__42045\
        );

    \I__9477\ : InMux
    port map (
            O => \N__42054\,
            I => \N__42042\
        );

    \I__9476\ : Odrv4
    port map (
            O => \N__42051\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__9475\ : Odrv4
    port map (
            O => \N__42048\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__42045\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__9473\ : LocalMux
    port map (
            O => \N__42042\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__9472\ : InMux
    port map (
            O => \N__42033\,
            I => \N__42030\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__42030\,
            I => \N__42026\
        );

    \I__9470\ : InMux
    port map (
            O => \N__42029\,
            I => \N__42023\
        );

    \I__9469\ : Span4Mux_h
    port map (
            O => \N__42026\,
            I => \N__42020\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__42023\,
            I => \N__42017\
        );

    \I__9467\ : Odrv4
    port map (
            O => \N__42020\,
            I => \phase_controller_inst1.N_231\
        );

    \I__9466\ : Odrv4
    port map (
            O => \N__42017\,
            I => \phase_controller_inst1.N_231\
        );

    \I__9465\ : CascadeMux
    port map (
            O => \N__42012\,
            I => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_\
        );

    \I__9464\ : InMux
    port map (
            O => \N__42009\,
            I => \N__42004\
        );

    \I__9463\ : InMux
    port map (
            O => \N__42008\,
            I => \N__42001\
        );

    \I__9462\ : InMux
    port map (
            O => \N__42007\,
            I => \N__41998\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__42004\,
            I => \N__41990\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__42001\,
            I => \N__41990\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__41998\,
            I => \N__41990\
        );

    \I__9458\ : InMux
    port map (
            O => \N__41997\,
            I => \N__41987\
        );

    \I__9457\ : Span4Mux_v
    port map (
            O => \N__41990\,
            I => \N__41984\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__41987\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__9455\ : Odrv4
    port map (
            O => \N__41984\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__9454\ : CascadeMux
    port map (
            O => \N__41979\,
            I => \N__41976\
        );

    \I__9453\ : InMux
    port map (
            O => \N__41976\,
            I => \N__41973\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__41973\,
            I => \N__41970\
        );

    \I__9451\ : Odrv4
    port map (
            O => \N__41970\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__9450\ : InMux
    port map (
            O => \N__41967\,
            I => \N__41964\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__41964\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__9448\ : InMux
    port map (
            O => \N__41961\,
            I => \N__41958\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__41958\,
            I => \N__41954\
        );

    \I__9446\ : InMux
    port map (
            O => \N__41957\,
            I => \N__41951\
        );

    \I__9445\ : Odrv12
    port map (
            O => \N__41954\,
            I => \delay_measurement_inst.elapsed_time_hc_26\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__41951\,
            I => \delay_measurement_inst.elapsed_time_hc_26\
        );

    \I__9443\ : InMux
    port map (
            O => \N__41946\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__9442\ : InMux
    port map (
            O => \N__41943\,
            I => \N__41940\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__41940\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__9440\ : InMux
    port map (
            O => \N__41937\,
            I => \bfn_17_11_0_\
        );

    \I__9439\ : InMux
    port map (
            O => \N__41934\,
            I => \N__41931\
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__41931\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__9437\ : InMux
    port map (
            O => \N__41928\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__9436\ : InMux
    port map (
            O => \N__41925\,
            I => \N__41922\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__41922\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__9434\ : InMux
    port map (
            O => \N__41919\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__9433\ : CascadeMux
    port map (
            O => \N__41916\,
            I => \N__41913\
        );

    \I__9432\ : InMux
    port map (
            O => \N__41913\,
            I => \N__41910\
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__41910\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30\
        );

    \I__9430\ : InMux
    port map (
            O => \N__41907\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__9429\ : InMux
    port map (
            O => \N__41904\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__9428\ : CascadeMux
    port map (
            O => \N__41901\,
            I => \N__41896\
        );

    \I__9427\ : CascadeMux
    port map (
            O => \N__41900\,
            I => \N__41889\
        );

    \I__9426\ : CascadeMux
    port map (
            O => \N__41899\,
            I => \N__41886\
        );

    \I__9425\ : InMux
    port map (
            O => \N__41896\,
            I => \N__41881\
        );

    \I__9424\ : InMux
    port map (
            O => \N__41895\,
            I => \N__41881\
        );

    \I__9423\ : CascadeMux
    port map (
            O => \N__41894\,
            I => \N__41876\
        );

    \I__9422\ : CascadeMux
    port map (
            O => \N__41893\,
            I => \N__41873\
        );

    \I__9421\ : CascadeMux
    port map (
            O => \N__41892\,
            I => \N__41870\
        );

    \I__9420\ : InMux
    port map (
            O => \N__41889\,
            I => \N__41866\
        );

    \I__9419\ : InMux
    port map (
            O => \N__41886\,
            I => \N__41863\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__41881\,
            I => \N__41860\
        );

    \I__9417\ : InMux
    port map (
            O => \N__41880\,
            I => \N__41857\
        );

    \I__9416\ : InMux
    port map (
            O => \N__41879\,
            I => \N__41854\
        );

    \I__9415\ : InMux
    port map (
            O => \N__41876\,
            I => \N__41849\
        );

    \I__9414\ : InMux
    port map (
            O => \N__41873\,
            I => \N__41842\
        );

    \I__9413\ : InMux
    port map (
            O => \N__41870\,
            I => \N__41842\
        );

    \I__9412\ : InMux
    port map (
            O => \N__41869\,
            I => \N__41842\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__41866\,
            I => \N__41839\
        );

    \I__9410\ : LocalMux
    port map (
            O => \N__41863\,
            I => \N__41836\
        );

    \I__9409\ : Span4Mux_v
    port map (
            O => \N__41860\,
            I => \N__41831\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__41857\,
            I => \N__41831\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__41854\,
            I => \N__41828\
        );

    \I__9406\ : InMux
    port map (
            O => \N__41853\,
            I => \N__41825\
        );

    \I__9405\ : CascadeMux
    port map (
            O => \N__41852\,
            I => \N__41821\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__41849\,
            I => \N__41818\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__41842\,
            I => \N__41815\
        );

    \I__9402\ : Span4Mux_v
    port map (
            O => \N__41839\,
            I => \N__41812\
        );

    \I__9401\ : Span4Mux_h
    port map (
            O => \N__41836\,
            I => \N__41807\
        );

    \I__9400\ : Span4Mux_h
    port map (
            O => \N__41831\,
            I => \N__41807\
        );

    \I__9399\ : Span4Mux_v
    port map (
            O => \N__41828\,
            I => \N__41802\
        );

    \I__9398\ : LocalMux
    port map (
            O => \N__41825\,
            I => \N__41802\
        );

    \I__9397\ : InMux
    port map (
            O => \N__41824\,
            I => \N__41799\
        );

    \I__9396\ : InMux
    port map (
            O => \N__41821\,
            I => \N__41795\
        );

    \I__9395\ : Span4Mux_v
    port map (
            O => \N__41818\,
            I => \N__41790\
        );

    \I__9394\ : Span4Mux_v
    port map (
            O => \N__41815\,
            I => \N__41790\
        );

    \I__9393\ : Span4Mux_h
    port map (
            O => \N__41812\,
            I => \N__41785\
        );

    \I__9392\ : Span4Mux_v
    port map (
            O => \N__41807\,
            I => \N__41785\
        );

    \I__9391\ : Span4Mux_v
    port map (
            O => \N__41802\,
            I => \N__41780\
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__41799\,
            I => \N__41780\
        );

    \I__9389\ : CascadeMux
    port map (
            O => \N__41798\,
            I => \N__41777\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__41795\,
            I => \N__41774\
        );

    \I__9387\ : Span4Mux_h
    port map (
            O => \N__41790\,
            I => \N__41771\
        );

    \I__9386\ : Span4Mux_h
    port map (
            O => \N__41785\,
            I => \N__41768\
        );

    \I__9385\ : Span4Mux_h
    port map (
            O => \N__41780\,
            I => \N__41765\
        );

    \I__9384\ : InMux
    port map (
            O => \N__41777\,
            I => \N__41762\
        );

    \I__9383\ : Odrv12
    port map (
            O => \N__41774\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__9382\ : Odrv4
    port map (
            O => \N__41771\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__9381\ : Odrv4
    port map (
            O => \N__41768\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__9380\ : Odrv4
    port map (
            O => \N__41765\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__41762\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__9378\ : CEMux
    port map (
            O => \N__41751\,
            I => \N__41736\
        );

    \I__9377\ : CEMux
    port map (
            O => \N__41750\,
            I => \N__41736\
        );

    \I__9376\ : CEMux
    port map (
            O => \N__41749\,
            I => \N__41736\
        );

    \I__9375\ : CEMux
    port map (
            O => \N__41748\,
            I => \N__41736\
        );

    \I__9374\ : CEMux
    port map (
            O => \N__41747\,
            I => \N__41736\
        );

    \I__9373\ : GlobalMux
    port map (
            O => \N__41736\,
            I => \N__41733\
        );

    \I__9372\ : gio2CtrlBuf
    port map (
            O => \N__41733\,
            I => \delay_measurement_inst.delay_hc_timer.N_335_i_g\
        );

    \I__9371\ : InMux
    port map (
            O => \N__41730\,
            I => \N__41727\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__41727\,
            I => \N__41722\
        );

    \I__9369\ : InMux
    port map (
            O => \N__41726\,
            I => \N__41717\
        );

    \I__9368\ : InMux
    port map (
            O => \N__41725\,
            I => \N__41717\
        );

    \I__9367\ : Odrv4
    port map (
            O => \N__41722\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__41717\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__9365\ : InMux
    port map (
            O => \N__41712\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__9364\ : InMux
    port map (
            O => \N__41709\,
            I => \N__41706\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__41706\,
            I => \N__41701\
        );

    \I__9362\ : InMux
    port map (
            O => \N__41705\,
            I => \N__41698\
        );

    \I__9361\ : CascadeMux
    port map (
            O => \N__41704\,
            I => \N__41695\
        );

    \I__9360\ : Span4Mux_h
    port map (
            O => \N__41701\,
            I => \N__41692\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__41698\,
            I => \N__41689\
        );

    \I__9358\ : InMux
    port map (
            O => \N__41695\,
            I => \N__41686\
        );

    \I__9357\ : Odrv4
    port map (
            O => \N__41692\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__9356\ : Odrv4
    port map (
            O => \N__41689\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__41686\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__9354\ : InMux
    port map (
            O => \N__41679\,
            I => \bfn_17_10_0_\
        );

    \I__9353\ : InMux
    port map (
            O => \N__41676\,
            I => \N__41670\
        );

    \I__9352\ : InMux
    port map (
            O => \N__41675\,
            I => \N__41670\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__41670\,
            I => \N__41667\
        );

    \I__9350\ : Odrv4
    port map (
            O => \N__41667\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9349\ : InMux
    port map (
            O => \N__41664\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__9348\ : InMux
    port map (
            O => \N__41661\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__9347\ : InMux
    port map (
            O => \N__41658\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__9346\ : InMux
    port map (
            O => \N__41655\,
            I => \N__41652\
        );

    \I__9345\ : LocalMux
    port map (
            O => \N__41652\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__9344\ : InMux
    port map (
            O => \N__41649\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__9343\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41643\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__41643\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_24\
        );

    \I__9341\ : InMux
    port map (
            O => \N__41640\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__9340\ : InMux
    port map (
            O => \N__41637\,
            I => \N__41634\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__41634\,
            I => \N__41631\
        );

    \I__9338\ : Span4Mux_h
    port map (
            O => \N__41631\,
            I => \N__41627\
        );

    \I__9337\ : InMux
    port map (
            O => \N__41630\,
            I => \N__41624\
        );

    \I__9336\ : Odrv4
    port map (
            O => \N__41627\,
            I => \delay_measurement_inst.elapsed_time_hc_25\
        );

    \I__9335\ : LocalMux
    port map (
            O => \N__41624\,
            I => \delay_measurement_inst.elapsed_time_hc_25\
        );

    \I__9334\ : InMux
    port map (
            O => \N__41619\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__9333\ : InMux
    port map (
            O => \N__41616\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__9332\ : InMux
    port map (
            O => \N__41613\,
            I => \N__41610\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__41610\,
            I => \N__41606\
        );

    \I__9330\ : CascadeMux
    port map (
            O => \N__41609\,
            I => \N__41603\
        );

    \I__9329\ : Span4Mux_h
    port map (
            O => \N__41606\,
            I => \N__41599\
        );

    \I__9328\ : InMux
    port map (
            O => \N__41603\,
            I => \N__41596\
        );

    \I__9327\ : InMux
    port map (
            O => \N__41602\,
            I => \N__41593\
        );

    \I__9326\ : Odrv4
    port map (
            O => \N__41599\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__41596\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__41593\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__9323\ : InMux
    port map (
            O => \N__41586\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__9322\ : InMux
    port map (
            O => \N__41583\,
            I => \N__41580\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__41580\,
            I => \N__41576\
        );

    \I__9320\ : InMux
    port map (
            O => \N__41579\,
            I => \N__41573\
        );

    \I__9319\ : Span4Mux_h
    port map (
            O => \N__41576\,
            I => \N__41569\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__41573\,
            I => \N__41566\
        );

    \I__9317\ : InMux
    port map (
            O => \N__41572\,
            I => \N__41563\
        );

    \I__9316\ : Odrv4
    port map (
            O => \N__41569\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__9315\ : Odrv4
    port map (
            O => \N__41566\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__41563\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__9313\ : InMux
    port map (
            O => \N__41556\,
            I => \bfn_17_9_0_\
        );

    \I__9312\ : InMux
    port map (
            O => \N__41553\,
            I => \N__41550\
        );

    \I__9311\ : LocalMux
    port map (
            O => \N__41550\,
            I => \N__41546\
        );

    \I__9310\ : CascadeMux
    port map (
            O => \N__41549\,
            I => \N__41543\
        );

    \I__9309\ : Span4Mux_h
    port map (
            O => \N__41546\,
            I => \N__41539\
        );

    \I__9308\ : InMux
    port map (
            O => \N__41543\,
            I => \N__41536\
        );

    \I__9307\ : InMux
    port map (
            O => \N__41542\,
            I => \N__41533\
        );

    \I__9306\ : Odrv4
    port map (
            O => \N__41539\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__41536\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__41533\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__9303\ : InMux
    port map (
            O => \N__41526\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__9302\ : InMux
    port map (
            O => \N__41523\,
            I => \N__41519\
        );

    \I__9301\ : CascadeMux
    port map (
            O => \N__41522\,
            I => \N__41515\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__41519\,
            I => \N__41512\
        );

    \I__9299\ : InMux
    port map (
            O => \N__41518\,
            I => \N__41509\
        );

    \I__9298\ : InMux
    port map (
            O => \N__41515\,
            I => \N__41506\
        );

    \I__9297\ : Odrv4
    port map (
            O => \N__41512\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__41509\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__41506\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__9294\ : InMux
    port map (
            O => \N__41499\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__9293\ : InMux
    port map (
            O => \N__41496\,
            I => \N__41493\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__41493\,
            I => \N__41487\
        );

    \I__9291\ : InMux
    port map (
            O => \N__41492\,
            I => \N__41482\
        );

    \I__9290\ : InMux
    port map (
            O => \N__41491\,
            I => \N__41482\
        );

    \I__9289\ : InMux
    port map (
            O => \N__41490\,
            I => \N__41479\
        );

    \I__9288\ : Odrv4
    port map (
            O => \N__41487\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__41482\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__41479\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__9285\ : InMux
    port map (
            O => \N__41472\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__9284\ : InMux
    port map (
            O => \N__41469\,
            I => \N__41466\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__41466\,
            I => \N__41457\
        );

    \I__9282\ : InMux
    port map (
            O => \N__41465\,
            I => \N__41450\
        );

    \I__9281\ : InMux
    port map (
            O => \N__41464\,
            I => \N__41450\
        );

    \I__9280\ : InMux
    port map (
            O => \N__41463\,
            I => \N__41450\
        );

    \I__9279\ : InMux
    port map (
            O => \N__41462\,
            I => \N__41443\
        );

    \I__9278\ : InMux
    port map (
            O => \N__41461\,
            I => \N__41443\
        );

    \I__9277\ : InMux
    port map (
            O => \N__41460\,
            I => \N__41443\
        );

    \I__9276\ : Odrv4
    port map (
            O => \N__41457\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__41450\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__9274\ : LocalMux
    port map (
            O => \N__41443\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__9273\ : InMux
    port map (
            O => \N__41436\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__9272\ : InMux
    port map (
            O => \N__41433\,
            I => \N__41430\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__41430\,
            I => \N__41425\
        );

    \I__9270\ : InMux
    port map (
            O => \N__41429\,
            I => \N__41422\
        );

    \I__9269\ : InMux
    port map (
            O => \N__41428\,
            I => \N__41419\
        );

    \I__9268\ : Odrv4
    port map (
            O => \N__41425\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__41422\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__41419\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__9265\ : InMux
    port map (
            O => \N__41412\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__9264\ : InMux
    port map (
            O => \N__41409\,
            I => \N__41406\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__41406\,
            I => \N__41401\
        );

    \I__9262\ : InMux
    port map (
            O => \N__41405\,
            I => \N__41396\
        );

    \I__9261\ : InMux
    port map (
            O => \N__41404\,
            I => \N__41396\
        );

    \I__9260\ : Odrv4
    port map (
            O => \N__41401\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__41396\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__9258\ : InMux
    port map (
            O => \N__41391\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__9257\ : CascadeMux
    port map (
            O => \N__41388\,
            I => \N__41385\
        );

    \I__9256\ : InMux
    port map (
            O => \N__41385\,
            I => \N__41382\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__41382\,
            I => \N__41379\
        );

    \I__9254\ : Span4Mux_v
    port map (
            O => \N__41379\,
            I => \N__41375\
        );

    \I__9253\ : InMux
    port map (
            O => \N__41378\,
            I => \N__41372\
        );

    \I__9252\ : Odrv4
    port map (
            O => \N__41375\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__41372\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__9250\ : CascadeMux
    port map (
            O => \N__41367\,
            I => \N__41364\
        );

    \I__9249\ : InMux
    port map (
            O => \N__41364\,
            I => \N__41359\
        );

    \I__9248\ : InMux
    port map (
            O => \N__41363\,
            I => \N__41356\
        );

    \I__9247\ : InMux
    port map (
            O => \N__41362\,
            I => \N__41353\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__41359\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__41356\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__41353\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__9243\ : CascadeMux
    port map (
            O => \N__41346\,
            I => \N__41343\
        );

    \I__9242\ : InMux
    port map (
            O => \N__41343\,
            I => \N__41340\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__41340\,
            I => \N__41337\
        );

    \I__9240\ : Span4Mux_h
    port map (
            O => \N__41337\,
            I => \N__41332\
        );

    \I__9239\ : InMux
    port map (
            O => \N__41336\,
            I => \N__41329\
        );

    \I__9238\ : InMux
    port map (
            O => \N__41335\,
            I => \N__41326\
        );

    \I__9237\ : Odrv4
    port map (
            O => \N__41332\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__9236\ : LocalMux
    port map (
            O => \N__41329\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__41326\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__9234\ : CascadeMux
    port map (
            O => \N__41319\,
            I => \N__41316\
        );

    \I__9233\ : InMux
    port map (
            O => \N__41316\,
            I => \N__41313\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__41313\,
            I => \N__41309\
        );

    \I__9231\ : CascadeMux
    port map (
            O => \N__41312\,
            I => \N__41306\
        );

    \I__9230\ : Span4Mux_h
    port map (
            O => \N__41309\,
            I => \N__41302\
        );

    \I__9229\ : InMux
    port map (
            O => \N__41306\,
            I => \N__41297\
        );

    \I__9228\ : InMux
    port map (
            O => \N__41305\,
            I => \N__41297\
        );

    \I__9227\ : Odrv4
    port map (
            O => \N__41302\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__41297\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__9225\ : InMux
    port map (
            O => \N__41292\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__9224\ : InMux
    port map (
            O => \N__41289\,
            I => \N__41286\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__41286\,
            I => \N__41282\
        );

    \I__9222\ : CascadeMux
    port map (
            O => \N__41285\,
            I => \N__41278\
        );

    \I__9221\ : Span4Mux_h
    port map (
            O => \N__41282\,
            I => \N__41275\
        );

    \I__9220\ : InMux
    port map (
            O => \N__41281\,
            I => \N__41272\
        );

    \I__9219\ : InMux
    port map (
            O => \N__41278\,
            I => \N__41269\
        );

    \I__9218\ : Odrv4
    port map (
            O => \N__41275\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__41272\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__9216\ : LocalMux
    port map (
            O => \N__41269\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__9215\ : InMux
    port map (
            O => \N__41262\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__9214\ : InMux
    port map (
            O => \N__41259\,
            I => \N__41254\
        );

    \I__9213\ : CascadeMux
    port map (
            O => \N__41258\,
            I => \N__41251\
        );

    \I__9212\ : CascadeMux
    port map (
            O => \N__41257\,
            I => \N__41247\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__41254\,
            I => \N__41244\
        );

    \I__9210\ : InMux
    port map (
            O => \N__41251\,
            I => \N__41239\
        );

    \I__9209\ : InMux
    port map (
            O => \N__41250\,
            I => \N__41239\
        );

    \I__9208\ : InMux
    port map (
            O => \N__41247\,
            I => \N__41236\
        );

    \I__9207\ : Span4Mux_h
    port map (
            O => \N__41244\,
            I => \N__41233\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__41239\,
            I => \N__41228\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__41236\,
            I => \N__41228\
        );

    \I__9204\ : Odrv4
    port map (
            O => \N__41233\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__9203\ : Odrv4
    port map (
            O => \N__41228\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__9202\ : InMux
    port map (
            O => \N__41223\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__9201\ : InMux
    port map (
            O => \N__41220\,
            I => \N__41217\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__41217\,
            I => \N__41214\
        );

    \I__9199\ : Span4Mux_h
    port map (
            O => \N__41214\,
            I => \N__41207\
        );

    \I__9198\ : InMux
    port map (
            O => \N__41213\,
            I => \N__41200\
        );

    \I__9197\ : InMux
    port map (
            O => \N__41212\,
            I => \N__41200\
        );

    \I__9196\ : InMux
    port map (
            O => \N__41211\,
            I => \N__41200\
        );

    \I__9195\ : InMux
    port map (
            O => \N__41210\,
            I => \N__41197\
        );

    \I__9194\ : Odrv4
    port map (
            O => \N__41207\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__9193\ : LocalMux
    port map (
            O => \N__41200\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__41197\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__9191\ : InMux
    port map (
            O => \N__41190\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__9190\ : InMux
    port map (
            O => \N__41187\,
            I => \N__41183\
        );

    \I__9189\ : CascadeMux
    port map (
            O => \N__41186\,
            I => \N__41177\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__41183\,
            I => \N__41174\
        );

    \I__9187\ : InMux
    port map (
            O => \N__41182\,
            I => \N__41167\
        );

    \I__9186\ : InMux
    port map (
            O => \N__41181\,
            I => \N__41167\
        );

    \I__9185\ : InMux
    port map (
            O => \N__41180\,
            I => \N__41167\
        );

    \I__9184\ : InMux
    port map (
            O => \N__41177\,
            I => \N__41164\
        );

    \I__9183\ : Odrv4
    port map (
            O => \N__41174\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__41167\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__41164\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__9180\ : InMux
    port map (
            O => \N__41157\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__9179\ : InMux
    port map (
            O => \N__41154\,
            I => \N__41151\
        );

    \I__9178\ : LocalMux
    port map (
            O => \N__41151\,
            I => \N__41146\
        );

    \I__9177\ : CascadeMux
    port map (
            O => \N__41150\,
            I => \N__41142\
        );

    \I__9176\ : CascadeMux
    port map (
            O => \N__41149\,
            I => \N__41139\
        );

    \I__9175\ : Span4Mux_h
    port map (
            O => \N__41146\,
            I => \N__41136\
        );

    \I__9174\ : InMux
    port map (
            O => \N__41145\,
            I => \N__41133\
        );

    \I__9173\ : InMux
    port map (
            O => \N__41142\,
            I => \N__41130\
        );

    \I__9172\ : InMux
    port map (
            O => \N__41139\,
            I => \N__41127\
        );

    \I__9171\ : Odrv4
    port map (
            O => \N__41136\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__41133\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__41130\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__41127\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__9167\ : InMux
    port map (
            O => \N__41118\,
            I => \N__41115\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__41115\,
            I => \N__41111\
        );

    \I__9165\ : InMux
    port map (
            O => \N__41114\,
            I => \N__41108\
        );

    \I__9164\ : Span4Mux_v
    port map (
            O => \N__41111\,
            I => \N__41105\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__41108\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9162\ : Odrv4
    port map (
            O => \N__41105\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9161\ : InMux
    port map (
            O => \N__41100\,
            I => \N__41097\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__41097\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_19\
        );

    \I__9159\ : InMux
    port map (
            O => \N__41094\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__9158\ : InMux
    port map (
            O => \N__41091\,
            I => \N__41086\
        );

    \I__9157\ : InMux
    port map (
            O => \N__41090\,
            I => \N__41081\
        );

    \I__9156\ : InMux
    port map (
            O => \N__41089\,
            I => \N__41081\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__41086\,
            I => \N__41078\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__41081\,
            I => \N__41075\
        );

    \I__9153\ : Span4Mux_h
    port map (
            O => \N__41078\,
            I => \N__41069\
        );

    \I__9152\ : Span4Mux_v
    port map (
            O => \N__41075\,
            I => \N__41066\
        );

    \I__9151\ : InMux
    port map (
            O => \N__41074\,
            I => \N__41063\
        );

    \I__9150\ : InMux
    port map (
            O => \N__41073\,
            I => \N__41058\
        );

    \I__9149\ : InMux
    port map (
            O => \N__41072\,
            I => \N__41058\
        );

    \I__9148\ : Span4Mux_v
    port map (
            O => \N__41069\,
            I => \N__41055\
        );

    \I__9147\ : Span4Mux_h
    port map (
            O => \N__41066\,
            I => \N__41050\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__41063\,
            I => \N__41050\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__41058\,
            I => \N__41047\
        );

    \I__9144\ : Odrv4
    port map (
            O => \N__41055\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9143\ : Odrv4
    port map (
            O => \N__41050\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9142\ : Odrv12
    port map (
            O => \N__41047\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9141\ : CascadeMux
    port map (
            O => \N__41040\,
            I => \N__41037\
        );

    \I__9140\ : InMux
    port map (
            O => \N__41037\,
            I => \N__41034\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__41034\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\
        );

    \I__9138\ : CascadeMux
    port map (
            O => \N__41031\,
            I => \N__41028\
        );

    \I__9137\ : InMux
    port map (
            O => \N__41028\,
            I => \N__41025\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__41025\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\
        );

    \I__9135\ : CascadeMux
    port map (
            O => \N__41022\,
            I => \N__41019\
        );

    \I__9134\ : InMux
    port map (
            O => \N__41019\,
            I => \N__41016\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__41016\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\
        );

    \I__9132\ : InMux
    port map (
            O => \N__41013\,
            I => \N__41010\
        );

    \I__9131\ : LocalMux
    port map (
            O => \N__41010\,
            I => \N__41007\
        );

    \I__9130\ : Odrv4
    port map (
            O => \N__41007\,
            I => delay_hc_input_c
        );

    \I__9129\ : InMux
    port map (
            O => \N__41004\,
            I => \N__41001\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__41001\,
            I => \N__40998\
        );

    \I__9127\ : Span4Mux_h
    port map (
            O => \N__40998\,
            I => \N__40995\
        );

    \I__9126\ : Span4Mux_v
    port map (
            O => \N__40995\,
            I => \N__40992\
        );

    \I__9125\ : Odrv4
    port map (
            O => \N__40992\,
            I => delay_hc_d1
        );

    \I__9124\ : InMux
    port map (
            O => \N__40989\,
            I => \N__40985\
        );

    \I__9123\ : InMux
    port map (
            O => \N__40988\,
            I => \N__40982\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__40985\,
            I => \N__40979\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__40982\,
            I => \N__40976\
        );

    \I__9120\ : Span4Mux_v
    port map (
            O => \N__40979\,
            I => \N__40973\
        );

    \I__9119\ : Span4Mux_v
    port map (
            O => \N__40976\,
            I => \N__40970\
        );

    \I__9118\ : Span4Mux_v
    port map (
            O => \N__40973\,
            I => \N__40967\
        );

    \I__9117\ : Span4Mux_h
    port map (
            O => \N__40970\,
            I => \N__40964\
        );

    \I__9116\ : Odrv4
    port map (
            O => \N__40967\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__9115\ : Odrv4
    port map (
            O => \N__40964\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__9114\ : InMux
    port map (
            O => \N__40959\,
            I => \N__40955\
        );

    \I__9113\ : InMux
    port map (
            O => \N__40958\,
            I => \N__40951\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__40955\,
            I => \N__40948\
        );

    \I__9111\ : InMux
    port map (
            O => \N__40954\,
            I => \N__40945\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__40951\,
            I => \N__40940\
        );

    \I__9109\ : Span4Mux_h
    port map (
            O => \N__40948\,
            I => \N__40940\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__40945\,
            I => \N__40937\
        );

    \I__9107\ : Span4Mux_v
    port map (
            O => \N__40940\,
            I => \N__40934\
        );

    \I__9106\ : Span4Mux_h
    port map (
            O => \N__40937\,
            I => \N__40931\
        );

    \I__9105\ : Span4Mux_h
    port map (
            O => \N__40934\,
            I => \N__40928\
        );

    \I__9104\ : Span4Mux_v
    port map (
            O => \N__40931\,
            I => \N__40925\
        );

    \I__9103\ : Odrv4
    port map (
            O => \N__40928\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__9102\ : Odrv4
    port map (
            O => \N__40925\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__9101\ : InMux
    port map (
            O => \N__40920\,
            I => \N__40917\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__40917\,
            I => \N__40913\
        );

    \I__9099\ : InMux
    port map (
            O => \N__40916\,
            I => \N__40908\
        );

    \I__9098\ : Span4Mux_h
    port map (
            O => \N__40913\,
            I => \N__40905\
        );

    \I__9097\ : InMux
    port map (
            O => \N__40912\,
            I => \N__40900\
        );

    \I__9096\ : InMux
    port map (
            O => \N__40911\,
            I => \N__40900\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__40908\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__9094\ : Odrv4
    port map (
            O => \N__40905\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__40900\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__9092\ : InMux
    port map (
            O => \N__40893\,
            I => \N__40890\
        );

    \I__9091\ : LocalMux
    port map (
            O => \N__40890\,
            I => \N__40887\
        );

    \I__9090\ : Span4Mux_v
    port map (
            O => \N__40887\,
            I => \N__40882\
        );

    \I__9089\ : InMux
    port map (
            O => \N__40886\,
            I => \N__40879\
        );

    \I__9088\ : InMux
    port map (
            O => \N__40885\,
            I => \N__40874\
        );

    \I__9087\ : Span4Mux_h
    port map (
            O => \N__40882\,
            I => \N__40871\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__40879\,
            I => \N__40868\
        );

    \I__9085\ : InMux
    port map (
            O => \N__40878\,
            I => \N__40865\
        );

    \I__9084\ : InMux
    port map (
            O => \N__40877\,
            I => \N__40862\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__40874\,
            I => \N__40859\
        );

    \I__9082\ : Span4Mux_h
    port map (
            O => \N__40871\,
            I => \N__40854\
        );

    \I__9081\ : Span4Mux_v
    port map (
            O => \N__40868\,
            I => \N__40854\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__40865\,
            I => \N__40851\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__40862\,
            I => \N__40844\
        );

    \I__9078\ : Span4Mux_v
    port map (
            O => \N__40859\,
            I => \N__40844\
        );

    \I__9077\ : Span4Mux_h
    port map (
            O => \N__40854\,
            I => \N__40844\
        );

    \I__9076\ : Span4Mux_h
    port map (
            O => \N__40851\,
            I => \N__40841\
        );

    \I__9075\ : Odrv4
    port map (
            O => \N__40844\,
            I => measured_delay_hc_2
        );

    \I__9074\ : Odrv4
    port map (
            O => \N__40841\,
            I => measured_delay_hc_2
        );

    \I__9073\ : InMux
    port map (
            O => \N__40836\,
            I => \N__40829\
        );

    \I__9072\ : InMux
    port map (
            O => \N__40835\,
            I => \N__40824\
        );

    \I__9071\ : InMux
    port map (
            O => \N__40834\,
            I => \N__40824\
        );

    \I__9070\ : CascadeMux
    port map (
            O => \N__40833\,
            I => \N__40815\
        );

    \I__9069\ : CascadeMux
    port map (
            O => \N__40832\,
            I => \N__40812\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__40829\,
            I => \N__40803\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__40824\,
            I => \N__40803\
        );

    \I__9066\ : InMux
    port map (
            O => \N__40823\,
            I => \N__40795\
        );

    \I__9065\ : InMux
    port map (
            O => \N__40822\,
            I => \N__40792\
        );

    \I__9064\ : InMux
    port map (
            O => \N__40821\,
            I => \N__40787\
        );

    \I__9063\ : InMux
    port map (
            O => \N__40820\,
            I => \N__40787\
        );

    \I__9062\ : CascadeMux
    port map (
            O => \N__40819\,
            I => \N__40781\
        );

    \I__9061\ : CascadeMux
    port map (
            O => \N__40818\,
            I => \N__40778\
        );

    \I__9060\ : InMux
    port map (
            O => \N__40815\,
            I => \N__40770\
        );

    \I__9059\ : InMux
    port map (
            O => \N__40812\,
            I => \N__40770\
        );

    \I__9058\ : InMux
    port map (
            O => \N__40811\,
            I => \N__40763\
        );

    \I__9057\ : InMux
    port map (
            O => \N__40810\,
            I => \N__40763\
        );

    \I__9056\ : InMux
    port map (
            O => \N__40809\,
            I => \N__40763\
        );

    \I__9055\ : InMux
    port map (
            O => \N__40808\,
            I => \N__40760\
        );

    \I__9054\ : Span4Mux_h
    port map (
            O => \N__40803\,
            I => \N__40756\
        );

    \I__9053\ : InMux
    port map (
            O => \N__40802\,
            I => \N__40753\
        );

    \I__9052\ : InMux
    port map (
            O => \N__40801\,
            I => \N__40750\
        );

    \I__9051\ : InMux
    port map (
            O => \N__40800\,
            I => \N__40745\
        );

    \I__9050\ : InMux
    port map (
            O => \N__40799\,
            I => \N__40745\
        );

    \I__9049\ : InMux
    port map (
            O => \N__40798\,
            I => \N__40737\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__40795\,
            I => \N__40730\
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__40792\,
            I => \N__40730\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__40787\,
            I => \N__40730\
        );

    \I__9045\ : InMux
    port map (
            O => \N__40786\,
            I => \N__40723\
        );

    \I__9044\ : InMux
    port map (
            O => \N__40785\,
            I => \N__40723\
        );

    \I__9043\ : InMux
    port map (
            O => \N__40784\,
            I => \N__40723\
        );

    \I__9042\ : InMux
    port map (
            O => \N__40781\,
            I => \N__40716\
        );

    \I__9041\ : InMux
    port map (
            O => \N__40778\,
            I => \N__40716\
        );

    \I__9040\ : InMux
    port map (
            O => \N__40777\,
            I => \N__40716\
        );

    \I__9039\ : InMux
    port map (
            O => \N__40776\,
            I => \N__40711\
        );

    \I__9038\ : InMux
    port map (
            O => \N__40775\,
            I => \N__40711\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__40770\,
            I => \N__40706\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__40763\,
            I => \N__40706\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__40760\,
            I => \N__40703\
        );

    \I__9034\ : InMux
    port map (
            O => \N__40759\,
            I => \N__40700\
        );

    \I__9033\ : Sp12to4
    port map (
            O => \N__40756\,
            I => \N__40691\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__40753\,
            I => \N__40691\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__40750\,
            I => \N__40691\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__40745\,
            I => \N__40691\
        );

    \I__9029\ : InMux
    port map (
            O => \N__40744\,
            I => \N__40684\
        );

    \I__9028\ : InMux
    port map (
            O => \N__40743\,
            I => \N__40684\
        );

    \I__9027\ : InMux
    port map (
            O => \N__40742\,
            I => \N__40684\
        );

    \I__9026\ : InMux
    port map (
            O => \N__40741\,
            I => \N__40679\
        );

    \I__9025\ : InMux
    port map (
            O => \N__40740\,
            I => \N__40679\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__40737\,
            I => \N__40674\
        );

    \I__9023\ : Span4Mux_v
    port map (
            O => \N__40730\,
            I => \N__40674\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__40723\,
            I => \N__40665\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__40716\,
            I => \N__40665\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__40711\,
            I => \N__40665\
        );

    \I__9019\ : Span4Mux_h
    port map (
            O => \N__40706\,
            I => \N__40665\
        );

    \I__9018\ : Span4Mux_h
    port map (
            O => \N__40703\,
            I => \N__40662\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__40700\,
            I => \N__40657\
        );

    \I__9016\ : Span12Mux_v
    port map (
            O => \N__40691\,
            I => \N__40657\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__40684\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__40679\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__9013\ : Odrv4
    port map (
            O => \N__40674\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__9012\ : Odrv4
    port map (
            O => \N__40665\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__9011\ : Odrv4
    port map (
            O => \N__40662\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__9010\ : Odrv12
    port map (
            O => \N__40657\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__9009\ : InMux
    port map (
            O => \N__40644\,
            I => \N__40641\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__40641\,
            I => \N__40636\
        );

    \I__9007\ : InMux
    port map (
            O => \N__40640\,
            I => \N__40631\
        );

    \I__9006\ : InMux
    port map (
            O => \N__40639\,
            I => \N__40631\
        );

    \I__9005\ : Span4Mux_h
    port map (
            O => \N__40636\,
            I => \N__40614\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__40631\,
            I => \N__40611\
        );

    \I__9003\ : InMux
    port map (
            O => \N__40630\,
            I => \N__40604\
        );

    \I__9002\ : InMux
    port map (
            O => \N__40629\,
            I => \N__40604\
        );

    \I__9001\ : InMux
    port map (
            O => \N__40628\,
            I => \N__40604\
        );

    \I__9000\ : InMux
    port map (
            O => \N__40627\,
            I => \N__40593\
        );

    \I__8999\ : InMux
    port map (
            O => \N__40626\,
            I => \N__40593\
        );

    \I__8998\ : InMux
    port map (
            O => \N__40625\,
            I => \N__40593\
        );

    \I__8997\ : InMux
    port map (
            O => \N__40624\,
            I => \N__40593\
        );

    \I__8996\ : InMux
    port map (
            O => \N__40623\,
            I => \N__40593\
        );

    \I__8995\ : InMux
    port map (
            O => \N__40622\,
            I => \N__40590\
        );

    \I__8994\ : InMux
    port map (
            O => \N__40621\,
            I => \N__40585\
        );

    \I__8993\ : InMux
    port map (
            O => \N__40620\,
            I => \N__40585\
        );

    \I__8992\ : InMux
    port map (
            O => \N__40619\,
            I => \N__40578\
        );

    \I__8991\ : InMux
    port map (
            O => \N__40618\,
            I => \N__40578\
        );

    \I__8990\ : InMux
    port map (
            O => \N__40617\,
            I => \N__40578\
        );

    \I__8989\ : Odrv4
    port map (
            O => \N__40614\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__8988\ : Odrv4
    port map (
            O => \N__40611\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__40604\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__40593\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__40590\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__40585\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__40578\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__8982\ : CascadeMux
    port map (
            O => \N__40563\,
            I => \N__40559\
        );

    \I__8981\ : CascadeMux
    port map (
            O => \N__40562\,
            I => \N__40556\
        );

    \I__8980\ : InMux
    port map (
            O => \N__40559\,
            I => \N__40551\
        );

    \I__8979\ : InMux
    port map (
            O => \N__40556\,
            I => \N__40548\
        );

    \I__8978\ : InMux
    port map (
            O => \N__40555\,
            I => \N__40545\
        );

    \I__8977\ : InMux
    port map (
            O => \N__40554\,
            I => \N__40542\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__40551\,
            I => \N__40537\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__40548\,
            I => \N__40534\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__40545\,
            I => \N__40531\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__40542\,
            I => \N__40528\
        );

    \I__8972\ : InMux
    port map (
            O => \N__40541\,
            I => \N__40525\
        );

    \I__8971\ : CascadeMux
    port map (
            O => \N__40540\,
            I => \N__40522\
        );

    \I__8970\ : Span4Mux_v
    port map (
            O => \N__40537\,
            I => \N__40519\
        );

    \I__8969\ : Span4Mux_v
    port map (
            O => \N__40534\,
            I => \N__40514\
        );

    \I__8968\ : Span4Mux_h
    port map (
            O => \N__40531\,
            I => \N__40514\
        );

    \I__8967\ : Span4Mux_h
    port map (
            O => \N__40528\,
            I => \N__40511\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__40525\,
            I => \N__40508\
        );

    \I__8965\ : InMux
    port map (
            O => \N__40522\,
            I => \N__40505\
        );

    \I__8964\ : Span4Mux_h
    port map (
            O => \N__40519\,
            I => \N__40500\
        );

    \I__8963\ : Span4Mux_v
    port map (
            O => \N__40514\,
            I => \N__40500\
        );

    \I__8962\ : Span4Mux_h
    port map (
            O => \N__40511\,
            I => \N__40497\
        );

    \I__8961\ : Span12Mux_h
    port map (
            O => \N__40508\,
            I => \N__40494\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__40505\,
            I => measured_delay_hc_15
        );

    \I__8959\ : Odrv4
    port map (
            O => \N__40500\,
            I => measured_delay_hc_15
        );

    \I__8958\ : Odrv4
    port map (
            O => \N__40497\,
            I => measured_delay_hc_15
        );

    \I__8957\ : Odrv12
    port map (
            O => \N__40494\,
            I => measured_delay_hc_15
        );

    \I__8956\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40481\
        );

    \I__8955\ : InMux
    port map (
            O => \N__40484\,
            I => \N__40478\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__40481\,
            I => \N__40475\
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__40478\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8952\ : Odrv12
    port map (
            O => \N__40475\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8951\ : InMux
    port map (
            O => \N__40470\,
            I => \N__40467\
        );

    \I__8950\ : LocalMux
    port map (
            O => \N__40467\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_12\
        );

    \I__8949\ : InMux
    port map (
            O => \N__40464\,
            I => \N__40460\
        );

    \I__8948\ : InMux
    port map (
            O => \N__40463\,
            I => \N__40457\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__40460\,
            I => \N__40454\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__40457\,
            I => \N__40451\
        );

    \I__8945\ : Odrv4
    port map (
            O => \N__40454\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8944\ : Odrv4
    port map (
            O => \N__40451\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8943\ : InMux
    port map (
            O => \N__40446\,
            I => \N__40443\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__40443\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_13\
        );

    \I__8941\ : CascadeMux
    port map (
            O => \N__40440\,
            I => \N__40437\
        );

    \I__8940\ : InMux
    port map (
            O => \N__40437\,
            I => \N__40434\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__40434\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\
        );

    \I__8938\ : InMux
    port map (
            O => \N__40431\,
            I => \N__40428\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__40428\,
            I => \N__40424\
        );

    \I__8936\ : InMux
    port map (
            O => \N__40427\,
            I => \N__40421\
        );

    \I__8935\ : Span4Mux_v
    port map (
            O => \N__40424\,
            I => \N__40416\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__40421\,
            I => \N__40416\
        );

    \I__8933\ : Odrv4
    port map (
            O => \N__40416\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8932\ : InMux
    port map (
            O => \N__40413\,
            I => \N__40410\
        );

    \I__8931\ : LocalMux
    port map (
            O => \N__40410\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_14\
        );

    \I__8930\ : CascadeMux
    port map (
            O => \N__40407\,
            I => \N__40404\
        );

    \I__8929\ : InMux
    port map (
            O => \N__40404\,
            I => \N__40401\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__40401\,
            I => \N__40398\
        );

    \I__8927\ : Odrv4
    port map (
            O => \N__40398\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\
        );

    \I__8926\ : InMux
    port map (
            O => \N__40395\,
            I => \N__40392\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__40392\,
            I => \N__40388\
        );

    \I__8924\ : InMux
    port map (
            O => \N__40391\,
            I => \N__40385\
        );

    \I__8923\ : Span4Mux_v
    port map (
            O => \N__40388\,
            I => \N__40380\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__40385\,
            I => \N__40380\
        );

    \I__8921\ : Odrv4
    port map (
            O => \N__40380\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8920\ : InMux
    port map (
            O => \N__40377\,
            I => \N__40374\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__40374\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_15\
        );

    \I__8918\ : InMux
    port map (
            O => \N__40371\,
            I => \N__40368\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__40368\,
            I => \N__40364\
        );

    \I__8916\ : InMux
    port map (
            O => \N__40367\,
            I => \N__40361\
        );

    \I__8915\ : Span4Mux_v
    port map (
            O => \N__40364\,
            I => \N__40358\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__40361\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8913\ : Odrv4
    port map (
            O => \N__40358\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8912\ : CascadeMux
    port map (
            O => \N__40353\,
            I => \N__40350\
        );

    \I__8911\ : InMux
    port map (
            O => \N__40350\,
            I => \N__40347\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__40347\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_16\
        );

    \I__8909\ : InMux
    port map (
            O => \N__40344\,
            I => \N__40341\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__40341\,
            I => \N__40337\
        );

    \I__8907\ : InMux
    port map (
            O => \N__40340\,
            I => \N__40334\
        );

    \I__8906\ : Span4Mux_v
    port map (
            O => \N__40337\,
            I => \N__40331\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__40334\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8904\ : Odrv4
    port map (
            O => \N__40331\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8903\ : InMux
    port map (
            O => \N__40326\,
            I => \N__40323\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__40323\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_17\
        );

    \I__8901\ : InMux
    port map (
            O => \N__40320\,
            I => \N__40317\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__40317\,
            I => \N__40313\
        );

    \I__8899\ : InMux
    port map (
            O => \N__40316\,
            I => \N__40310\
        );

    \I__8898\ : Span4Mux_v
    port map (
            O => \N__40313\,
            I => \N__40307\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__40310\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8896\ : Odrv4
    port map (
            O => \N__40307\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8895\ : InMux
    port map (
            O => \N__40302\,
            I => \N__40299\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__40299\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_18\
        );

    \I__8893\ : InMux
    port map (
            O => \N__40296\,
            I => \N__40292\
        );

    \I__8892\ : InMux
    port map (
            O => \N__40295\,
            I => \N__40289\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__40292\,
            I => \N__40286\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__40289\,
            I => \N__40283\
        );

    \I__8889\ : Odrv4
    port map (
            O => \N__40286\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8888\ : Odrv4
    port map (
            O => \N__40283\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8887\ : InMux
    port map (
            O => \N__40278\,
            I => \N__40275\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__40275\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_4\
        );

    \I__8885\ : CascadeMux
    port map (
            O => \N__40272\,
            I => \N__40269\
        );

    \I__8884\ : InMux
    port map (
            O => \N__40269\,
            I => \N__40266\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__40266\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\
        );

    \I__8882\ : InMux
    port map (
            O => \N__40263\,
            I => \N__40260\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__40260\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_5\
        );

    \I__8880\ : InMux
    port map (
            O => \N__40257\,
            I => \N__40254\
        );

    \I__8879\ : LocalMux
    port map (
            O => \N__40254\,
            I => \N__40250\
        );

    \I__8878\ : InMux
    port map (
            O => \N__40253\,
            I => \N__40247\
        );

    \I__8877\ : Span4Mux_v
    port map (
            O => \N__40250\,
            I => \N__40242\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__40247\,
            I => \N__40242\
        );

    \I__8875\ : Odrv4
    port map (
            O => \N__40242\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8874\ : InMux
    port map (
            O => \N__40239\,
            I => \N__40236\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__40236\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_6\
        );

    \I__8872\ : InMux
    port map (
            O => \N__40233\,
            I => \N__40229\
        );

    \I__8871\ : InMux
    port map (
            O => \N__40232\,
            I => \N__40226\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__40229\,
            I => \N__40223\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__40226\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8868\ : Odrv12
    port map (
            O => \N__40223\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8867\ : InMux
    port map (
            O => \N__40218\,
            I => \N__40215\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__40215\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_7\
        );

    \I__8865\ : CascadeMux
    port map (
            O => \N__40212\,
            I => \N__40209\
        );

    \I__8864\ : InMux
    port map (
            O => \N__40209\,
            I => \N__40206\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__40206\,
            I => \N__40203\
        );

    \I__8862\ : Odrv4
    port map (
            O => \N__40203\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\
        );

    \I__8861\ : InMux
    port map (
            O => \N__40200\,
            I => \N__40197\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__40197\,
            I => \N__40193\
        );

    \I__8859\ : InMux
    port map (
            O => \N__40196\,
            I => \N__40190\
        );

    \I__8858\ : Span4Mux_v
    port map (
            O => \N__40193\,
            I => \N__40187\
        );

    \I__8857\ : LocalMux
    port map (
            O => \N__40190\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8856\ : Odrv4
    port map (
            O => \N__40187\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8855\ : InMux
    port map (
            O => \N__40182\,
            I => \N__40179\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__40179\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_8\
        );

    \I__8853\ : InMux
    port map (
            O => \N__40176\,
            I => \N__40172\
        );

    \I__8852\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40169\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__40172\,
            I => \N__40166\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__40169\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8849\ : Odrv12
    port map (
            O => \N__40166\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8848\ : InMux
    port map (
            O => \N__40161\,
            I => \N__40158\
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__40158\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_9\
        );

    \I__8846\ : InMux
    port map (
            O => \N__40155\,
            I => \N__40151\
        );

    \I__8845\ : InMux
    port map (
            O => \N__40154\,
            I => \N__40148\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__40151\,
            I => \N__40145\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__40148\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8842\ : Odrv12
    port map (
            O => \N__40145\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8841\ : InMux
    port map (
            O => \N__40140\,
            I => \N__40137\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__40137\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_10\
        );

    \I__8839\ : InMux
    port map (
            O => \N__40134\,
            I => \N__40130\
        );

    \I__8838\ : InMux
    port map (
            O => \N__40133\,
            I => \N__40127\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__40130\,
            I => \N__40124\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__40127\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8835\ : Odrv12
    port map (
            O => \N__40124\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8834\ : InMux
    port map (
            O => \N__40119\,
            I => \N__40116\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__40116\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_11\
        );

    \I__8832\ : InMux
    port map (
            O => \N__40113\,
            I => \N__40109\
        );

    \I__8831\ : InMux
    port map (
            O => \N__40112\,
            I => \N__40106\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__40109\,
            I => \N__40103\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__40106\,
            I => \N__40099\
        );

    \I__8828\ : Span4Mux_h
    port map (
            O => \N__40103\,
            I => \N__40096\
        );

    \I__8827\ : InMux
    port map (
            O => \N__40102\,
            I => \N__40093\
        );

    \I__8826\ : Span4Mux_h
    port map (
            O => \N__40099\,
            I => \N__40090\
        );

    \I__8825\ : Odrv4
    port map (
            O => \N__40096\,
            I => measured_delay_tr_2
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__40093\,
            I => measured_delay_tr_2
        );

    \I__8823\ : Odrv4
    port map (
            O => \N__40090\,
            I => measured_delay_tr_2
        );

    \I__8822\ : InMux
    port map (
            O => \N__40083\,
            I => \N__40080\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__40080\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\
        );

    \I__8820\ : InMux
    port map (
            O => \N__40077\,
            I => \N__40074\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__40074\,
            I => \N__40070\
        );

    \I__8818\ : CascadeMux
    port map (
            O => \N__40073\,
            I => \N__40067\
        );

    \I__8817\ : Span4Mux_h
    port map (
            O => \N__40070\,
            I => \N__40064\
        );

    \I__8816\ : InMux
    port map (
            O => \N__40067\,
            I => \N__40061\
        );

    \I__8815\ : Odrv4
    port map (
            O => \N__40064\,
            I => measured_delay_tr_1
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__40061\,
            I => measured_delay_tr_1
        );

    \I__8813\ : CascadeMux
    port map (
            O => \N__40056\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1_cascade_\
        );

    \I__8812\ : InMux
    port map (
            O => \N__40053\,
            I => \N__40050\
        );

    \I__8811\ : LocalMux
    port map (
            O => \N__40050\,
            I => \N__40042\
        );

    \I__8810\ : InMux
    port map (
            O => \N__40049\,
            I => \N__40037\
        );

    \I__8809\ : InMux
    port map (
            O => \N__40048\,
            I => \N__40037\
        );

    \I__8808\ : InMux
    port map (
            O => \N__40047\,
            I => \N__40030\
        );

    \I__8807\ : InMux
    port map (
            O => \N__40046\,
            I => \N__40030\
        );

    \I__8806\ : InMux
    port map (
            O => \N__40045\,
            I => \N__40030\
        );

    \I__8805\ : Span4Mux_v
    port map (
            O => \N__40042\,
            I => \N__40025\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__40037\,
            I => \N__40025\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__40030\,
            I => \phase_controller_inst1.stoper_tr.N_20_li\
        );

    \I__8802\ : Odrv4
    port map (
            O => \N__40025\,
            I => \phase_controller_inst1.stoper_tr.N_20_li\
        );

    \I__8801\ : CascadeMux
    port map (
            O => \N__40020\,
            I => \N__40016\
        );

    \I__8800\ : CascadeMux
    port map (
            O => \N__40019\,
            I => \N__40011\
        );

    \I__8799\ : InMux
    port map (
            O => \N__40016\,
            I => \N__40007\
        );

    \I__8798\ : InMux
    port map (
            O => \N__40015\,
            I => \N__40002\
        );

    \I__8797\ : InMux
    port map (
            O => \N__40014\,
            I => \N__40002\
        );

    \I__8796\ : InMux
    port map (
            O => \N__40011\,
            I => \N__39999\
        );

    \I__8795\ : InMux
    port map (
            O => \N__40010\,
            I => \N__39996\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__40007\,
            I => \N__39991\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__40002\,
            I => \N__39991\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__39999\,
            I => \N__39984\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__39996\,
            I => \N__39984\
        );

    \I__8790\ : Span4Mux_v
    port map (
            O => \N__39991\,
            I => \N__39984\
        );

    \I__8789\ : Odrv4
    port map (
            O => \N__39984\,
            I => measured_delay_tr_3
        );

    \I__8788\ : InMux
    port map (
            O => \N__39981\,
            I => \N__39978\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__39978\,
            I => \N__39973\
        );

    \I__8786\ : InMux
    port map (
            O => \N__39977\,
            I => \N__39969\
        );

    \I__8785\ : InMux
    port map (
            O => \N__39976\,
            I => \N__39966\
        );

    \I__8784\ : Span4Mux_v
    port map (
            O => \N__39973\,
            I => \N__39963\
        );

    \I__8783\ : InMux
    port map (
            O => \N__39972\,
            I => \N__39960\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__39969\,
            I => \N__39957\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__39966\,
            I => \N__39952\
        );

    \I__8780\ : Span4Mux_v
    port map (
            O => \N__39963\,
            I => \N__39952\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__39960\,
            I => \N__39947\
        );

    \I__8778\ : Span4Mux_h
    port map (
            O => \N__39957\,
            I => \N__39947\
        );

    \I__8777\ : Odrv4
    port map (
            O => \N__39952\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8776\ : Odrv4
    port map (
            O => \N__39947\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8775\ : InMux
    port map (
            O => \N__39942\,
            I => \N__39908\
        );

    \I__8774\ : InMux
    port map (
            O => \N__39941\,
            I => \N__39908\
        );

    \I__8773\ : InMux
    port map (
            O => \N__39940\,
            I => \N__39908\
        );

    \I__8772\ : InMux
    port map (
            O => \N__39939\,
            I => \N__39908\
        );

    \I__8771\ : InMux
    port map (
            O => \N__39938\,
            I => \N__39899\
        );

    \I__8770\ : InMux
    port map (
            O => \N__39937\,
            I => \N__39899\
        );

    \I__8769\ : InMux
    port map (
            O => \N__39936\,
            I => \N__39899\
        );

    \I__8768\ : InMux
    port map (
            O => \N__39935\,
            I => \N__39899\
        );

    \I__8767\ : InMux
    port map (
            O => \N__39934\,
            I => \N__39890\
        );

    \I__8766\ : InMux
    port map (
            O => \N__39933\,
            I => \N__39890\
        );

    \I__8765\ : InMux
    port map (
            O => \N__39932\,
            I => \N__39890\
        );

    \I__8764\ : InMux
    port map (
            O => \N__39931\,
            I => \N__39890\
        );

    \I__8763\ : InMux
    port map (
            O => \N__39930\,
            I => \N__39877\
        );

    \I__8762\ : InMux
    port map (
            O => \N__39929\,
            I => \N__39877\
        );

    \I__8761\ : InMux
    port map (
            O => \N__39928\,
            I => \N__39877\
        );

    \I__8760\ : InMux
    port map (
            O => \N__39927\,
            I => \N__39877\
        );

    \I__8759\ : InMux
    port map (
            O => \N__39926\,
            I => \N__39868\
        );

    \I__8758\ : InMux
    port map (
            O => \N__39925\,
            I => \N__39868\
        );

    \I__8757\ : InMux
    port map (
            O => \N__39924\,
            I => \N__39868\
        );

    \I__8756\ : InMux
    port map (
            O => \N__39923\,
            I => \N__39868\
        );

    \I__8755\ : InMux
    port map (
            O => \N__39922\,
            I => \N__39863\
        );

    \I__8754\ : InMux
    port map (
            O => \N__39921\,
            I => \N__39863\
        );

    \I__8753\ : InMux
    port map (
            O => \N__39920\,
            I => \N__39854\
        );

    \I__8752\ : InMux
    port map (
            O => \N__39919\,
            I => \N__39854\
        );

    \I__8751\ : InMux
    port map (
            O => \N__39918\,
            I => \N__39854\
        );

    \I__8750\ : InMux
    port map (
            O => \N__39917\,
            I => \N__39854\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__39908\,
            I => \N__39847\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__39899\,
            I => \N__39847\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__39890\,
            I => \N__39847\
        );

    \I__8746\ : InMux
    port map (
            O => \N__39889\,
            I => \N__39838\
        );

    \I__8745\ : InMux
    port map (
            O => \N__39888\,
            I => \N__39838\
        );

    \I__8744\ : InMux
    port map (
            O => \N__39887\,
            I => \N__39838\
        );

    \I__8743\ : InMux
    port map (
            O => \N__39886\,
            I => \N__39838\
        );

    \I__8742\ : LocalMux
    port map (
            O => \N__39877\,
            I => \N__39835\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__39868\,
            I => \N__39830\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__39863\,
            I => \N__39830\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__39854\,
            I => \N__39827\
        );

    \I__8738\ : Span4Mux_v
    port map (
            O => \N__39847\,
            I => \N__39824\
        );

    \I__8737\ : LocalMux
    port map (
            O => \N__39838\,
            I => \N__39815\
        );

    \I__8736\ : Span4Mux_h
    port map (
            O => \N__39835\,
            I => \N__39815\
        );

    \I__8735\ : Span4Mux_v
    port map (
            O => \N__39830\,
            I => \N__39815\
        );

    \I__8734\ : Span4Mux_v
    port map (
            O => \N__39827\,
            I => \N__39815\
        );

    \I__8733\ : Odrv4
    port map (
            O => \N__39824\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__8732\ : Odrv4
    port map (
            O => \N__39815\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__8731\ : CascadeMux
    port map (
            O => \N__39810\,
            I => \N__39807\
        );

    \I__8730\ : InMux
    port map (
            O => \N__39807\,
            I => \N__39804\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__39804\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\
        );

    \I__8728\ : CascadeMux
    port map (
            O => \N__39801\,
            I => \N__39798\
        );

    \I__8727\ : InMux
    port map (
            O => \N__39798\,
            I => \N__39794\
        );

    \I__8726\ : InMux
    port map (
            O => \N__39797\,
            I => \N__39790\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__39794\,
            I => \N__39787\
        );

    \I__8724\ : InMux
    port map (
            O => \N__39793\,
            I => \N__39784\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__39790\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8722\ : Odrv12
    port map (
            O => \N__39787\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__39784\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8720\ : InMux
    port map (
            O => \N__39777\,
            I => \N__39774\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__39774\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_1\
        );

    \I__8718\ : CascadeMux
    port map (
            O => \N__39771\,
            I => \N__39768\
        );

    \I__8717\ : InMux
    port map (
            O => \N__39768\,
            I => \N__39765\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__39765\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\
        );

    \I__8715\ : InMux
    port map (
            O => \N__39762\,
            I => \N__39758\
        );

    \I__8714\ : InMux
    port map (
            O => \N__39761\,
            I => \N__39755\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__39758\,
            I => \N__39752\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__39755\,
            I => \N__39749\
        );

    \I__8711\ : Odrv4
    port map (
            O => \N__39752\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8710\ : Odrv4
    port map (
            O => \N__39749\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8709\ : InMux
    port map (
            O => \N__39744\,
            I => \N__39741\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__39741\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_2\
        );

    \I__8707\ : CascadeMux
    port map (
            O => \N__39738\,
            I => \N__39735\
        );

    \I__8706\ : InMux
    port map (
            O => \N__39735\,
            I => \N__39731\
        );

    \I__8705\ : InMux
    port map (
            O => \N__39734\,
            I => \N__39728\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__39731\,
            I => \N__39725\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__39728\,
            I => \N__39722\
        );

    \I__8702\ : Odrv4
    port map (
            O => \N__39725\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8701\ : Odrv4
    port map (
            O => \N__39722\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8700\ : CascadeMux
    port map (
            O => \N__39717\,
            I => \N__39714\
        );

    \I__8699\ : InMux
    port map (
            O => \N__39714\,
            I => \N__39711\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__39711\,
            I => \N__39708\
        );

    \I__8697\ : Odrv4
    port map (
            O => \N__39708\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\
        );

    \I__8696\ : InMux
    port map (
            O => \N__39705\,
            I => \N__39702\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__39702\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_3\
        );

    \I__8694\ : InMux
    port map (
            O => \N__39699\,
            I => \N__39695\
        );

    \I__8693\ : InMux
    port map (
            O => \N__39698\,
            I => \N__39692\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__39695\,
            I => \N__39689\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__39692\,
            I => \N__39686\
        );

    \I__8690\ : Span4Mux_h
    port map (
            O => \N__39689\,
            I => \N__39683\
        );

    \I__8689\ : Span4Mux_h
    port map (
            O => \N__39686\,
            I => \N__39680\
        );

    \I__8688\ : Odrv4
    port map (
            O => \N__39683\,
            I => \delay_measurement_inst.N_284_1\
        );

    \I__8687\ : Odrv4
    port map (
            O => \N__39680\,
            I => \delay_measurement_inst.N_284_1\
        );

    \I__8686\ : InMux
    port map (
            O => \N__39675\,
            I => \N__39672\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__39672\,
            I => \N__39666\
        );

    \I__8684\ : InMux
    port map (
            O => \N__39671\,
            I => \N__39662\
        );

    \I__8683\ : InMux
    port map (
            O => \N__39670\,
            I => \N__39657\
        );

    \I__8682\ : InMux
    port map (
            O => \N__39669\,
            I => \N__39657\
        );

    \I__8681\ : Span4Mux_h
    port map (
            O => \N__39666\,
            I => \N__39654\
        );

    \I__8680\ : InMux
    port map (
            O => \N__39665\,
            I => \N__39650\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__39662\,
            I => \N__39647\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__39657\,
            I => \N__39644\
        );

    \I__8677\ : Span4Mux_v
    port map (
            O => \N__39654\,
            I => \N__39640\
        );

    \I__8676\ : InMux
    port map (
            O => \N__39653\,
            I => \N__39637\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__39650\,
            I => \N__39630\
        );

    \I__8674\ : Span4Mux_v
    port map (
            O => \N__39647\,
            I => \N__39630\
        );

    \I__8673\ : Span4Mux_h
    port map (
            O => \N__39644\,
            I => \N__39630\
        );

    \I__8672\ : InMux
    port map (
            O => \N__39643\,
            I => \N__39627\
        );

    \I__8671\ : Odrv4
    port map (
            O => \N__39640\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__39637\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__8669\ : Odrv4
    port map (
            O => \N__39630\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__39627\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__8667\ : InMux
    port map (
            O => \N__39618\,
            I => \N__39615\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__39615\,
            I => \N__39611\
        );

    \I__8665\ : InMux
    port map (
            O => \N__39614\,
            I => \N__39608\
        );

    \I__8664\ : Span4Mux_v
    port map (
            O => \N__39611\,
            I => \N__39603\
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__39608\,
            I => \N__39603\
        );

    \I__8662\ : Span4Mux_h
    port map (
            O => \N__39603\,
            I => \N__39599\
        );

    \I__8661\ : InMux
    port map (
            O => \N__39602\,
            I => \N__39596\
        );

    \I__8660\ : Odrv4
    port map (
            O => \N__39599\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__39596\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i\
        );

    \I__8658\ : InMux
    port map (
            O => \N__39591\,
            I => \N__39588\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__39588\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\
        );

    \I__8656\ : InMux
    port map (
            O => \N__39585\,
            I => \N__39582\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__39582\,
            I => \N__39579\
        );

    \I__8654\ : Span4Mux_v
    port map (
            O => \N__39579\,
            I => \N__39576\
        );

    \I__8653\ : Span4Mux_h
    port map (
            O => \N__39576\,
            I => \N__39571\
        );

    \I__8652\ : InMux
    port map (
            O => \N__39575\,
            I => \N__39568\
        );

    \I__8651\ : InMux
    port map (
            O => \N__39574\,
            I => \N__39565\
        );

    \I__8650\ : Odrv4
    port map (
            O => \N__39571\,
            I => measured_delay_tr_8
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__39568\,
            I => measured_delay_tr_8
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__39565\,
            I => measured_delay_tr_8
        );

    \I__8647\ : InMux
    port map (
            O => \N__39558\,
            I => \N__39555\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__39555\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\
        );

    \I__8645\ : InMux
    port map (
            O => \N__39552\,
            I => \N__39549\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__39549\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\
        );

    \I__8643\ : InMux
    port map (
            O => \N__39546\,
            I => \N__39543\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__39543\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\
        );

    \I__8641\ : InMux
    port map (
            O => \N__39540\,
            I => \N__39537\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__39537\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\
        );

    \I__8639\ : InMux
    port map (
            O => \N__39534\,
            I => \N__39531\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__39531\,
            I => \N__39525\
        );

    \I__8637\ : InMux
    port map (
            O => \N__39530\,
            I => \N__39520\
        );

    \I__8636\ : InMux
    port map (
            O => \N__39529\,
            I => \N__39520\
        );

    \I__8635\ : InMux
    port map (
            O => \N__39528\,
            I => \N__39517\
        );

    \I__8634\ : Span4Mux_h
    port map (
            O => \N__39525\,
            I => \N__39514\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__39520\,
            I => \N__39511\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__39517\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__8631\ : Odrv4
    port map (
            O => \N__39514\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__8630\ : Odrv12
    port map (
            O => \N__39511\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__8629\ : InMux
    port map (
            O => \N__39504\,
            I => \N__39501\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__39501\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\
        );

    \I__8627\ : InMux
    port map (
            O => \N__39498\,
            I => \N__39495\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__39495\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\
        );

    \I__8625\ : InMux
    port map (
            O => \N__39492\,
            I => \N__39489\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__39489\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\
        );

    \I__8623\ : InMux
    port map (
            O => \N__39486\,
            I => \N__39483\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__39483\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\
        );

    \I__8621\ : CascadeMux
    port map (
            O => \N__39480\,
            I => \N__39477\
        );

    \I__8620\ : InMux
    port map (
            O => \N__39477\,
            I => \N__39474\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__39474\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\
        );

    \I__8618\ : InMux
    port map (
            O => \N__39471\,
            I => \N__39468\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__39468\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_15\
        );

    \I__8616\ : CascadeMux
    port map (
            O => \N__39465\,
            I => \N__39462\
        );

    \I__8615\ : InMux
    port map (
            O => \N__39462\,
            I => \N__39459\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__39459\,
            I => \N__39456\
        );

    \I__8613\ : Odrv4
    port map (
            O => \N__39456\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\
        );

    \I__8612\ : InMux
    port map (
            O => \N__39453\,
            I => \N__39450\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__39450\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_16\
        );

    \I__8610\ : CascadeMux
    port map (
            O => \N__39447\,
            I => \N__39444\
        );

    \I__8609\ : InMux
    port map (
            O => \N__39444\,
            I => \N__39441\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__39441\,
            I => \N__39438\
        );

    \I__8607\ : Span4Mux_h
    port map (
            O => \N__39438\,
            I => \N__39435\
        );

    \I__8606\ : Odrv4
    port map (
            O => \N__39435\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\
        );

    \I__8605\ : InMux
    port map (
            O => \N__39432\,
            I => \N__39429\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__39429\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_17\
        );

    \I__8603\ : CascadeMux
    port map (
            O => \N__39426\,
            I => \N__39423\
        );

    \I__8602\ : InMux
    port map (
            O => \N__39423\,
            I => \N__39420\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__39420\,
            I => \N__39417\
        );

    \I__8600\ : Span4Mux_h
    port map (
            O => \N__39417\,
            I => \N__39414\
        );

    \I__8599\ : Odrv4
    port map (
            O => \N__39414\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\
        );

    \I__8598\ : InMux
    port map (
            O => \N__39411\,
            I => \N__39408\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__39408\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_18\
        );

    \I__8596\ : CascadeMux
    port map (
            O => \N__39405\,
            I => \N__39402\
        );

    \I__8595\ : InMux
    port map (
            O => \N__39402\,
            I => \N__39399\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__39399\,
            I => \N__39396\
        );

    \I__8593\ : Span4Mux_h
    port map (
            O => \N__39396\,
            I => \N__39393\
        );

    \I__8592\ : Odrv4
    port map (
            O => \N__39393\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\
        );

    \I__8591\ : InMux
    port map (
            O => \N__39390\,
            I => \N__39387\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__39387\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_19\
        );

    \I__8589\ : InMux
    port map (
            O => \N__39384\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__8588\ : CascadeMux
    port map (
            O => \N__39381\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\
        );

    \I__8587\ : InMux
    port map (
            O => \N__39378\,
            I => \N__39375\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__39375\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__8585\ : CascadeMux
    port map (
            O => \N__39372\,
            I => \N__39369\
        );

    \I__8584\ : InMux
    port map (
            O => \N__39369\,
            I => \N__39366\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__39366\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\
        );

    \I__8582\ : InMux
    port map (
            O => \N__39363\,
            I => \N__39360\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__39360\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_7\
        );

    \I__8580\ : CascadeMux
    port map (
            O => \N__39357\,
            I => \N__39354\
        );

    \I__8579\ : InMux
    port map (
            O => \N__39354\,
            I => \N__39351\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__39351\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\
        );

    \I__8577\ : InMux
    port map (
            O => \N__39348\,
            I => \N__39345\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__39345\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_8\
        );

    \I__8575\ : CascadeMux
    port map (
            O => \N__39342\,
            I => \N__39339\
        );

    \I__8574\ : InMux
    port map (
            O => \N__39339\,
            I => \N__39336\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__39336\,
            I => \N__39333\
        );

    \I__8572\ : Odrv12
    port map (
            O => \N__39333\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\
        );

    \I__8571\ : InMux
    port map (
            O => \N__39330\,
            I => \N__39327\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__39327\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_9\
        );

    \I__8569\ : CascadeMux
    port map (
            O => \N__39324\,
            I => \N__39321\
        );

    \I__8568\ : InMux
    port map (
            O => \N__39321\,
            I => \N__39318\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__39318\,
            I => \N__39315\
        );

    \I__8566\ : Odrv4
    port map (
            O => \N__39315\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\
        );

    \I__8565\ : InMux
    port map (
            O => \N__39312\,
            I => \N__39309\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__39309\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_10\
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__39306\,
            I => \N__39303\
        );

    \I__8562\ : InMux
    port map (
            O => \N__39303\,
            I => \N__39300\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__39300\,
            I => \N__39297\
        );

    \I__8560\ : Span4Mux_h
    port map (
            O => \N__39297\,
            I => \N__39294\
        );

    \I__8559\ : Span4Mux_h
    port map (
            O => \N__39294\,
            I => \N__39291\
        );

    \I__8558\ : Odrv4
    port map (
            O => \N__39291\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\
        );

    \I__8557\ : InMux
    port map (
            O => \N__39288\,
            I => \N__39285\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__39285\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_11\
        );

    \I__8555\ : CascadeMux
    port map (
            O => \N__39282\,
            I => \N__39279\
        );

    \I__8554\ : InMux
    port map (
            O => \N__39279\,
            I => \N__39276\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__39276\,
            I => \N__39273\
        );

    \I__8552\ : Span4Mux_h
    port map (
            O => \N__39273\,
            I => \N__39270\
        );

    \I__8551\ : Odrv4
    port map (
            O => \N__39270\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\
        );

    \I__8550\ : InMux
    port map (
            O => \N__39267\,
            I => \N__39264\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__39264\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_12\
        );

    \I__8548\ : InMux
    port map (
            O => \N__39261\,
            I => \N__39258\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__39258\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\
        );

    \I__8546\ : CascadeMux
    port map (
            O => \N__39255\,
            I => \N__39252\
        );

    \I__8545\ : InMux
    port map (
            O => \N__39252\,
            I => \N__39249\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__39249\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_13\
        );

    \I__8543\ : CascadeMux
    port map (
            O => \N__39246\,
            I => \N__39243\
        );

    \I__8542\ : InMux
    port map (
            O => \N__39243\,
            I => \N__39240\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__39240\,
            I => \N__39237\
        );

    \I__8540\ : Odrv4
    port map (
            O => \N__39237\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\
        );

    \I__8539\ : InMux
    port map (
            O => \N__39234\,
            I => \N__39231\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__39231\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_14\
        );

    \I__8537\ : InMux
    port map (
            O => \N__39228\,
            I => \N__39225\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__39225\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\
        );

    \I__8535\ : InMux
    port map (
            O => \N__39222\,
            I => \N__39219\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__39219\,
            I => \N__39216\
        );

    \I__8533\ : Odrv12
    port map (
            O => \N__39216\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_6\
        );

    \I__8532\ : CascadeMux
    port map (
            O => \N__39213\,
            I => \N__39210\
        );

    \I__8531\ : InMux
    port map (
            O => \N__39210\,
            I => \N__39207\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__39207\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_0\
        );

    \I__8529\ : CascadeMux
    port map (
            O => \N__39204\,
            I => \N__39201\
        );

    \I__8528\ : InMux
    port map (
            O => \N__39201\,
            I => \N__39198\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__39198\,
            I => \N__39195\
        );

    \I__8526\ : Odrv4
    port map (
            O => \N__39195\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\
        );

    \I__8525\ : InMux
    port map (
            O => \N__39192\,
            I => \N__39189\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__39189\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_1\
        );

    \I__8523\ : CascadeMux
    port map (
            O => \N__39186\,
            I => \N__39183\
        );

    \I__8522\ : InMux
    port map (
            O => \N__39183\,
            I => \N__39180\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__39180\,
            I => \N__39177\
        );

    \I__8520\ : Odrv4
    port map (
            O => \N__39177\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\
        );

    \I__8519\ : InMux
    port map (
            O => \N__39174\,
            I => \N__39171\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__39171\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_2\
        );

    \I__8517\ : CascadeMux
    port map (
            O => \N__39168\,
            I => \N__39165\
        );

    \I__8516\ : InMux
    port map (
            O => \N__39165\,
            I => \N__39162\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__39162\,
            I => \N__39159\
        );

    \I__8514\ : Odrv4
    port map (
            O => \N__39159\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\
        );

    \I__8513\ : InMux
    port map (
            O => \N__39156\,
            I => \N__39153\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__39153\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_3\
        );

    \I__8511\ : CascadeMux
    port map (
            O => \N__39150\,
            I => \N__39147\
        );

    \I__8510\ : InMux
    port map (
            O => \N__39147\,
            I => \N__39144\
        );

    \I__8509\ : LocalMux
    port map (
            O => \N__39144\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\
        );

    \I__8508\ : InMux
    port map (
            O => \N__39141\,
            I => \N__39138\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__39138\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_4\
        );

    \I__8506\ : CascadeMux
    port map (
            O => \N__39135\,
            I => \N__39132\
        );

    \I__8505\ : InMux
    port map (
            O => \N__39132\,
            I => \N__39129\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__39129\,
            I => \N__39126\
        );

    \I__8503\ : Odrv4
    port map (
            O => \N__39126\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\
        );

    \I__8502\ : InMux
    port map (
            O => \N__39123\,
            I => \N__39120\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__39120\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_5\
        );

    \I__8500\ : CascadeMux
    port map (
            O => \N__39117\,
            I => \N__39114\
        );

    \I__8499\ : InMux
    port map (
            O => \N__39114\,
            I => \N__39111\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__39111\,
            I => \N__39108\
        );

    \I__8497\ : Odrv4
    port map (
            O => \N__39108\,
            I => \phase_controller_slave.stoper_hc.target_timeZ1Z_6\
        );

    \I__8496\ : InMux
    port map (
            O => \N__39105\,
            I => \N__39102\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__39102\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_6\
        );

    \I__8494\ : CascadeMux
    port map (
            O => \N__39099\,
            I => \N__39096\
        );

    \I__8493\ : InMux
    port map (
            O => \N__39096\,
            I => \N__39093\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__39093\,
            I => \N__39090\
        );

    \I__8491\ : Odrv4
    port map (
            O => \N__39090\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1\
        );

    \I__8490\ : CascadeMux
    port map (
            O => \N__39087\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1_cascade_\
        );

    \I__8489\ : InMux
    port map (
            O => \N__39084\,
            I => \N__39081\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__39081\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0\
        );

    \I__8487\ : InMux
    port map (
            O => \N__39078\,
            I => \N__39074\
        );

    \I__8486\ : InMux
    port map (
            O => \N__39077\,
            I => \N__39071\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__39074\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__39071\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\
        );

    \I__8483\ : InMux
    port map (
            O => \N__39066\,
            I => \N__39063\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__39063\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_0\
        );

    \I__8481\ : InMux
    port map (
            O => \N__39060\,
            I => \N__39057\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__39057\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4\
        );

    \I__8479\ : CascadeMux
    port map (
            O => \N__39054\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_3_cascade_\
        );

    \I__8478\ : InMux
    port map (
            O => \N__39051\,
            I => \N__39048\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__39048\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30\
        );

    \I__8476\ : CascadeMux
    port map (
            O => \N__39045\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_cascade_\
        );

    \I__8475\ : InMux
    port map (
            O => \N__39042\,
            I => \N__39034\
        );

    \I__8474\ : InMux
    port map (
            O => \N__39041\,
            I => \N__39031\
        );

    \I__8473\ : InMux
    port map (
            O => \N__39040\,
            I => \N__39022\
        );

    \I__8472\ : InMux
    port map (
            O => \N__39039\,
            I => \N__39022\
        );

    \I__8471\ : InMux
    port map (
            O => \N__39038\,
            I => \N__39019\
        );

    \I__8470\ : InMux
    port map (
            O => \N__39037\,
            I => \N__39016\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__39034\,
            I => \N__39010\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__39031\,
            I => \N__39010\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39030\,
            I => \N__39007\
        );

    \I__8466\ : InMux
    port map (
            O => \N__39029\,
            I => \N__38998\
        );

    \I__8465\ : InMux
    port map (
            O => \N__39028\,
            I => \N__38998\
        );

    \I__8464\ : InMux
    port map (
            O => \N__39027\,
            I => \N__38998\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__39022\,
            I => \N__38995\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__39019\,
            I => \N__38990\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__39016\,
            I => \N__38990\
        );

    \I__8460\ : InMux
    port map (
            O => \N__39015\,
            I => \N__38987\
        );

    \I__8459\ : Span4Mux_h
    port map (
            O => \N__39010\,
            I => \N__38982\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__39007\,
            I => \N__38982\
        );

    \I__8457\ : InMux
    port map (
            O => \N__39006\,
            I => \N__38979\
        );

    \I__8456\ : InMux
    port map (
            O => \N__39005\,
            I => \N__38976\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__38998\,
            I => \N__38973\
        );

    \I__8454\ : Span4Mux_v
    port map (
            O => \N__38995\,
            I => \N__38966\
        );

    \I__8453\ : Span4Mux_v
    port map (
            O => \N__38990\,
            I => \N__38966\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__38987\,
            I => \N__38966\
        );

    \I__8451\ : Span4Mux_h
    port map (
            O => \N__38982\,
            I => \N__38961\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__38979\,
            I => \N__38961\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__38976\,
            I => \N__38958\
        );

    \I__8448\ : Span4Mux_v
    port map (
            O => \N__38973\,
            I => \N__38955\
        );

    \I__8447\ : Span4Mux_h
    port map (
            O => \N__38966\,
            I => \N__38948\
        );

    \I__8446\ : Span4Mux_v
    port map (
            O => \N__38961\,
            I => \N__38948\
        );

    \I__8445\ : Span4Mux_v
    port map (
            O => \N__38958\,
            I => \N__38948\
        );

    \I__8444\ : Odrv4
    port map (
            O => \N__38955\,
            I => \delay_measurement_inst.delay_hc_reg3lt31_0\
        );

    \I__8443\ : Odrv4
    port map (
            O => \N__38948\,
            I => \delay_measurement_inst.delay_hc_reg3lt31_0\
        );

    \I__8442\ : InMux
    port map (
            O => \N__38943\,
            I => \N__38940\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__38940\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_4\
        );

    \I__8440\ : CascadeMux
    port map (
            O => \N__38937\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_5_cascade_\
        );

    \I__8439\ : CascadeMux
    port map (
            O => \N__38934\,
            I => \N__38931\
        );

    \I__8438\ : InMux
    port map (
            O => \N__38931\,
            I => \N__38928\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__38928\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt13_0\
        );

    \I__8436\ : InMux
    port map (
            O => \N__38925\,
            I => \N__38922\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__38922\,
            I => \N__38919\
        );

    \I__8434\ : Odrv4
    port map (
            O => \N__38919\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt19\
        );

    \I__8433\ : CascadeMux
    port map (
            O => \N__38916\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_\
        );

    \I__8432\ : InMux
    port map (
            O => \N__38913\,
            I => \N__38910\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__38910\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\
        );

    \I__8430\ : InMux
    port map (
            O => \N__38907\,
            I => \N__38904\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__38904\,
            I => \N__38901\
        );

    \I__8428\ : Odrv4
    port map (
            O => \N__38901\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclt31_0\
        );

    \I__8427\ : InMux
    port map (
            O => \N__38898\,
            I => \N__38895\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__38895\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_7\
        );

    \I__8425\ : InMux
    port map (
            O => \N__38892\,
            I => \N__38889\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__38889\,
            I => \N__38886\
        );

    \I__8423\ : Odrv4
    port map (
            O => \N__38886\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3\
        );

    \I__8422\ : InMux
    port map (
            O => \N__38883\,
            I => \N__38880\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__38880\,
            I => \N__38877\
        );

    \I__8420\ : Odrv4
    port map (
            O => \N__38877\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1\
        );

    \I__8419\ : CascadeMux
    port map (
            O => \N__38874\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz_cascade_\
        );

    \I__8418\ : CascadeMux
    port map (
            O => \N__38871\,
            I => \N__38866\
        );

    \I__8417\ : InMux
    port map (
            O => \N__38870\,
            I => \N__38863\
        );

    \I__8416\ : InMux
    port map (
            O => \N__38869\,
            I => \N__38860\
        );

    \I__8415\ : InMux
    port map (
            O => \N__38866\,
            I => \N__38857\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__38863\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__38860\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__38857\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__8411\ : InMux
    port map (
            O => \N__38850\,
            I => \bfn_15_22_0_\
        );

    \I__8410\ : CascadeMux
    port map (
            O => \N__38847\,
            I => \N__38842\
        );

    \I__8409\ : InMux
    port map (
            O => \N__38846\,
            I => \N__38839\
        );

    \I__8408\ : InMux
    port map (
            O => \N__38845\,
            I => \N__38836\
        );

    \I__8407\ : InMux
    port map (
            O => \N__38842\,
            I => \N__38833\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__38839\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__38836\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__38833\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__8403\ : InMux
    port map (
            O => \N__38826\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__8402\ : CascadeMux
    port map (
            O => \N__38823\,
            I => \N__38818\
        );

    \I__8401\ : InMux
    port map (
            O => \N__38822\,
            I => \N__38815\
        );

    \I__8400\ : InMux
    port map (
            O => \N__38821\,
            I => \N__38812\
        );

    \I__8399\ : InMux
    port map (
            O => \N__38818\,
            I => \N__38809\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__38815\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__38812\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__38809\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__8395\ : InMux
    port map (
            O => \N__38802\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__8394\ : CascadeMux
    port map (
            O => \N__38799\,
            I => \N__38794\
        );

    \I__8393\ : InMux
    port map (
            O => \N__38798\,
            I => \N__38791\
        );

    \I__8392\ : InMux
    port map (
            O => \N__38797\,
            I => \N__38788\
        );

    \I__8391\ : InMux
    port map (
            O => \N__38794\,
            I => \N__38785\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__38791\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__38788\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__38785\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__8387\ : InMux
    port map (
            O => \N__38778\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__8386\ : CascadeMux
    port map (
            O => \N__38775\,
            I => \N__38771\
        );

    \I__8385\ : InMux
    port map (
            O => \N__38774\,
            I => \N__38768\
        );

    \I__8384\ : InMux
    port map (
            O => \N__38771\,
            I => \N__38765\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__38768\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__38765\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__8381\ : InMux
    port map (
            O => \N__38760\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__8380\ : InMux
    port map (
            O => \N__38757\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__8379\ : CascadeMux
    port map (
            O => \N__38754\,
            I => \N__38750\
        );

    \I__8378\ : InMux
    port map (
            O => \N__38753\,
            I => \N__38747\
        );

    \I__8377\ : InMux
    port map (
            O => \N__38750\,
            I => \N__38744\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__38747\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__38744\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__8374\ : CEMux
    port map (
            O => \N__38739\,
            I => \N__38736\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__38736\,
            I => \N__38733\
        );

    \I__8372\ : Span4Mux_v
    port map (
            O => \N__38733\,
            I => \N__38728\
        );

    \I__8371\ : CEMux
    port map (
            O => \N__38732\,
            I => \N__38725\
        );

    \I__8370\ : CEMux
    port map (
            O => \N__38731\,
            I => \N__38721\
        );

    \I__8369\ : Span4Mux_h
    port map (
            O => \N__38728\,
            I => \N__38716\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__38725\,
            I => \N__38716\
        );

    \I__8367\ : CEMux
    port map (
            O => \N__38724\,
            I => \N__38713\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__38721\,
            I => \N__38710\
        );

    \I__8365\ : Span4Mux_v
    port map (
            O => \N__38716\,
            I => \N__38707\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__38713\,
            I => \N__38702\
        );

    \I__8363\ : Span4Mux_v
    port map (
            O => \N__38710\,
            I => \N__38702\
        );

    \I__8362\ : Odrv4
    port map (
            O => \N__38707\,
            I => \delay_measurement_inst.delay_tr_timer.N_338_i\
        );

    \I__8361\ : Odrv4
    port map (
            O => \N__38702\,
            I => \delay_measurement_inst.delay_tr_timer.N_338_i\
        );

    \I__8360\ : CascadeMux
    port map (
            O => \N__38697\,
            I => \N__38692\
        );

    \I__8359\ : InMux
    port map (
            O => \N__38696\,
            I => \N__38689\
        );

    \I__8358\ : InMux
    port map (
            O => \N__38695\,
            I => \N__38686\
        );

    \I__8357\ : InMux
    port map (
            O => \N__38692\,
            I => \N__38683\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__38689\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__38686\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__38683\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__8353\ : InMux
    port map (
            O => \N__38676\,
            I => \bfn_15_21_0_\
        );

    \I__8352\ : CascadeMux
    port map (
            O => \N__38673\,
            I => \N__38668\
        );

    \I__8351\ : InMux
    port map (
            O => \N__38672\,
            I => \N__38665\
        );

    \I__8350\ : InMux
    port map (
            O => \N__38671\,
            I => \N__38662\
        );

    \I__8349\ : InMux
    port map (
            O => \N__38668\,
            I => \N__38659\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__38665\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__38662\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__38659\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__8345\ : InMux
    port map (
            O => \N__38652\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__8344\ : CascadeMux
    port map (
            O => \N__38649\,
            I => \N__38644\
        );

    \I__8343\ : InMux
    port map (
            O => \N__38648\,
            I => \N__38641\
        );

    \I__8342\ : InMux
    port map (
            O => \N__38647\,
            I => \N__38638\
        );

    \I__8341\ : InMux
    port map (
            O => \N__38644\,
            I => \N__38635\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__38641\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__38638\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__38635\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__8337\ : InMux
    port map (
            O => \N__38628\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__8336\ : CascadeMux
    port map (
            O => \N__38625\,
            I => \N__38620\
        );

    \I__8335\ : InMux
    port map (
            O => \N__38624\,
            I => \N__38617\
        );

    \I__8334\ : InMux
    port map (
            O => \N__38623\,
            I => \N__38614\
        );

    \I__8333\ : InMux
    port map (
            O => \N__38620\,
            I => \N__38611\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__38617\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__38614\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__38611\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__8329\ : InMux
    port map (
            O => \N__38604\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__8328\ : CascadeMux
    port map (
            O => \N__38601\,
            I => \N__38596\
        );

    \I__8327\ : InMux
    port map (
            O => \N__38600\,
            I => \N__38593\
        );

    \I__8326\ : InMux
    port map (
            O => \N__38599\,
            I => \N__38590\
        );

    \I__8325\ : InMux
    port map (
            O => \N__38596\,
            I => \N__38587\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__38593\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__38590\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__38587\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__8321\ : InMux
    port map (
            O => \N__38580\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__8320\ : CascadeMux
    port map (
            O => \N__38577\,
            I => \N__38572\
        );

    \I__8319\ : InMux
    port map (
            O => \N__38576\,
            I => \N__38569\
        );

    \I__8318\ : InMux
    port map (
            O => \N__38575\,
            I => \N__38566\
        );

    \I__8317\ : InMux
    port map (
            O => \N__38572\,
            I => \N__38563\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__38569\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__38566\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__38563\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__8313\ : InMux
    port map (
            O => \N__38556\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__8312\ : CascadeMux
    port map (
            O => \N__38553\,
            I => \N__38548\
        );

    \I__8311\ : InMux
    port map (
            O => \N__38552\,
            I => \N__38545\
        );

    \I__8310\ : InMux
    port map (
            O => \N__38551\,
            I => \N__38542\
        );

    \I__8309\ : InMux
    port map (
            O => \N__38548\,
            I => \N__38539\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__38545\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__38542\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__38539\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__8305\ : InMux
    port map (
            O => \N__38532\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__8304\ : CascadeMux
    port map (
            O => \N__38529\,
            I => \N__38524\
        );

    \I__8303\ : InMux
    port map (
            O => \N__38528\,
            I => \N__38521\
        );

    \I__8302\ : InMux
    port map (
            O => \N__38527\,
            I => \N__38518\
        );

    \I__8301\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38515\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__38521\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__38518\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__38515\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__8297\ : InMux
    port map (
            O => \N__38508\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__8296\ : CascadeMux
    port map (
            O => \N__38505\,
            I => \N__38500\
        );

    \I__8295\ : InMux
    port map (
            O => \N__38504\,
            I => \N__38497\
        );

    \I__8294\ : InMux
    port map (
            O => \N__38503\,
            I => \N__38494\
        );

    \I__8293\ : InMux
    port map (
            O => \N__38500\,
            I => \N__38491\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__38497\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__38494\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__38491\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__8289\ : InMux
    port map (
            O => \N__38484\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__8288\ : CascadeMux
    port map (
            O => \N__38481\,
            I => \N__38476\
        );

    \I__8287\ : InMux
    port map (
            O => \N__38480\,
            I => \N__38473\
        );

    \I__8286\ : InMux
    port map (
            O => \N__38479\,
            I => \N__38470\
        );

    \I__8285\ : InMux
    port map (
            O => \N__38476\,
            I => \N__38467\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__38473\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__38470\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__38467\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__8281\ : InMux
    port map (
            O => \N__38460\,
            I => \bfn_15_20_0_\
        );

    \I__8280\ : CascadeMux
    port map (
            O => \N__38457\,
            I => \N__38452\
        );

    \I__8279\ : InMux
    port map (
            O => \N__38456\,
            I => \N__38449\
        );

    \I__8278\ : InMux
    port map (
            O => \N__38455\,
            I => \N__38446\
        );

    \I__8277\ : InMux
    port map (
            O => \N__38452\,
            I => \N__38443\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__38449\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__8275\ : LocalMux
    port map (
            O => \N__38446\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__38443\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__8273\ : InMux
    port map (
            O => \N__38436\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__8272\ : CascadeMux
    port map (
            O => \N__38433\,
            I => \N__38428\
        );

    \I__8271\ : InMux
    port map (
            O => \N__38432\,
            I => \N__38425\
        );

    \I__8270\ : InMux
    port map (
            O => \N__38431\,
            I => \N__38422\
        );

    \I__8269\ : InMux
    port map (
            O => \N__38428\,
            I => \N__38419\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__38425\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__38422\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__38419\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__8265\ : InMux
    port map (
            O => \N__38412\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__8264\ : CascadeMux
    port map (
            O => \N__38409\,
            I => \N__38404\
        );

    \I__8263\ : InMux
    port map (
            O => \N__38408\,
            I => \N__38401\
        );

    \I__8262\ : InMux
    port map (
            O => \N__38407\,
            I => \N__38398\
        );

    \I__8261\ : InMux
    port map (
            O => \N__38404\,
            I => \N__38395\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__38401\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__38398\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__38395\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__8257\ : InMux
    port map (
            O => \N__38388\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__8256\ : CascadeMux
    port map (
            O => \N__38385\,
            I => \N__38380\
        );

    \I__8255\ : InMux
    port map (
            O => \N__38384\,
            I => \N__38377\
        );

    \I__8254\ : InMux
    port map (
            O => \N__38383\,
            I => \N__38374\
        );

    \I__8253\ : InMux
    port map (
            O => \N__38380\,
            I => \N__38371\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__38377\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__38374\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__38371\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__8249\ : InMux
    port map (
            O => \N__38364\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__8248\ : CascadeMux
    port map (
            O => \N__38361\,
            I => \N__38356\
        );

    \I__8247\ : InMux
    port map (
            O => \N__38360\,
            I => \N__38353\
        );

    \I__8246\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38350\
        );

    \I__8245\ : InMux
    port map (
            O => \N__38356\,
            I => \N__38347\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__38353\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__38350\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__38347\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__8241\ : InMux
    port map (
            O => \N__38340\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__8240\ : CascadeMux
    port map (
            O => \N__38337\,
            I => \N__38332\
        );

    \I__8239\ : InMux
    port map (
            O => \N__38336\,
            I => \N__38329\
        );

    \I__8238\ : InMux
    port map (
            O => \N__38335\,
            I => \N__38326\
        );

    \I__8237\ : InMux
    port map (
            O => \N__38332\,
            I => \N__38323\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__38329\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__38326\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__38323\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__8233\ : InMux
    port map (
            O => \N__38316\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__8232\ : CascadeMux
    port map (
            O => \N__38313\,
            I => \N__38308\
        );

    \I__8231\ : InMux
    port map (
            O => \N__38312\,
            I => \N__38305\
        );

    \I__8230\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38302\
        );

    \I__8229\ : InMux
    port map (
            O => \N__38308\,
            I => \N__38299\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__38305\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__38302\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__38299\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__8225\ : InMux
    port map (
            O => \N__38292\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__8224\ : InMux
    port map (
            O => \N__38289\,
            I => \N__38286\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__38286\,
            I => \N__38283\
        );

    \I__8222\ : Span4Mux_v
    port map (
            O => \N__38283\,
            I => \N__38278\
        );

    \I__8221\ : InMux
    port map (
            O => \N__38282\,
            I => \N__38275\
        );

    \I__8220\ : InMux
    port map (
            O => \N__38281\,
            I => \N__38272\
        );

    \I__8219\ : Odrv4
    port map (
            O => \N__38278\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__38275\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__38272\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__8216\ : InMux
    port map (
            O => \N__38265\,
            I => \bfn_15_19_0_\
        );

    \I__8215\ : InMux
    port map (
            O => \N__38262\,
            I => \N__38259\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__38259\,
            I => \N__38256\
        );

    \I__8213\ : Span4Mux_v
    port map (
            O => \N__38256\,
            I => \N__38251\
        );

    \I__8212\ : InMux
    port map (
            O => \N__38255\,
            I => \N__38248\
        );

    \I__8211\ : InMux
    port map (
            O => \N__38254\,
            I => \N__38245\
        );

    \I__8210\ : Odrv4
    port map (
            O => \N__38251\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__38248\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__38245\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__8207\ : InMux
    port map (
            O => \N__38238\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__8206\ : CascadeMux
    port map (
            O => \N__38235\,
            I => \N__38230\
        );

    \I__8205\ : InMux
    port map (
            O => \N__38234\,
            I => \N__38227\
        );

    \I__8204\ : InMux
    port map (
            O => \N__38233\,
            I => \N__38224\
        );

    \I__8203\ : InMux
    port map (
            O => \N__38230\,
            I => \N__38221\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__38227\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__38224\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__38221\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__8199\ : InMux
    port map (
            O => \N__38214\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__8198\ : CascadeMux
    port map (
            O => \N__38211\,
            I => \N__38206\
        );

    \I__8197\ : InMux
    port map (
            O => \N__38210\,
            I => \N__38203\
        );

    \I__8196\ : InMux
    port map (
            O => \N__38209\,
            I => \N__38200\
        );

    \I__8195\ : InMux
    port map (
            O => \N__38206\,
            I => \N__38197\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__38203\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__38200\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__38197\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__8191\ : InMux
    port map (
            O => \N__38190\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__38187\,
            I => \N__38182\
        );

    \I__8189\ : InMux
    port map (
            O => \N__38186\,
            I => \N__38179\
        );

    \I__8188\ : InMux
    port map (
            O => \N__38185\,
            I => \N__38176\
        );

    \I__8187\ : InMux
    port map (
            O => \N__38182\,
            I => \N__38173\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__38179\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__38176\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__38173\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__8183\ : InMux
    port map (
            O => \N__38166\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__8182\ : CascadeMux
    port map (
            O => \N__38163\,
            I => \N__38158\
        );

    \I__8181\ : InMux
    port map (
            O => \N__38162\,
            I => \N__38155\
        );

    \I__8180\ : InMux
    port map (
            O => \N__38161\,
            I => \N__38152\
        );

    \I__8179\ : InMux
    port map (
            O => \N__38158\,
            I => \N__38149\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__38155\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__38152\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__38149\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__8175\ : InMux
    port map (
            O => \N__38142\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__8174\ : CascadeMux
    port map (
            O => \N__38139\,
            I => \N__38134\
        );

    \I__8173\ : InMux
    port map (
            O => \N__38138\,
            I => \N__38131\
        );

    \I__8172\ : InMux
    port map (
            O => \N__38137\,
            I => \N__38128\
        );

    \I__8171\ : InMux
    port map (
            O => \N__38134\,
            I => \N__38125\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__38131\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__38128\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__38125\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__8167\ : InMux
    port map (
            O => \N__38118\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__8166\ : CascadeMux
    port map (
            O => \N__38115\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__8165\ : InMux
    port map (
            O => \N__38112\,
            I => \N__38109\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__38109\,
            I => \N__38106\
        );

    \I__8163\ : Odrv4
    port map (
            O => \N__38106\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\
        );

    \I__8162\ : InMux
    port map (
            O => \N__38103\,
            I => \N__38100\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__38100\,
            I => \N__38097\
        );

    \I__8160\ : Odrv4
    port map (
            O => \N__38097\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\
        );

    \I__8159\ : InMux
    port map (
            O => \N__38094\,
            I => \N__38091\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__38091\,
            I => \N__38088\
        );

    \I__8157\ : Odrv4
    port map (
            O => \N__38088\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\
        );

    \I__8156\ : InMux
    port map (
            O => \N__38085\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__8155\ : InMux
    port map (
            O => \N__38082\,
            I => \N__38079\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__38079\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\
        );

    \I__8153\ : InMux
    port map (
            O => \N__38076\,
            I => \N__38072\
        );

    \I__8152\ : CascadeMux
    port map (
            O => \N__38075\,
            I => \N__38069\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__38072\,
            I => \N__38066\
        );

    \I__8150\ : InMux
    port map (
            O => \N__38069\,
            I => \N__38063\
        );

    \I__8149\ : Span4Mux_v
    port map (
            O => \N__38066\,
            I => \N__38057\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__38063\,
            I => \N__38057\
        );

    \I__8147\ : InMux
    port map (
            O => \N__38062\,
            I => \N__38053\
        );

    \I__8146\ : Span4Mux_h
    port map (
            O => \N__38057\,
            I => \N__38050\
        );

    \I__8145\ : InMux
    port map (
            O => \N__38056\,
            I => \N__38047\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__38053\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__8143\ : Odrv4
    port map (
            O => \N__38050\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__38047\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__8141\ : InMux
    port map (
            O => \N__38040\,
            I => \N__38037\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__38037\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\
        );

    \I__8139\ : InMux
    port map (
            O => \N__38034\,
            I => \N__38031\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__38031\,
            I => \N__38028\
        );

    \I__8137\ : Odrv12
    port map (
            O => \N__38028\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\
        );

    \I__8136\ : InMux
    port map (
            O => \N__38025\,
            I => \N__38022\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__38022\,
            I => \N__38019\
        );

    \I__8134\ : Odrv4
    port map (
            O => \N__38019\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\
        );

    \I__8133\ : InMux
    port map (
            O => \N__38016\,
            I => \N__38013\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__38013\,
            I => \N__38010\
        );

    \I__8131\ : Odrv4
    port map (
            O => \N__38010\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\
        );

    \I__8130\ : InMux
    port map (
            O => \N__38007\,
            I => \N__38004\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__38004\,
            I => \N__38001\
        );

    \I__8128\ : Odrv4
    port map (
            O => \N__38001\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\
        );

    \I__8127\ : InMux
    port map (
            O => \N__37998\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__8126\ : InMux
    port map (
            O => \N__37995\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__8125\ : InMux
    port map (
            O => \N__37992\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__8124\ : InMux
    port map (
            O => \N__37989\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__8123\ : InMux
    port map (
            O => \N__37986\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__8122\ : InMux
    port map (
            O => \N__37983\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__8121\ : InMux
    port map (
            O => \N__37980\,
            I => \N__37977\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__37977\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\
        );

    \I__8119\ : InMux
    port map (
            O => \N__37974\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__8118\ : InMux
    port map (
            O => \N__37971\,
            I => \bfn_15_15_0_\
        );

    \I__8117\ : InMux
    port map (
            O => \N__37968\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__8116\ : InMux
    port map (
            O => \N__37965\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__8115\ : InMux
    port map (
            O => \N__37962\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__8114\ : InMux
    port map (
            O => \N__37959\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__8113\ : InMux
    port map (
            O => \N__37956\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__8112\ : InMux
    port map (
            O => \N__37953\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__8111\ : InMux
    port map (
            O => \N__37950\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__8110\ : InMux
    port map (
            O => \N__37947\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__8109\ : InMux
    port map (
            O => \N__37944\,
            I => \bfn_15_14_0_\
        );

    \I__8108\ : InMux
    port map (
            O => \N__37941\,
            I => \N__37937\
        );

    \I__8107\ : CascadeMux
    port map (
            O => \N__37940\,
            I => \N__37933\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__37937\,
            I => \N__37929\
        );

    \I__8105\ : InMux
    port map (
            O => \N__37936\,
            I => \N__37925\
        );

    \I__8104\ : InMux
    port map (
            O => \N__37933\,
            I => \N__37922\
        );

    \I__8103\ : CascadeMux
    port map (
            O => \N__37932\,
            I => \N__37919\
        );

    \I__8102\ : Span4Mux_h
    port map (
            O => \N__37929\,
            I => \N__37916\
        );

    \I__8101\ : InMux
    port map (
            O => \N__37928\,
            I => \N__37913\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__37925\,
            I => \N__37910\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__37922\,
            I => \N__37907\
        );

    \I__8098\ : InMux
    port map (
            O => \N__37919\,
            I => \N__37904\
        );

    \I__8097\ : Span4Mux_v
    port map (
            O => \N__37916\,
            I => \N__37899\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__37913\,
            I => \N__37899\
        );

    \I__8095\ : Span4Mux_h
    port map (
            O => \N__37910\,
            I => \N__37894\
        );

    \I__8094\ : Span4Mux_h
    port map (
            O => \N__37907\,
            I => \N__37894\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__37904\,
            I => measured_delay_hc_8
        );

    \I__8092\ : Odrv4
    port map (
            O => \N__37899\,
            I => measured_delay_hc_8
        );

    \I__8091\ : Odrv4
    port map (
            O => \N__37894\,
            I => measured_delay_hc_8
        );

    \I__8090\ : InMux
    port map (
            O => \N__37887\,
            I => \N__37876\
        );

    \I__8089\ : InMux
    port map (
            O => \N__37886\,
            I => \N__37876\
        );

    \I__8088\ : InMux
    port map (
            O => \N__37885\,
            I => \N__37871\
        );

    \I__8087\ : InMux
    port map (
            O => \N__37884\,
            I => \N__37871\
        );

    \I__8086\ : CascadeMux
    port map (
            O => \N__37883\,
            I => \N__37866\
        );

    \I__8085\ : InMux
    port map (
            O => \N__37882\,
            I => \N__37862\
        );

    \I__8084\ : InMux
    port map (
            O => \N__37881\,
            I => \N__37859\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__37876\,
            I => \N__37856\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__37871\,
            I => \N__37853\
        );

    \I__8081\ : CascadeMux
    port map (
            O => \N__37870\,
            I => \N__37849\
        );

    \I__8080\ : CascadeMux
    port map (
            O => \N__37869\,
            I => \N__37845\
        );

    \I__8079\ : InMux
    port map (
            O => \N__37866\,
            I => \N__37836\
        );

    \I__8078\ : InMux
    port map (
            O => \N__37865\,
            I => \N__37836\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__37862\,
            I => \N__37833\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__37859\,
            I => \N__37830\
        );

    \I__8075\ : Span4Mux_h
    port map (
            O => \N__37856\,
            I => \N__37827\
        );

    \I__8074\ : Span4Mux_h
    port map (
            O => \N__37853\,
            I => \N__37824\
        );

    \I__8073\ : InMux
    port map (
            O => \N__37852\,
            I => \N__37821\
        );

    \I__8072\ : InMux
    port map (
            O => \N__37849\,
            I => \N__37818\
        );

    \I__8071\ : InMux
    port map (
            O => \N__37848\,
            I => \N__37815\
        );

    \I__8070\ : InMux
    port map (
            O => \N__37845\,
            I => \N__37810\
        );

    \I__8069\ : InMux
    port map (
            O => \N__37844\,
            I => \N__37810\
        );

    \I__8068\ : InMux
    port map (
            O => \N__37843\,
            I => \N__37805\
        );

    \I__8067\ : InMux
    port map (
            O => \N__37842\,
            I => \N__37805\
        );

    \I__8066\ : CascadeMux
    port map (
            O => \N__37841\,
            I => \N__37802\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__37836\,
            I => \N__37795\
        );

    \I__8064\ : Span4Mux_h
    port map (
            O => \N__37833\,
            I => \N__37795\
        );

    \I__8063\ : Span4Mux_v
    port map (
            O => \N__37830\,
            I => \N__37795\
        );

    \I__8062\ : Span4Mux_h
    port map (
            O => \N__37827\,
            I => \N__37790\
        );

    \I__8061\ : Span4Mux_v
    port map (
            O => \N__37824\,
            I => \N__37790\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__37821\,
            I => \N__37785\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__37818\,
            I => \N__37785\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__37815\,
            I => \N__37782\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__37810\,
            I => \N__37777\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__37805\,
            I => \N__37777\
        );

    \I__8055\ : InMux
    port map (
            O => \N__37802\,
            I => \N__37774\
        );

    \I__8054\ : Span4Mux_v
    port map (
            O => \N__37795\,
            I => \N__37771\
        );

    \I__8053\ : Span4Mux_v
    port map (
            O => \N__37790\,
            I => \N__37766\
        );

    \I__8052\ : Span4Mux_h
    port map (
            O => \N__37785\,
            I => \N__37766\
        );

    \I__8051\ : Span4Mux_h
    port map (
            O => \N__37782\,
            I => \N__37761\
        );

    \I__8050\ : Span4Mux_h
    port map (
            O => \N__37777\,
            I => \N__37761\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__37774\,
            I => measured_delay_hc_31
        );

    \I__8048\ : Odrv4
    port map (
            O => \N__37771\,
            I => measured_delay_hc_31
        );

    \I__8047\ : Odrv4
    port map (
            O => \N__37766\,
            I => measured_delay_hc_31
        );

    \I__8046\ : Odrv4
    port map (
            O => \N__37761\,
            I => measured_delay_hc_31
        );

    \I__8045\ : InMux
    port map (
            O => \N__37752\,
            I => \N__37748\
        );

    \I__8044\ : InMux
    port map (
            O => \N__37751\,
            I => \N__37744\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__37748\,
            I => \N__37740\
        );

    \I__8042\ : CascadeMux
    port map (
            O => \N__37747\,
            I => \N__37736\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__37744\,
            I => \N__37733\
        );

    \I__8040\ : InMux
    port map (
            O => \N__37743\,
            I => \N__37730\
        );

    \I__8039\ : Span4Mux_v
    port map (
            O => \N__37740\,
            I => \N__37727\
        );

    \I__8038\ : CascadeMux
    port map (
            O => \N__37739\,
            I => \N__37724\
        );

    \I__8037\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37721\
        );

    \I__8036\ : Span4Mux_h
    port map (
            O => \N__37733\,
            I => \N__37718\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__37730\,
            I => \N__37715\
        );

    \I__8034\ : Span4Mux_h
    port map (
            O => \N__37727\,
            I => \N__37712\
        );

    \I__8033\ : InMux
    port map (
            O => \N__37724\,
            I => \N__37709\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__37721\,
            I => measured_delay_hc_5
        );

    \I__8031\ : Odrv4
    port map (
            O => \N__37718\,
            I => measured_delay_hc_5
        );

    \I__8030\ : Odrv12
    port map (
            O => \N__37715\,
            I => measured_delay_hc_5
        );

    \I__8029\ : Odrv4
    port map (
            O => \N__37712\,
            I => measured_delay_hc_5
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__37709\,
            I => measured_delay_hc_5
        );

    \I__8027\ : InMux
    port map (
            O => \N__37698\,
            I => \N__37692\
        );

    \I__8026\ : InMux
    port map (
            O => \N__37697\,
            I => \N__37684\
        );

    \I__8025\ : InMux
    port map (
            O => \N__37696\,
            I => \N__37684\
        );

    \I__8024\ : InMux
    port map (
            O => \N__37695\,
            I => \N__37677\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__37692\,
            I => \N__37674\
        );

    \I__8022\ : InMux
    port map (
            O => \N__37691\,
            I => \N__37669\
        );

    \I__8021\ : InMux
    port map (
            O => \N__37690\,
            I => \N__37669\
        );

    \I__8020\ : InMux
    port map (
            O => \N__37689\,
            I => \N__37663\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__37684\,
            I => \N__37660\
        );

    \I__8018\ : InMux
    port map (
            O => \N__37683\,
            I => \N__37653\
        );

    \I__8017\ : InMux
    port map (
            O => \N__37682\,
            I => \N__37653\
        );

    \I__8016\ : InMux
    port map (
            O => \N__37681\,
            I => \N__37653\
        );

    \I__8015\ : InMux
    port map (
            O => \N__37680\,
            I => \N__37642\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__37677\,
            I => \N__37637\
        );

    \I__8013\ : Span4Mux_h
    port map (
            O => \N__37674\,
            I => \N__37637\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__37669\,
            I => \N__37634\
        );

    \I__8011\ : InMux
    port map (
            O => \N__37668\,
            I => \N__37627\
        );

    \I__8010\ : InMux
    port map (
            O => \N__37667\,
            I => \N__37627\
        );

    \I__8009\ : InMux
    port map (
            O => \N__37666\,
            I => \N__37627\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__37663\,
            I => \N__37624\
        );

    \I__8007\ : Span4Mux_v
    port map (
            O => \N__37660\,
            I => \N__37619\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__37653\,
            I => \N__37619\
        );

    \I__8005\ : InMux
    port map (
            O => \N__37652\,
            I => \N__37614\
        );

    \I__8004\ : InMux
    port map (
            O => \N__37651\,
            I => \N__37614\
        );

    \I__8003\ : InMux
    port map (
            O => \N__37650\,
            I => \N__37601\
        );

    \I__8002\ : InMux
    port map (
            O => \N__37649\,
            I => \N__37601\
        );

    \I__8001\ : InMux
    port map (
            O => \N__37648\,
            I => \N__37601\
        );

    \I__8000\ : InMux
    port map (
            O => \N__37647\,
            I => \N__37601\
        );

    \I__7999\ : InMux
    port map (
            O => \N__37646\,
            I => \N__37601\
        );

    \I__7998\ : InMux
    port map (
            O => \N__37645\,
            I => \N__37601\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__37642\,
            I => \N__37598\
        );

    \I__7996\ : Span4Mux_v
    port map (
            O => \N__37637\,
            I => \N__37595\
        );

    \I__7995\ : Span4Mux_h
    port map (
            O => \N__37634\,
            I => \N__37592\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__37627\,
            I => \N__37589\
        );

    \I__7993\ : Span4Mux_v
    port map (
            O => \N__37624\,
            I => \N__37582\
        );

    \I__7992\ : Span4Mux_h
    port map (
            O => \N__37619\,
            I => \N__37582\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__37614\,
            I => \N__37582\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__37601\,
            I => \N__37579\
        );

    \I__7989\ : Odrv12
    port map (
            O => \N__37598\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7988\ : Odrv4
    port map (
            O => \N__37595\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7987\ : Odrv4
    port map (
            O => \N__37592\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7986\ : Odrv12
    port map (
            O => \N__37589\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7985\ : Odrv4
    port map (
            O => \N__37582\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7984\ : Odrv12
    port map (
            O => \N__37579\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7983\ : CascadeMux
    port map (
            O => \N__37566\,
            I => \N__37563\
        );

    \I__7982\ : InMux
    port map (
            O => \N__37563\,
            I => \N__37557\
        );

    \I__7981\ : CascadeMux
    port map (
            O => \N__37562\,
            I => \N__37554\
        );

    \I__7980\ : InMux
    port map (
            O => \N__37561\,
            I => \N__37551\
        );

    \I__7979\ : CascadeMux
    port map (
            O => \N__37560\,
            I => \N__37547\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__37557\,
            I => \N__37544\
        );

    \I__7977\ : InMux
    port map (
            O => \N__37554\,
            I => \N__37541\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__37551\,
            I => \N__37538\
        );

    \I__7975\ : CascadeMux
    port map (
            O => \N__37550\,
            I => \N__37535\
        );

    \I__7974\ : InMux
    port map (
            O => \N__37547\,
            I => \N__37532\
        );

    \I__7973\ : Span4Mux_h
    port map (
            O => \N__37544\,
            I => \N__37527\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__37541\,
            I => \N__37527\
        );

    \I__7971\ : Span4Mux_h
    port map (
            O => \N__37538\,
            I => \N__37524\
        );

    \I__7970\ : InMux
    port map (
            O => \N__37535\,
            I => \N__37521\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__37532\,
            I => measured_delay_hc_13
        );

    \I__7968\ : Odrv4
    port map (
            O => \N__37527\,
            I => measured_delay_hc_13
        );

    \I__7967\ : Odrv4
    port map (
            O => \N__37524\,
            I => measured_delay_hc_13
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__37521\,
            I => measured_delay_hc_13
        );

    \I__7965\ : InMux
    port map (
            O => \N__37512\,
            I => \N__37499\
        );

    \I__7964\ : InMux
    port map (
            O => \N__37511\,
            I => \N__37499\
        );

    \I__7963\ : InMux
    port map (
            O => \N__37510\,
            I => \N__37499\
        );

    \I__7962\ : InMux
    port map (
            O => \N__37509\,
            I => \N__37499\
        );

    \I__7961\ : InMux
    port map (
            O => \N__37508\,
            I => \N__37496\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__37499\,
            I => \N__37492\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__37496\,
            I => \N__37489\
        );

    \I__7958\ : InMux
    port map (
            O => \N__37495\,
            I => \N__37486\
        );

    \I__7957\ : Span4Mux_v
    port map (
            O => \N__37492\,
            I => \N__37478\
        );

    \I__7956\ : Span4Mux_h
    port map (
            O => \N__37489\,
            I => \N__37478\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__37486\,
            I => \N__37478\
        );

    \I__7954\ : InMux
    port map (
            O => \N__37485\,
            I => \N__37475\
        );

    \I__7953\ : Span4Mux_h
    port map (
            O => \N__37478\,
            I => \N__37464\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__37475\,
            I => \N__37464\
        );

    \I__7951\ : InMux
    port map (
            O => \N__37474\,
            I => \N__37461\
        );

    \I__7950\ : InMux
    port map (
            O => \N__37473\,
            I => \N__37452\
        );

    \I__7949\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37452\
        );

    \I__7948\ : InMux
    port map (
            O => \N__37471\,
            I => \N__37452\
        );

    \I__7947\ : InMux
    port map (
            O => \N__37470\,
            I => \N__37452\
        );

    \I__7946\ : InMux
    port map (
            O => \N__37469\,
            I => \N__37449\
        );

    \I__7945\ : Odrv4
    port map (
            O => \N__37464\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__37461\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__37452\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__37449\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0\
        );

    \I__7941\ : CascadeMux
    port map (
            O => \N__37440\,
            I => \N__37433\
        );

    \I__7940\ : CascadeMux
    port map (
            O => \N__37439\,
            I => \N__37430\
        );

    \I__7939\ : CascadeMux
    port map (
            O => \N__37438\,
            I => \N__37425\
        );

    \I__7938\ : CascadeMux
    port map (
            O => \N__37437\,
            I => \N__37418\
        );

    \I__7937\ : CascadeMux
    port map (
            O => \N__37436\,
            I => \N__37413\
        );

    \I__7936\ : InMux
    port map (
            O => \N__37433\,
            I => \N__37402\
        );

    \I__7935\ : InMux
    port map (
            O => \N__37430\,
            I => \N__37402\
        );

    \I__7934\ : InMux
    port map (
            O => \N__37429\,
            I => \N__37402\
        );

    \I__7933\ : InMux
    port map (
            O => \N__37428\,
            I => \N__37389\
        );

    \I__7932\ : InMux
    port map (
            O => \N__37425\,
            I => \N__37389\
        );

    \I__7931\ : InMux
    port map (
            O => \N__37424\,
            I => \N__37389\
        );

    \I__7930\ : InMux
    port map (
            O => \N__37423\,
            I => \N__37389\
        );

    \I__7929\ : InMux
    port map (
            O => \N__37422\,
            I => \N__37389\
        );

    \I__7928\ : InMux
    port map (
            O => \N__37421\,
            I => \N__37389\
        );

    \I__7927\ : InMux
    port map (
            O => \N__37418\,
            I => \N__37378\
        );

    \I__7926\ : InMux
    port map (
            O => \N__37417\,
            I => \N__37378\
        );

    \I__7925\ : InMux
    port map (
            O => \N__37416\,
            I => \N__37378\
        );

    \I__7924\ : InMux
    port map (
            O => \N__37413\,
            I => \N__37378\
        );

    \I__7923\ : InMux
    port map (
            O => \N__37412\,
            I => \N__37378\
        );

    \I__7922\ : InMux
    port map (
            O => \N__37411\,
            I => \N__37375\
        );

    \I__7921\ : InMux
    port map (
            O => \N__37410\,
            I => \N__37368\
        );

    \I__7920\ : CascadeMux
    port map (
            O => \N__37409\,
            I => \N__37362\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__37402\,
            I => \N__37358\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__37389\,
            I => \N__37353\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__37378\,
            I => \N__37353\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__37375\,
            I => \N__37350\
        );

    \I__7915\ : InMux
    port map (
            O => \N__37374\,
            I => \N__37346\
        );

    \I__7914\ : InMux
    port map (
            O => \N__37373\,
            I => \N__37339\
        );

    \I__7913\ : InMux
    port map (
            O => \N__37372\,
            I => \N__37339\
        );

    \I__7912\ : InMux
    port map (
            O => \N__37371\,
            I => \N__37339\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__37368\,
            I => \N__37336\
        );

    \I__7910\ : CascadeMux
    port map (
            O => \N__37367\,
            I => \N__37333\
        );

    \I__7909\ : CascadeMux
    port map (
            O => \N__37366\,
            I => \N__37330\
        );

    \I__7908\ : CascadeMux
    port map (
            O => \N__37365\,
            I => \N__37325\
        );

    \I__7907\ : InMux
    port map (
            O => \N__37362\,
            I => \N__37318\
        );

    \I__7906\ : InMux
    port map (
            O => \N__37361\,
            I => \N__37315\
        );

    \I__7905\ : Span4Mux_v
    port map (
            O => \N__37358\,
            I => \N__37310\
        );

    \I__7904\ : Span4Mux_v
    port map (
            O => \N__37353\,
            I => \N__37310\
        );

    \I__7903\ : Span4Mux_h
    port map (
            O => \N__37350\,
            I => \N__37307\
        );

    \I__7902\ : InMux
    port map (
            O => \N__37349\,
            I => \N__37304\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__37346\,
            I => \N__37299\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__37339\,
            I => \N__37299\
        );

    \I__7899\ : Span4Mux_h
    port map (
            O => \N__37336\,
            I => \N__37296\
        );

    \I__7898\ : InMux
    port map (
            O => \N__37333\,
            I => \N__37293\
        );

    \I__7897\ : InMux
    port map (
            O => \N__37330\,
            I => \N__37288\
        );

    \I__7896\ : InMux
    port map (
            O => \N__37329\,
            I => \N__37288\
        );

    \I__7895\ : InMux
    port map (
            O => \N__37328\,
            I => \N__37275\
        );

    \I__7894\ : InMux
    port map (
            O => \N__37325\,
            I => \N__37275\
        );

    \I__7893\ : InMux
    port map (
            O => \N__37324\,
            I => \N__37275\
        );

    \I__7892\ : InMux
    port map (
            O => \N__37323\,
            I => \N__37275\
        );

    \I__7891\ : InMux
    port map (
            O => \N__37322\,
            I => \N__37275\
        );

    \I__7890\ : InMux
    port map (
            O => \N__37321\,
            I => \N__37275\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__37318\,
            I => \N__37270\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__37315\,
            I => \N__37270\
        );

    \I__7887\ : Span4Mux_h
    port map (
            O => \N__37310\,
            I => \N__37267\
        );

    \I__7886\ : Span4Mux_h
    port map (
            O => \N__37307\,
            I => \N__37264\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__37304\,
            I => \N__37257\
        );

    \I__7884\ : Span4Mux_h
    port map (
            O => \N__37299\,
            I => \N__37257\
        );

    \I__7883\ : Span4Mux_h
    port map (
            O => \N__37296\,
            I => \N__37257\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__37293\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__37288\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__37275\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7879\ : Odrv4
    port map (
            O => \N__37270\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7878\ : Odrv4
    port map (
            O => \N__37267\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7877\ : Odrv4
    port map (
            O => \N__37264\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7876\ : Odrv4
    port map (
            O => \N__37257\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7875\ : CascadeMux
    port map (
            O => \N__37242\,
            I => \N__37238\
        );

    \I__7874\ : CascadeMux
    port map (
            O => \N__37241\,
            I => \N__37235\
        );

    \I__7873\ : InMux
    port map (
            O => \N__37238\,
            I => \N__37230\
        );

    \I__7872\ : InMux
    port map (
            O => \N__37235\,
            I => \N__37227\
        );

    \I__7871\ : InMux
    port map (
            O => \N__37234\,
            I => \N__37224\
        );

    \I__7870\ : CascadeMux
    port map (
            O => \N__37233\,
            I => \N__37220\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__37230\,
            I => \N__37217\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__37227\,
            I => \N__37214\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__37224\,
            I => \N__37211\
        );

    \I__7866\ : InMux
    port map (
            O => \N__37223\,
            I => \N__37208\
        );

    \I__7865\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37205\
        );

    \I__7864\ : Span4Mux_h
    port map (
            O => \N__37217\,
            I => \N__37196\
        );

    \I__7863\ : Span4Mux_h
    port map (
            O => \N__37214\,
            I => \N__37196\
        );

    \I__7862\ : Span4Mux_v
    port map (
            O => \N__37211\,
            I => \N__37196\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__37208\,
            I => \N__37196\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__37205\,
            I => measured_delay_hc_7
        );

    \I__7859\ : Odrv4
    port map (
            O => \N__37196\,
            I => measured_delay_hc_7
        );

    \I__7858\ : InMux
    port map (
            O => \N__37191\,
            I => \N__37181\
        );

    \I__7857\ : InMux
    port map (
            O => \N__37190\,
            I => \N__37181\
        );

    \I__7856\ : InMux
    port map (
            O => \N__37189\,
            I => \N__37176\
        );

    \I__7855\ : InMux
    port map (
            O => \N__37188\,
            I => \N__37176\
        );

    \I__7854\ : InMux
    port map (
            O => \N__37187\,
            I => \N__37173\
        );

    \I__7853\ : InMux
    port map (
            O => \N__37186\,
            I => \N__37170\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__37181\,
            I => \N__37163\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__37176\,
            I => \N__37163\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__37173\,
            I => \N__37163\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__37170\,
            I => \N__37157\
        );

    \I__7848\ : Span4Mux_v
    port map (
            O => \N__37163\,
            I => \N__37150\
        );

    \I__7847\ : InMux
    port map (
            O => \N__37162\,
            I => \N__37145\
        );

    \I__7846\ : InMux
    port map (
            O => \N__37161\,
            I => \N__37145\
        );

    \I__7845\ : InMux
    port map (
            O => \N__37160\,
            I => \N__37142\
        );

    \I__7844\ : Span4Mux_v
    port map (
            O => \N__37157\,
            I => \N__37138\
        );

    \I__7843\ : InMux
    port map (
            O => \N__37156\,
            I => \N__37133\
        );

    \I__7842\ : InMux
    port map (
            O => \N__37155\,
            I => \N__37133\
        );

    \I__7841\ : InMux
    port map (
            O => \N__37154\,
            I => \N__37128\
        );

    \I__7840\ : InMux
    port map (
            O => \N__37153\,
            I => \N__37128\
        );

    \I__7839\ : Span4Mux_h
    port map (
            O => \N__37150\,
            I => \N__37121\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__37145\,
            I => \N__37121\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__37142\,
            I => \N__37121\
        );

    \I__7836\ : InMux
    port map (
            O => \N__37141\,
            I => \N__37118\
        );

    \I__7835\ : Odrv4
    port map (
            O => \N__37138\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__37133\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__37128\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0\
        );

    \I__7832\ : Odrv4
    port map (
            O => \N__37121\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__37118\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0\
        );

    \I__7830\ : CEMux
    port map (
            O => \N__37107\,
            I => \N__37103\
        );

    \I__7829\ : CEMux
    port map (
            O => \N__37106\,
            I => \N__37100\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__37103\,
            I => \N__37096\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__37100\,
            I => \N__37093\
        );

    \I__7826\ : CEMux
    port map (
            O => \N__37099\,
            I => \N__37088\
        );

    \I__7825\ : Span4Mux_v
    port map (
            O => \N__37096\,
            I => \N__37083\
        );

    \I__7824\ : Span4Mux_v
    port map (
            O => \N__37093\,
            I => \N__37083\
        );

    \I__7823\ : CEMux
    port map (
            O => \N__37092\,
            I => \N__37080\
        );

    \I__7822\ : CEMux
    port map (
            O => \N__37091\,
            I => \N__37077\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__37088\,
            I => \N__37074\
        );

    \I__7820\ : Span4Mux_h
    port map (
            O => \N__37083\,
            I => \N__37071\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__37080\,
            I => \N__37068\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__37077\,
            I => \N__37065\
        );

    \I__7817\ : Span4Mux_v
    port map (
            O => \N__37074\,
            I => \N__37062\
        );

    \I__7816\ : Span4Mux_h
    port map (
            O => \N__37071\,
            I => \N__37057\
        );

    \I__7815\ : Span4Mux_v
    port map (
            O => \N__37068\,
            I => \N__37057\
        );

    \I__7814\ : Span4Mux_v
    port map (
            O => \N__37065\,
            I => \N__37052\
        );

    \I__7813\ : Span4Mux_v
    port map (
            O => \N__37062\,
            I => \N__37052\
        );

    \I__7812\ : Odrv4
    port map (
            O => \N__37057\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__7811\ : Odrv4
    port map (
            O => \N__37052\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__7810\ : InMux
    port map (
            O => \N__37047\,
            I => \N__37043\
        );

    \I__7809\ : InMux
    port map (
            O => \N__37046\,
            I => \N__37039\
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__37043\,
            I => \N__37033\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37042\,
            I => \N__37030\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__37039\,
            I => \N__37027\
        );

    \I__7805\ : InMux
    port map (
            O => \N__37038\,
            I => \N__37024\
        );

    \I__7804\ : InMux
    port map (
            O => \N__37037\,
            I => \N__37021\
        );

    \I__7803\ : InMux
    port map (
            O => \N__37036\,
            I => \N__37018\
        );

    \I__7802\ : Span4Mux_h
    port map (
            O => \N__37033\,
            I => \N__37013\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__37030\,
            I => \N__37013\
        );

    \I__7800\ : Span12Mux_s8_v
    port map (
            O => \N__37027\,
            I => \N__37010\
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__37024\,
            I => \N__37007\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__37021\,
            I => \N__37004\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__37018\,
            I => measured_delay_hc_9
        );

    \I__7796\ : Odrv4
    port map (
            O => \N__37013\,
            I => measured_delay_hc_9
        );

    \I__7795\ : Odrv12
    port map (
            O => \N__37010\,
            I => measured_delay_hc_9
        );

    \I__7794\ : Odrv12
    port map (
            O => \N__37007\,
            I => measured_delay_hc_9
        );

    \I__7793\ : Odrv4
    port map (
            O => \N__37004\,
            I => measured_delay_hc_9
        );

    \I__7792\ : CascadeMux
    port map (
            O => \N__36993\,
            I => \N__36989\
        );

    \I__7791\ : InMux
    port map (
            O => \N__36992\,
            I => \N__36986\
        );

    \I__7790\ : InMux
    port map (
            O => \N__36989\,
            I => \N__36982\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__36986\,
            I => \N__36979\
        );

    \I__7788\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36975\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__36982\,
            I => \N__36972\
        );

    \I__7786\ : Span4Mux_h
    port map (
            O => \N__36979\,
            I => \N__36969\
        );

    \I__7785\ : InMux
    port map (
            O => \N__36978\,
            I => \N__36966\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__36975\,
            I => measured_delay_hc_0
        );

    \I__7783\ : Odrv12
    port map (
            O => \N__36972\,
            I => measured_delay_hc_0
        );

    \I__7782\ : Odrv4
    port map (
            O => \N__36969\,
            I => measured_delay_hc_0
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__36966\,
            I => measured_delay_hc_0
        );

    \I__7780\ : InMux
    port map (
            O => \N__36957\,
            I => \N__36952\
        );

    \I__7779\ : CascadeMux
    port map (
            O => \N__36956\,
            I => \N__36948\
        );

    \I__7778\ : CascadeMux
    port map (
            O => \N__36955\,
            I => \N__36945\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__36952\,
            I => \N__36942\
        );

    \I__7776\ : InMux
    port map (
            O => \N__36951\,
            I => \N__36939\
        );

    \I__7775\ : InMux
    port map (
            O => \N__36948\,
            I => \N__36935\
        );

    \I__7774\ : InMux
    port map (
            O => \N__36945\,
            I => \N__36932\
        );

    \I__7773\ : Span4Mux_h
    port map (
            O => \N__36942\,
            I => \N__36927\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__36939\,
            I => \N__36927\
        );

    \I__7771\ : InMux
    port map (
            O => \N__36938\,
            I => \N__36924\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__36935\,
            I => measured_delay_hc_6
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__36932\,
            I => measured_delay_hc_6
        );

    \I__7768\ : Odrv4
    port map (
            O => \N__36927\,
            I => measured_delay_hc_6
        );

    \I__7767\ : LocalMux
    port map (
            O => \N__36924\,
            I => measured_delay_hc_6
        );

    \I__7766\ : InMux
    port map (
            O => \N__36915\,
            I => \N__36910\
        );

    \I__7765\ : InMux
    port map (
            O => \N__36914\,
            I => \N__36906\
        );

    \I__7764\ : InMux
    port map (
            O => \N__36913\,
            I => \N__36903\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__36910\,
            I => \N__36900\
        );

    \I__7762\ : InMux
    port map (
            O => \N__36909\,
            I => \N__36896\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__36906\,
            I => \N__36893\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__36903\,
            I => \N__36888\
        );

    \I__7759\ : Span4Mux_v
    port map (
            O => \N__36900\,
            I => \N__36888\
        );

    \I__7758\ : InMux
    port map (
            O => \N__36899\,
            I => \N__36885\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__36896\,
            I => measured_delay_hc_1
        );

    \I__7756\ : Odrv12
    port map (
            O => \N__36893\,
            I => measured_delay_hc_1
        );

    \I__7755\ : Odrv4
    port map (
            O => \N__36888\,
            I => measured_delay_hc_1
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__36885\,
            I => measured_delay_hc_1
        );

    \I__7753\ : InMux
    port map (
            O => \N__36876\,
            I => \N__36872\
        );

    \I__7752\ : InMux
    port map (
            O => \N__36875\,
            I => \N__36868\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__36872\,
            I => \N__36864\
        );

    \I__7750\ : InMux
    port map (
            O => \N__36871\,
            I => \N__36861\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__36868\,
            I => \N__36858\
        );

    \I__7748\ : InMux
    port map (
            O => \N__36867\,
            I => \N__36854\
        );

    \I__7747\ : Span4Mux_v
    port map (
            O => \N__36864\,
            I => \N__36851\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__36861\,
            I => \N__36848\
        );

    \I__7745\ : Span4Mux_v
    port map (
            O => \N__36858\,
            I => \N__36845\
        );

    \I__7744\ : InMux
    port map (
            O => \N__36857\,
            I => \N__36842\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__36854\,
            I => measured_delay_hc_3
        );

    \I__7742\ : Odrv4
    port map (
            O => \N__36851\,
            I => measured_delay_hc_3
        );

    \I__7741\ : Odrv12
    port map (
            O => \N__36848\,
            I => measured_delay_hc_3
        );

    \I__7740\ : Odrv4
    port map (
            O => \N__36845\,
            I => measured_delay_hc_3
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__36842\,
            I => measured_delay_hc_3
        );

    \I__7738\ : InMux
    port map (
            O => \N__36831\,
            I => \N__36828\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__36828\,
            I => \N__36821\
        );

    \I__7736\ : InMux
    port map (
            O => \N__36827\,
            I => \N__36818\
        );

    \I__7735\ : InMux
    port map (
            O => \N__36826\,
            I => \N__36815\
        );

    \I__7734\ : InMux
    port map (
            O => \N__36825\,
            I => \N__36812\
        );

    \I__7733\ : InMux
    port map (
            O => \N__36824\,
            I => \N__36809\
        );

    \I__7732\ : Span12Mux_s8_v
    port map (
            O => \N__36821\,
            I => \N__36804\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__36818\,
            I => \N__36804\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__36815\,
            I => \N__36801\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__36812\,
            I => measured_delay_hc_4
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__36809\,
            I => measured_delay_hc_4
        );

    \I__7727\ : Odrv12
    port map (
            O => \N__36804\,
            I => measured_delay_hc_4
        );

    \I__7726\ : Odrv4
    port map (
            O => \N__36801\,
            I => measured_delay_hc_4
        );

    \I__7725\ : InMux
    port map (
            O => \N__36792\,
            I => \N__36788\
        );

    \I__7724\ : InMux
    port map (
            O => \N__36791\,
            I => \N__36785\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__36788\,
            I => \N__36779\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__36785\,
            I => \N__36779\
        );

    \I__7721\ : InMux
    port map (
            O => \N__36784\,
            I => \N__36776\
        );

    \I__7720\ : Span4Mux_v
    port map (
            O => \N__36779\,
            I => \N__36769\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__36776\,
            I => \N__36769\
        );

    \I__7718\ : InMux
    port map (
            O => \N__36775\,
            I => \N__36766\
        );

    \I__7717\ : InMux
    port map (
            O => \N__36774\,
            I => \N__36763\
        );

    \I__7716\ : Span4Mux_h
    port map (
            O => \N__36769\,
            I => \N__36760\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__36766\,
            I => measured_delay_hc_16
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__36763\,
            I => measured_delay_hc_16
        );

    \I__7713\ : Odrv4
    port map (
            O => \N__36760\,
            I => measured_delay_hc_16
        );

    \I__7712\ : InMux
    port map (
            O => \N__36753\,
            I => \N__36746\
        );

    \I__7711\ : InMux
    port map (
            O => \N__36752\,
            I => \N__36743\
        );

    \I__7710\ : InMux
    port map (
            O => \N__36751\,
            I => \N__36740\
        );

    \I__7709\ : CascadeMux
    port map (
            O => \N__36750\,
            I => \N__36737\
        );

    \I__7708\ : InMux
    port map (
            O => \N__36749\,
            I => \N__36734\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__36746\,
            I => \N__36731\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__36743\,
            I => \N__36728\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__36740\,
            I => \N__36725\
        );

    \I__7704\ : InMux
    port map (
            O => \N__36737\,
            I => \N__36722\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__36734\,
            I => \N__36719\
        );

    \I__7702\ : Span4Mux_h
    port map (
            O => \N__36731\,
            I => \N__36716\
        );

    \I__7701\ : Span4Mux_h
    port map (
            O => \N__36728\,
            I => \N__36711\
        );

    \I__7700\ : Span4Mux_h
    port map (
            O => \N__36725\,
            I => \N__36711\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__36722\,
            I => measured_delay_hc_14
        );

    \I__7698\ : Odrv4
    port map (
            O => \N__36719\,
            I => measured_delay_hc_14
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__36716\,
            I => measured_delay_hc_14
        );

    \I__7696\ : Odrv4
    port map (
            O => \N__36711\,
            I => measured_delay_hc_14
        );

    \I__7695\ : InMux
    port map (
            O => \N__36702\,
            I => \N__36698\
        );

    \I__7694\ : InMux
    port map (
            O => \N__36701\,
            I => \N__36694\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__36698\,
            I => \N__36690\
        );

    \I__7692\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36687\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__36694\,
            I => \N__36684\
        );

    \I__7690\ : InMux
    port map (
            O => \N__36693\,
            I => \N__36680\
        );

    \I__7689\ : Span4Mux_h
    port map (
            O => \N__36690\,
            I => \N__36675\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__36687\,
            I => \N__36675\
        );

    \I__7687\ : Span4Mux_v
    port map (
            O => \N__36684\,
            I => \N__36672\
        );

    \I__7686\ : InMux
    port map (
            O => \N__36683\,
            I => \N__36669\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__36680\,
            I => measured_delay_hc_10
        );

    \I__7684\ : Odrv4
    port map (
            O => \N__36675\,
            I => measured_delay_hc_10
        );

    \I__7683\ : Odrv4
    port map (
            O => \N__36672\,
            I => measured_delay_hc_10
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__36669\,
            I => measured_delay_hc_10
        );

    \I__7681\ : CascadeMux
    port map (
            O => \N__36660\,
            I => \N__36657\
        );

    \I__7680\ : InMux
    port map (
            O => \N__36657\,
            I => \N__36652\
        );

    \I__7679\ : InMux
    port map (
            O => \N__36656\,
            I => \N__36649\
        );

    \I__7678\ : InMux
    port map (
            O => \N__36655\,
            I => \N__36645\
        );

    \I__7677\ : LocalMux
    port map (
            O => \N__36652\,
            I => \N__36640\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__36649\,
            I => \N__36640\
        );

    \I__7675\ : CascadeMux
    port map (
            O => \N__36648\,
            I => \N__36637\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__36645\,
            I => \N__36634\
        );

    \I__7673\ : Span4Mux_v
    port map (
            O => \N__36640\,
            I => \N__36631\
        );

    \I__7672\ : InMux
    port map (
            O => \N__36637\,
            I => \N__36627\
        );

    \I__7671\ : Span12Mux_h
    port map (
            O => \N__36634\,
            I => \N__36624\
        );

    \I__7670\ : Span4Mux_h
    port map (
            O => \N__36631\,
            I => \N__36621\
        );

    \I__7669\ : InMux
    port map (
            O => \N__36630\,
            I => \N__36618\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__36627\,
            I => measured_delay_hc_11
        );

    \I__7667\ : Odrv12
    port map (
            O => \N__36624\,
            I => measured_delay_hc_11
        );

    \I__7666\ : Odrv4
    port map (
            O => \N__36621\,
            I => measured_delay_hc_11
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__36618\,
            I => measured_delay_hc_11
        );

    \I__7664\ : InMux
    port map (
            O => \N__36609\,
            I => \N__36603\
        );

    \I__7663\ : CascadeMux
    port map (
            O => \N__36608\,
            I => \N__36600\
        );

    \I__7662\ : InMux
    port map (
            O => \N__36607\,
            I => \N__36597\
        );

    \I__7661\ : InMux
    port map (
            O => \N__36606\,
            I => \N__36594\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__36603\,
            I => \N__36591\
        );

    \I__7659\ : InMux
    port map (
            O => \N__36600\,
            I => \N__36587\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__36597\,
            I => \N__36584\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__36594\,
            I => \N__36581\
        );

    \I__7656\ : Span4Mux_h
    port map (
            O => \N__36591\,
            I => \N__36578\
        );

    \I__7655\ : InMux
    port map (
            O => \N__36590\,
            I => \N__36575\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__36587\,
            I => measured_delay_hc_12
        );

    \I__7653\ : Odrv4
    port map (
            O => \N__36584\,
            I => measured_delay_hc_12
        );

    \I__7652\ : Odrv12
    port map (
            O => \N__36581\,
            I => measured_delay_hc_12
        );

    \I__7651\ : Odrv4
    port map (
            O => \N__36578\,
            I => measured_delay_hc_12
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__36575\,
            I => measured_delay_hc_12
        );

    \I__7649\ : InMux
    port map (
            O => \N__36564\,
            I => \N__36559\
        );

    \I__7648\ : InMux
    port map (
            O => \N__36563\,
            I => \N__36555\
        );

    \I__7647\ : InMux
    port map (
            O => \N__36562\,
            I => \N__36552\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__36559\,
            I => \N__36548\
        );

    \I__7645\ : InMux
    port map (
            O => \N__36558\,
            I => \N__36545\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__36555\,
            I => \N__36540\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__36552\,
            I => \N__36540\
        );

    \I__7642\ : CascadeMux
    port map (
            O => \N__36551\,
            I => \N__36537\
        );

    \I__7641\ : Span4Mux_h
    port map (
            O => \N__36548\,
            I => \N__36532\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__36545\,
            I => \N__36532\
        );

    \I__7639\ : Span4Mux_v
    port map (
            O => \N__36540\,
            I => \N__36529\
        );

    \I__7638\ : InMux
    port map (
            O => \N__36537\,
            I => \N__36526\
        );

    \I__7637\ : Span4Mux_v
    port map (
            O => \N__36532\,
            I => \N__36521\
        );

    \I__7636\ : Span4Mux_h
    port map (
            O => \N__36529\,
            I => \N__36521\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__36526\,
            I => measured_delay_hc_19
        );

    \I__7634\ : Odrv4
    port map (
            O => \N__36521\,
            I => measured_delay_hc_19
        );

    \I__7633\ : CascadeMux
    port map (
            O => \N__36516\,
            I => \N__36513\
        );

    \I__7632\ : InMux
    port map (
            O => \N__36513\,
            I => \N__36509\
        );

    \I__7631\ : CascadeMux
    port map (
            O => \N__36512\,
            I => \N__36505\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__36509\,
            I => \N__36502\
        );

    \I__7629\ : InMux
    port map (
            O => \N__36508\,
            I => \N__36497\
        );

    \I__7628\ : InMux
    port map (
            O => \N__36505\,
            I => \N__36494\
        );

    \I__7627\ : Span4Mux_h
    port map (
            O => \N__36502\,
            I => \N__36491\
        );

    \I__7626\ : InMux
    port map (
            O => \N__36501\,
            I => \N__36488\
        );

    \I__7625\ : InMux
    port map (
            O => \N__36500\,
            I => \N__36485\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__36497\,
            I => \N__36480\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__36494\,
            I => \N__36480\
        );

    \I__7622\ : Span4Mux_h
    port map (
            O => \N__36491\,
            I => \N__36477\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__36488\,
            I => measured_delay_hc_17
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__36485\,
            I => measured_delay_hc_17
        );

    \I__7619\ : Odrv12
    port map (
            O => \N__36480\,
            I => measured_delay_hc_17
        );

    \I__7618\ : Odrv4
    port map (
            O => \N__36477\,
            I => measured_delay_hc_17
        );

    \I__7617\ : InMux
    port map (
            O => \N__36468\,
            I => \N__36465\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__36465\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\
        );

    \I__7615\ : InMux
    port map (
            O => \N__36462\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__7614\ : InMux
    port map (
            O => \N__36459\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__7613\ : CascadeMux
    port map (
            O => \N__36456\,
            I => \N__36449\
        );

    \I__7612\ : CascadeMux
    port map (
            O => \N__36455\,
            I => \N__36443\
        );

    \I__7611\ : CascadeMux
    port map (
            O => \N__36454\,
            I => \N__36440\
        );

    \I__7610\ : InMux
    port map (
            O => \N__36453\,
            I => \N__36416\
        );

    \I__7609\ : InMux
    port map (
            O => \N__36452\,
            I => \N__36416\
        );

    \I__7608\ : InMux
    port map (
            O => \N__36449\,
            I => \N__36416\
        );

    \I__7607\ : InMux
    port map (
            O => \N__36448\,
            I => \N__36416\
        );

    \I__7606\ : InMux
    port map (
            O => \N__36447\,
            I => \N__36416\
        );

    \I__7605\ : InMux
    port map (
            O => \N__36446\,
            I => \N__36416\
        );

    \I__7604\ : InMux
    port map (
            O => \N__36443\,
            I => \N__36405\
        );

    \I__7603\ : InMux
    port map (
            O => \N__36440\,
            I => \N__36405\
        );

    \I__7602\ : InMux
    port map (
            O => \N__36439\,
            I => \N__36405\
        );

    \I__7601\ : InMux
    port map (
            O => \N__36438\,
            I => \N__36405\
        );

    \I__7600\ : InMux
    port map (
            O => \N__36437\,
            I => \N__36405\
        );

    \I__7599\ : InMux
    port map (
            O => \N__36436\,
            I => \N__36400\
        );

    \I__7598\ : InMux
    port map (
            O => \N__36435\,
            I => \N__36400\
        );

    \I__7597\ : InMux
    port map (
            O => \N__36434\,
            I => \N__36395\
        );

    \I__7596\ : InMux
    port map (
            O => \N__36433\,
            I => \N__36395\
        );

    \I__7595\ : InMux
    port map (
            O => \N__36432\,
            I => \N__36392\
        );

    \I__7594\ : InMux
    port map (
            O => \N__36431\,
            I => \N__36385\
        );

    \I__7593\ : InMux
    port map (
            O => \N__36430\,
            I => \N__36385\
        );

    \I__7592\ : InMux
    port map (
            O => \N__36429\,
            I => \N__36385\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__36416\,
            I => \N__36376\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__36405\,
            I => \N__36376\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__36400\,
            I => \N__36376\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__36395\,
            I => \N__36376\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__36392\,
            I => \N__36369\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__36385\,
            I => \N__36369\
        );

    \I__7585\ : Span4Mux_v
    port map (
            O => \N__36376\,
            I => \N__36369\
        );

    \I__7584\ : Odrv4
    port map (
            O => \N__36369\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__7583\ : CEMux
    port map (
            O => \N__36366\,
            I => \N__36362\
        );

    \I__7582\ : CEMux
    port map (
            O => \N__36365\,
            I => \N__36359\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__36362\,
            I => \N__36356\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__36359\,
            I => \N__36352\
        );

    \I__7579\ : Span4Mux_v
    port map (
            O => \N__36356\,
            I => \N__36349\
        );

    \I__7578\ : CEMux
    port map (
            O => \N__36355\,
            I => \N__36344\
        );

    \I__7577\ : Span4Mux_h
    port map (
            O => \N__36352\,
            I => \N__36341\
        );

    \I__7576\ : Span4Mux_h
    port map (
            O => \N__36349\,
            I => \N__36338\
        );

    \I__7575\ : CEMux
    port map (
            O => \N__36348\,
            I => \N__36335\
        );

    \I__7574\ : CEMux
    port map (
            O => \N__36347\,
            I => \N__36332\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__36344\,
            I => \N__36329\
        );

    \I__7572\ : Odrv4
    port map (
            O => \N__36341\,
            I => \delay_measurement_inst.delay_tr_timer.N_337_i\
        );

    \I__7571\ : Odrv4
    port map (
            O => \N__36338\,
            I => \delay_measurement_inst.delay_tr_timer.N_337_i\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__36335\,
            I => \delay_measurement_inst.delay_tr_timer.N_337_i\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__36332\,
            I => \delay_measurement_inst.delay_tr_timer.N_337_i\
        );

    \I__7568\ : Odrv4
    port map (
            O => \N__36329\,
            I => \delay_measurement_inst.delay_tr_timer.N_337_i\
        );

    \I__7567\ : InMux
    port map (
            O => \N__36318\,
            I => \N__36315\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__36315\,
            I => \N__36312\
        );

    \I__7565\ : Odrv4
    port map (
            O => \N__36312\,
            I => delay_tr_input_c
        );

    \I__7564\ : InMux
    port map (
            O => \N__36309\,
            I => \N__36306\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__36306\,
            I => delay_tr_d1
        );

    \I__7562\ : InMux
    port map (
            O => \N__36303\,
            I => \N__36298\
        );

    \I__7561\ : InMux
    port map (
            O => \N__36302\,
            I => \N__36295\
        );

    \I__7560\ : InMux
    port map (
            O => \N__36301\,
            I => \N__36292\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__36298\,
            I => \N__36288\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__36295\,
            I => \N__36285\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__36292\,
            I => \N__36282\
        );

    \I__7556\ : InMux
    port map (
            O => \N__36291\,
            I => \N__36279\
        );

    \I__7555\ : Span4Mux_v
    port map (
            O => \N__36288\,
            I => \N__36272\
        );

    \I__7554\ : Span4Mux_h
    port map (
            O => \N__36285\,
            I => \N__36272\
        );

    \I__7553\ : Span4Mux_v
    port map (
            O => \N__36282\,
            I => \N__36272\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__36279\,
            I => \N__36269\
        );

    \I__7551\ : Sp12to4
    port map (
            O => \N__36272\,
            I => \N__36264\
        );

    \I__7550\ : Span12Mux_h
    port map (
            O => \N__36269\,
            I => \N__36264\
        );

    \I__7549\ : Odrv12
    port map (
            O => \N__36264\,
            I => delay_tr_d2
        );

    \I__7548\ : InMux
    port map (
            O => \N__36261\,
            I => \N__36258\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__36258\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__7546\ : InMux
    port map (
            O => \N__36255\,
            I => \N__36252\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__36252\,
            I => \N__36249\
        );

    \I__7544\ : Odrv4
    port map (
            O => \N__36249\,
            I => \phase_controller_inst1.N_228\
        );

    \I__7543\ : CascadeMux
    port map (
            O => \N__36246\,
            I => \N__36231\
        );

    \I__7542\ : CascadeMux
    port map (
            O => \N__36245\,
            I => \N__36224\
        );

    \I__7541\ : CascadeMux
    port map (
            O => \N__36244\,
            I => \N__36221\
        );

    \I__7540\ : CascadeMux
    port map (
            O => \N__36243\,
            I => \N__36218\
        );

    \I__7539\ : CascadeMux
    port map (
            O => \N__36242\,
            I => \N__36215\
        );

    \I__7538\ : InMux
    port map (
            O => \N__36241\,
            I => \N__36212\
        );

    \I__7537\ : CascadeMux
    port map (
            O => \N__36240\,
            I => \N__36209\
        );

    \I__7536\ : CascadeMux
    port map (
            O => \N__36239\,
            I => \N__36206\
        );

    \I__7535\ : CascadeMux
    port map (
            O => \N__36238\,
            I => \N__36203\
        );

    \I__7534\ : CascadeMux
    port map (
            O => \N__36237\,
            I => \N__36194\
        );

    \I__7533\ : CascadeMux
    port map (
            O => \N__36236\,
            I => \N__36191\
        );

    \I__7532\ : CascadeMux
    port map (
            O => \N__36235\,
            I => \N__36188\
        );

    \I__7531\ : CascadeMux
    port map (
            O => \N__36234\,
            I => \N__36185\
        );

    \I__7530\ : InMux
    port map (
            O => \N__36231\,
            I => \N__36182\
        );

    \I__7529\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36179\
        );

    \I__7528\ : InMux
    port map (
            O => \N__36229\,
            I => \N__36163\
        );

    \I__7527\ : InMux
    port map (
            O => \N__36228\,
            I => \N__36163\
        );

    \I__7526\ : InMux
    port map (
            O => \N__36227\,
            I => \N__36163\
        );

    \I__7525\ : InMux
    port map (
            O => \N__36224\,
            I => \N__36163\
        );

    \I__7524\ : InMux
    port map (
            O => \N__36221\,
            I => \N__36163\
        );

    \I__7523\ : InMux
    port map (
            O => \N__36218\,
            I => \N__36163\
        );

    \I__7522\ : InMux
    port map (
            O => \N__36215\,
            I => \N__36163\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__36212\,
            I => \N__36160\
        );

    \I__7520\ : InMux
    port map (
            O => \N__36209\,
            I => \N__36157\
        );

    \I__7519\ : InMux
    port map (
            O => \N__36206\,
            I => \N__36146\
        );

    \I__7518\ : InMux
    port map (
            O => \N__36203\,
            I => \N__36146\
        );

    \I__7517\ : InMux
    port map (
            O => \N__36202\,
            I => \N__36146\
        );

    \I__7516\ : InMux
    port map (
            O => \N__36201\,
            I => \N__36146\
        );

    \I__7515\ : InMux
    port map (
            O => \N__36200\,
            I => \N__36146\
        );

    \I__7514\ : InMux
    port map (
            O => \N__36199\,
            I => \N__36131\
        );

    \I__7513\ : InMux
    port map (
            O => \N__36198\,
            I => \N__36131\
        );

    \I__7512\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36131\
        );

    \I__7511\ : InMux
    port map (
            O => \N__36194\,
            I => \N__36131\
        );

    \I__7510\ : InMux
    port map (
            O => \N__36191\,
            I => \N__36131\
        );

    \I__7509\ : InMux
    port map (
            O => \N__36188\,
            I => \N__36131\
        );

    \I__7508\ : InMux
    port map (
            O => \N__36185\,
            I => \N__36131\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__36182\,
            I => \N__36128\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__36179\,
            I => \N__36125\
        );

    \I__7505\ : CascadeMux
    port map (
            O => \N__36178\,
            I => \N__36122\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__36163\,
            I => \N__36119\
        );

    \I__7503\ : Span4Mux_v
    port map (
            O => \N__36160\,
            I => \N__36116\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__36157\,
            I => \N__36105\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__36146\,
            I => \N__36105\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__36131\,
            I => \N__36105\
        );

    \I__7499\ : Span4Mux_v
    port map (
            O => \N__36128\,
            I => \N__36105\
        );

    \I__7498\ : Span4Mux_h
    port map (
            O => \N__36125\,
            I => \N__36105\
        );

    \I__7497\ : InMux
    port map (
            O => \N__36122\,
            I => \N__36102\
        );

    \I__7496\ : Span4Mux_h
    port map (
            O => \N__36119\,
            I => \N__36099\
        );

    \I__7495\ : Span4Mux_h
    port map (
            O => \N__36116\,
            I => \N__36096\
        );

    \I__7494\ : Span4Mux_v
    port map (
            O => \N__36105\,
            I => \N__36093\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__36102\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7492\ : Odrv4
    port map (
            O => \N__36099\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7491\ : Odrv4
    port map (
            O => \N__36096\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7490\ : Odrv4
    port map (
            O => \N__36093\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7489\ : InMux
    port map (
            O => \N__36084\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__7488\ : InMux
    port map (
            O => \N__36081\,
            I => \N__36078\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__36078\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__7486\ : InMux
    port map (
            O => \N__36075\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__7485\ : InMux
    port map (
            O => \N__36072\,
            I => \N__36069\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__36069\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__7483\ : InMux
    port map (
            O => \N__36066\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__7482\ : CascadeMux
    port map (
            O => \N__36063\,
            I => \N__36060\
        );

    \I__7481\ : InMux
    port map (
            O => \N__36060\,
            I => \N__36057\
        );

    \I__7480\ : LocalMux
    port map (
            O => \N__36057\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36054\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__7478\ : InMux
    port map (
            O => \N__36051\,
            I => \N__36048\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__36048\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__7476\ : InMux
    port map (
            O => \N__36045\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__7475\ : InMux
    port map (
            O => \N__36042\,
            I => \N__36039\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__36039\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__7473\ : InMux
    port map (
            O => \N__36036\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__7472\ : InMux
    port map (
            O => \N__36033\,
            I => \N__36030\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__36030\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__7470\ : InMux
    port map (
            O => \N__36027\,
            I => \bfn_14_23_0_\
        );

    \I__7469\ : CascadeMux
    port map (
            O => \N__36024\,
            I => \N__36021\
        );

    \I__7468\ : InMux
    port map (
            O => \N__36021\,
            I => \N__36018\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__36018\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__7466\ : InMux
    port map (
            O => \N__36015\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__7465\ : InMux
    port map (
            O => \N__36012\,
            I => \N__36009\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__36009\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__7463\ : InMux
    port map (
            O => \N__36006\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__7462\ : InMux
    port map (
            O => \N__36003\,
            I => \N__35999\
        );

    \I__7461\ : CascadeMux
    port map (
            O => \N__36002\,
            I => \N__35996\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__35999\,
            I => \N__35993\
        );

    \I__7459\ : InMux
    port map (
            O => \N__35996\,
            I => \N__35990\
        );

    \I__7458\ : Span4Mux_v
    port map (
            O => \N__35993\,
            I => \N__35987\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__35990\,
            I => \N__35984\
        );

    \I__7456\ : Odrv4
    port map (
            O => \N__35987\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__7455\ : Odrv4
    port map (
            O => \N__35984\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__7454\ : InMux
    port map (
            O => \N__35979\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__7453\ : InMux
    port map (
            O => \N__35976\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__7452\ : InMux
    port map (
            O => \N__35973\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__7451\ : InMux
    port map (
            O => \N__35970\,
            I => \N__35967\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__35967\,
            I => \N__35962\
        );

    \I__7449\ : InMux
    port map (
            O => \N__35966\,
            I => \N__35959\
        );

    \I__7448\ : InMux
    port map (
            O => \N__35965\,
            I => \N__35956\
        );

    \I__7447\ : Span4Mux_h
    port map (
            O => \N__35962\,
            I => \N__35951\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__35959\,
            I => \N__35951\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__35956\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__7444\ : Odrv4
    port map (
            O => \N__35951\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__7443\ : InMux
    port map (
            O => \N__35946\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__7442\ : CascadeMux
    port map (
            O => \N__35943\,
            I => \N__35939\
        );

    \I__7441\ : InMux
    port map (
            O => \N__35942\,
            I => \N__35936\
        );

    \I__7440\ : InMux
    port map (
            O => \N__35939\,
            I => \N__35933\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__35936\,
            I => \N__35929\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__35933\,
            I => \N__35926\
        );

    \I__7437\ : InMux
    port map (
            O => \N__35932\,
            I => \N__35923\
        );

    \I__7436\ : Span4Mux_v
    port map (
            O => \N__35929\,
            I => \N__35920\
        );

    \I__7435\ : Span4Mux_h
    port map (
            O => \N__35926\,
            I => \N__35917\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__35923\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__7433\ : Odrv4
    port map (
            O => \N__35920\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__7432\ : Odrv4
    port map (
            O => \N__35917\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__7431\ : InMux
    port map (
            O => \N__35910\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__7430\ : InMux
    port map (
            O => \N__35907\,
            I => \N__35901\
        );

    \I__7429\ : InMux
    port map (
            O => \N__35906\,
            I => \N__35901\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__35901\,
            I => \N__35897\
        );

    \I__7427\ : InMux
    port map (
            O => \N__35900\,
            I => \N__35894\
        );

    \I__7426\ : Span4Mux_h
    port map (
            O => \N__35897\,
            I => \N__35891\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__35894\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__7424\ : Odrv4
    port map (
            O => \N__35891\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__7423\ : InMux
    port map (
            O => \N__35886\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__7422\ : CascadeMux
    port map (
            O => \N__35883\,
            I => \N__35879\
        );

    \I__7421\ : InMux
    port map (
            O => \N__35882\,
            I => \N__35873\
        );

    \I__7420\ : InMux
    port map (
            O => \N__35879\,
            I => \N__35873\
        );

    \I__7419\ : InMux
    port map (
            O => \N__35878\,
            I => \N__35870\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__35873\,
            I => \N__35867\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__35870\,
            I => \N__35862\
        );

    \I__7416\ : Span4Mux_h
    port map (
            O => \N__35867\,
            I => \N__35862\
        );

    \I__7415\ : Odrv4
    port map (
            O => \N__35862\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__7414\ : InMux
    port map (
            O => \N__35859\,
            I => \bfn_14_22_0_\
        );

    \I__7413\ : CascadeMux
    port map (
            O => \N__35856\,
            I => \N__35853\
        );

    \I__7412\ : InMux
    port map (
            O => \N__35853\,
            I => \N__35850\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__35850\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__7410\ : InMux
    port map (
            O => \N__35847\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__7409\ : InMux
    port map (
            O => \N__35844\,
            I => \N__35841\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__35841\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__7407\ : InMux
    port map (
            O => \N__35838\,
            I => \N__35834\
        );

    \I__7406\ : InMux
    port map (
            O => \N__35837\,
            I => \N__35831\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__35834\,
            I => \N__35826\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__35831\,
            I => \N__35826\
        );

    \I__7403\ : Odrv4
    port map (
            O => \N__35826\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__7402\ : InMux
    port map (
            O => \N__35823\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__7401\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35814\
        );

    \I__7400\ : InMux
    port map (
            O => \N__35819\,
            I => \N__35809\
        );

    \I__7399\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35809\
        );

    \I__7398\ : InMux
    port map (
            O => \N__35817\,
            I => \N__35806\
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__35814\,
            I => \N__35803\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__35809\,
            I => \N__35798\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__35806\,
            I => \N__35798\
        );

    \I__7394\ : Odrv4
    port map (
            O => \N__35803\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__7393\ : Odrv4
    port map (
            O => \N__35798\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__7392\ : InMux
    port map (
            O => \N__35793\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__7391\ : InMux
    port map (
            O => \N__35790\,
            I => \N__35786\
        );

    \I__7390\ : InMux
    port map (
            O => \N__35789\,
            I => \N__35783\
        );

    \I__7389\ : LocalMux
    port map (
            O => \N__35786\,
            I => \N__35780\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__35783\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__7387\ : Odrv12
    port map (
            O => \N__35780\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__7386\ : InMux
    port map (
            O => \N__35775\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__7385\ : CascadeMux
    port map (
            O => \N__35772\,
            I => \N__35769\
        );

    \I__7384\ : InMux
    port map (
            O => \N__35769\,
            I => \N__35765\
        );

    \I__7383\ : InMux
    port map (
            O => \N__35768\,
            I => \N__35762\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__35765\,
            I => \N__35759\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__35762\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__7380\ : Odrv4
    port map (
            O => \N__35759\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__7379\ : InMux
    port map (
            O => \N__35754\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__7378\ : CascadeMux
    port map (
            O => \N__35751\,
            I => \N__35746\
        );

    \I__7377\ : InMux
    port map (
            O => \N__35750\,
            I => \N__35742\
        );

    \I__7376\ : CascadeMux
    port map (
            O => \N__35749\,
            I => \N__35738\
        );

    \I__7375\ : InMux
    port map (
            O => \N__35746\,
            I => \N__35735\
        );

    \I__7374\ : InMux
    port map (
            O => \N__35745\,
            I => \N__35732\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__35742\,
            I => \N__35729\
        );

    \I__7372\ : InMux
    port map (
            O => \N__35741\,
            I => \N__35726\
        );

    \I__7371\ : InMux
    port map (
            O => \N__35738\,
            I => \N__35723\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__35735\,
            I => \N__35718\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__35732\,
            I => \N__35718\
        );

    \I__7368\ : Span4Mux_h
    port map (
            O => \N__35729\,
            I => \N__35713\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__35726\,
            I => \N__35713\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__35723\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__7365\ : Odrv4
    port map (
            O => \N__35718\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__7364\ : Odrv4
    port map (
            O => \N__35713\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__7363\ : InMux
    port map (
            O => \N__35706\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__7362\ : InMux
    port map (
            O => \N__35703\,
            I => \N__35699\
        );

    \I__7361\ : InMux
    port map (
            O => \N__35702\,
            I => \N__35696\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__35699\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__35696\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__7358\ : InMux
    port map (
            O => \N__35691\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__7357\ : InMux
    port map (
            O => \N__35688\,
            I => \N__35684\
        );

    \I__7356\ : InMux
    port map (
            O => \N__35687\,
            I => \N__35681\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__35684\,
            I => \N__35678\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__35681\,
            I => \N__35675\
        );

    \I__7353\ : Odrv4
    port map (
            O => \N__35678\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__7352\ : Odrv4
    port map (
            O => \N__35675\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__7351\ : InMux
    port map (
            O => \N__35670\,
            I => \bfn_14_21_0_\
        );

    \I__7350\ : InMux
    port map (
            O => \N__35667\,
            I => \N__35664\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__35664\,
            I => \N__35660\
        );

    \I__7348\ : InMux
    port map (
            O => \N__35663\,
            I => \N__35657\
        );

    \I__7347\ : Span4Mux_h
    port map (
            O => \N__35660\,
            I => \N__35654\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__35657\,
            I => \N__35651\
        );

    \I__7345\ : Odrv4
    port map (
            O => \N__35654\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__7344\ : Odrv4
    port map (
            O => \N__35651\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__7343\ : InMux
    port map (
            O => \N__35646\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__7342\ : CascadeMux
    port map (
            O => \N__35643\,
            I => \delay_measurement_inst.N_333_cascade_\
        );

    \I__7341\ : InMux
    port map (
            O => \N__35640\,
            I => \N__35636\
        );

    \I__7340\ : InMux
    port map (
            O => \N__35639\,
            I => \N__35633\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__35636\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__35633\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__7337\ : InMux
    port map (
            O => \N__35628\,
            I => \N__35623\
        );

    \I__7336\ : InMux
    port map (
            O => \N__35627\,
            I => \N__35620\
        );

    \I__7335\ : InMux
    port map (
            O => \N__35626\,
            I => \N__35617\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__35623\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__35620\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__35617\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__7331\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35595\
        );

    \I__7330\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35595\
        );

    \I__7329\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35595\
        );

    \I__7328\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35595\
        );

    \I__7327\ : InMux
    port map (
            O => \N__35606\,
            I => \N__35595\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__35595\,
            I => \delay_measurement_inst.N_333\
        );

    \I__7325\ : InMux
    port map (
            O => \N__35592\,
            I => \N__35588\
        );

    \I__7324\ : InMux
    port map (
            O => \N__35591\,
            I => \N__35585\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__35588\,
            I => \N__35580\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__35585\,
            I => \N__35580\
        );

    \I__7321\ : Span4Mux_v
    port map (
            O => \N__35580\,
            I => \N__35577\
        );

    \I__7320\ : Span4Mux_h
    port map (
            O => \N__35577\,
            I => \N__35573\
        );

    \I__7319\ : InMux
    port map (
            O => \N__35576\,
            I => \N__35570\
        );

    \I__7318\ : Odrv4
    port map (
            O => \N__35573\,
            I => \delay_measurement_inst.N_328\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__35570\,
            I => \delay_measurement_inst.N_328\
        );

    \I__7316\ : CascadeMux
    port map (
            O => \N__35565\,
            I => \N__35558\
        );

    \I__7315\ : CascadeMux
    port map (
            O => \N__35564\,
            I => \N__35554\
        );

    \I__7314\ : CascadeMux
    port map (
            O => \N__35563\,
            I => \N__35551\
        );

    \I__7313\ : InMux
    port map (
            O => \N__35562\,
            I => \N__35544\
        );

    \I__7312\ : InMux
    port map (
            O => \N__35561\,
            I => \N__35544\
        );

    \I__7311\ : InMux
    port map (
            O => \N__35558\,
            I => \N__35541\
        );

    \I__7310\ : InMux
    port map (
            O => \N__35557\,
            I => \N__35530\
        );

    \I__7309\ : InMux
    port map (
            O => \N__35554\,
            I => \N__35530\
        );

    \I__7308\ : InMux
    port map (
            O => \N__35551\,
            I => \N__35530\
        );

    \I__7307\ : InMux
    port map (
            O => \N__35550\,
            I => \N__35530\
        );

    \I__7306\ : InMux
    port map (
            O => \N__35549\,
            I => \N__35530\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__35544\,
            I => \N__35527\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__35541\,
            I => \N__35522\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__35530\,
            I => \N__35522\
        );

    \I__7302\ : Span4Mux_h
    port map (
            O => \N__35527\,
            I => \N__35519\
        );

    \I__7301\ : Span4Mux_v
    port map (
            O => \N__35522\,
            I => \N__35516\
        );

    \I__7300\ : Odrv4
    port map (
            O => \N__35519\,
            I => \delay_measurement_inst.N_324\
        );

    \I__7299\ : Odrv4
    port map (
            O => \N__35516\,
            I => \delay_measurement_inst.N_324\
        );

    \I__7298\ : CEMux
    port map (
            O => \N__35511\,
            I => \N__35504\
        );

    \I__7297\ : CEMux
    port map (
            O => \N__35510\,
            I => \N__35501\
        );

    \I__7296\ : CEMux
    port map (
            O => \N__35509\,
            I => \N__35498\
        );

    \I__7295\ : CEMux
    port map (
            O => \N__35508\,
            I => \N__35495\
        );

    \I__7294\ : CEMux
    port map (
            O => \N__35507\,
            I => \N__35492\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__35504\,
            I => \N__35489\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__35501\,
            I => \N__35486\
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__35498\,
            I => \N__35483\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__35495\,
            I => \N__35480\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__35492\,
            I => \N__35477\
        );

    \I__7288\ : Span4Mux_v
    port map (
            O => \N__35489\,
            I => \N__35472\
        );

    \I__7287\ : Span4Mux_h
    port map (
            O => \N__35486\,
            I => \N__35472\
        );

    \I__7286\ : Span4Mux_v
    port map (
            O => \N__35483\,
            I => \N__35467\
        );

    \I__7285\ : Span4Mux_h
    port map (
            O => \N__35480\,
            I => \N__35467\
        );

    \I__7284\ : Odrv12
    port map (
            O => \N__35477\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__7283\ : Odrv4
    port map (
            O => \N__35472\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__7282\ : Odrv4
    port map (
            O => \N__35467\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__7281\ : CascadeMux
    port map (
            O => \N__35460\,
            I => \N__35456\
        );

    \I__7280\ : CascadeMux
    port map (
            O => \N__35459\,
            I => \N__35453\
        );

    \I__7279\ : InMux
    port map (
            O => \N__35456\,
            I => \N__35449\
        );

    \I__7278\ : InMux
    port map (
            O => \N__35453\,
            I => \N__35444\
        );

    \I__7277\ : InMux
    port map (
            O => \N__35452\,
            I => \N__35444\
        );

    \I__7276\ : LocalMux
    port map (
            O => \N__35449\,
            I => \N__35439\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__35444\,
            I => \N__35439\
        );

    \I__7274\ : Odrv4
    port map (
            O => \N__35439\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__7273\ : InMux
    port map (
            O => \N__35436\,
            I => \N__35432\
        );

    \I__7272\ : InMux
    port map (
            O => \N__35435\,
            I => \N__35429\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__35432\,
            I => \N__35426\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__35429\,
            I => \N__35423\
        );

    \I__7269\ : Odrv12
    port map (
            O => \N__35426\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__7268\ : Odrv4
    port map (
            O => \N__35423\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__7267\ : InMux
    port map (
            O => \N__35418\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__7266\ : CascadeMux
    port map (
            O => \N__35415\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_\
        );

    \I__7265\ : CascadeMux
    port map (
            O => \N__35412\,
            I => \N__35407\
        );

    \I__7264\ : InMux
    port map (
            O => \N__35411\,
            I => \N__35403\
        );

    \I__7263\ : InMux
    port map (
            O => \N__35410\,
            I => \N__35400\
        );

    \I__7262\ : InMux
    port map (
            O => \N__35407\,
            I => \N__35395\
        );

    \I__7261\ : InMux
    port map (
            O => \N__35406\,
            I => \N__35395\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__35403\,
            I => \N__35392\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__35400\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__35395\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__7257\ : Odrv4
    port map (
            O => \N__35392\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__7256\ : InMux
    port map (
            O => \N__35385\,
            I => \N__35380\
        );

    \I__7255\ : InMux
    port map (
            O => \N__35384\,
            I => \N__35377\
        );

    \I__7254\ : InMux
    port map (
            O => \N__35383\,
            I => \N__35374\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__35380\,
            I => \N__35371\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__35377\,
            I => \N__35366\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__35374\,
            I => \N__35366\
        );

    \I__7250\ : Span4Mux_h
    port map (
            O => \N__35371\,
            I => \N__35361\
        );

    \I__7249\ : Span4Mux_v
    port map (
            O => \N__35366\,
            I => \N__35361\
        );

    \I__7248\ : Span4Mux_h
    port map (
            O => \N__35361\,
            I => \N__35358\
        );

    \I__7247\ : Sp12to4
    port map (
            O => \N__35358\,
            I => \N__35355\
        );

    \I__7246\ : Odrv12
    port map (
            O => \N__35355\,
            I => \il_min_comp2_D2\
        );

    \I__7245\ : InMux
    port map (
            O => \N__35352\,
            I => \N__35349\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__35349\,
            I => \N__35346\
        );

    \I__7243\ : Odrv4
    port map (
            O => \N__35346\,
            I => \phase_controller_slave.start_timer_tr_0_sqmuxa\
        );

    \I__7242\ : InMux
    port map (
            O => \N__35343\,
            I => \N__35340\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__35340\,
            I => \N__35336\
        );

    \I__7240\ : InMux
    port map (
            O => \N__35339\,
            I => \N__35333\
        );

    \I__7239\ : Span4Mux_h
    port map (
            O => \N__35336\,
            I => \N__35329\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__35333\,
            I => \N__35326\
        );

    \I__7237\ : InMux
    port map (
            O => \N__35332\,
            I => \N__35323\
        );

    \I__7236\ : Span4Mux_v
    port map (
            O => \N__35329\,
            I => \N__35320\
        );

    \I__7235\ : Odrv4
    port map (
            O => \N__35326\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__35323\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7233\ : Odrv4
    port map (
            O => \N__35320\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7232\ : InMux
    port map (
            O => \N__35313\,
            I => \N__35309\
        );

    \I__7231\ : InMux
    port map (
            O => \N__35312\,
            I => \N__35306\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__35309\,
            I => \N__35303\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__35306\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7228\ : Odrv12
    port map (
            O => \N__35303\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7227\ : CascadeMux
    port map (
            O => \N__35298\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6_cascade_\
        );

    \I__7226\ : CascadeMux
    port map (
            O => \N__35295\,
            I => \N__35291\
        );

    \I__7225\ : InMux
    port map (
            O => \N__35294\,
            I => \N__35282\
        );

    \I__7224\ : InMux
    port map (
            O => \N__35291\,
            I => \N__35279\
        );

    \I__7223\ : InMux
    port map (
            O => \N__35290\,
            I => \N__35276\
        );

    \I__7222\ : InMux
    port map (
            O => \N__35289\,
            I => \N__35273\
        );

    \I__7221\ : InMux
    port map (
            O => \N__35288\,
            I => \N__35270\
        );

    \I__7220\ : InMux
    port map (
            O => \N__35287\,
            I => \N__35265\
        );

    \I__7219\ : InMux
    port map (
            O => \N__35286\,
            I => \N__35265\
        );

    \I__7218\ : InMux
    port map (
            O => \N__35285\,
            I => \N__35262\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__35282\,
            I => \N__35259\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__35279\,
            I => \N__35256\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__35276\,
            I => \N__35251\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__35273\,
            I => \N__35251\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__35270\,
            I => \delay_measurement_inst.N_358\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__35265\,
            I => \delay_measurement_inst.N_358\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__35262\,
            I => \delay_measurement_inst.N_358\
        );

    \I__7210\ : Odrv4
    port map (
            O => \N__35259\,
            I => \delay_measurement_inst.N_358\
        );

    \I__7209\ : Odrv12
    port map (
            O => \N__35256\,
            I => \delay_measurement_inst.N_358\
        );

    \I__7208\ : Odrv4
    port map (
            O => \N__35251\,
            I => \delay_measurement_inst.N_358\
        );

    \I__7207\ : InMux
    port map (
            O => \N__35238\,
            I => \N__35232\
        );

    \I__7206\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35232\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__35232\,
            I => \delay_measurement_inst.delay_tr_timer.N_331\
        );

    \I__7204\ : CascadeMux
    port map (
            O => \N__35229\,
            I => \delay_measurement_inst.delay_tr_timer.N_331_cascade_\
        );

    \I__7203\ : CascadeMux
    port map (
            O => \N__35226\,
            I => \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa_cascade_\
        );

    \I__7202\ : CascadeMux
    port map (
            O => \N__35223\,
            I => \N__35219\
        );

    \I__7201\ : InMux
    port map (
            O => \N__35222\,
            I => \N__35211\
        );

    \I__7200\ : InMux
    port map (
            O => \N__35219\,
            I => \N__35211\
        );

    \I__7199\ : InMux
    port map (
            O => \N__35218\,
            I => \N__35211\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__35211\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__7197\ : InMux
    port map (
            O => \N__35208\,
            I => \N__35202\
        );

    \I__7196\ : InMux
    port map (
            O => \N__35207\,
            I => \N__35202\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__35202\,
            I => \phase_controller_slave.stateZ0Z_0\
        );

    \I__7194\ : InMux
    port map (
            O => \N__35199\,
            I => \N__35194\
        );

    \I__7193\ : InMux
    port map (
            O => \N__35198\,
            I => \N__35189\
        );

    \I__7192\ : InMux
    port map (
            O => \N__35197\,
            I => \N__35189\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__35194\,
            I => \N__35186\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__35189\,
            I => \N__35183\
        );

    \I__7189\ : Span4Mux_v
    port map (
            O => \N__35186\,
            I => \N__35178\
        );

    \I__7188\ : Span4Mux_v
    port map (
            O => \N__35183\,
            I => \N__35178\
        );

    \I__7187\ : Span4Mux_v
    port map (
            O => \N__35178\,
            I => \N__35175\
        );

    \I__7186\ : Odrv4
    port map (
            O => \N__35175\,
            I => \il_max_comp2_D2\
        );

    \I__7185\ : InMux
    port map (
            O => \N__35172\,
            I => \N__35169\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__35169\,
            I => \phase_controller_slave.N_211\
        );

    \I__7183\ : CascadeMux
    port map (
            O => \N__35166\,
            I => \N__35162\
        );

    \I__7182\ : CascadeMux
    port map (
            O => \N__35165\,
            I => \N__35158\
        );

    \I__7181\ : InMux
    port map (
            O => \N__35162\,
            I => \N__35151\
        );

    \I__7180\ : InMux
    port map (
            O => \N__35161\,
            I => \N__35151\
        );

    \I__7179\ : InMux
    port map (
            O => \N__35158\,
            I => \N__35148\
        );

    \I__7178\ : InMux
    port map (
            O => \N__35157\,
            I => \N__35143\
        );

    \I__7177\ : InMux
    port map (
            O => \N__35156\,
            I => \N__35143\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__35151\,
            I => \N__35140\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__35148\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__35143\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__7173\ : Odrv4
    port map (
            O => \N__35140\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__7172\ : InMux
    port map (
            O => \N__35133\,
            I => \N__35129\
        );

    \I__7171\ : InMux
    port map (
            O => \N__35132\,
            I => \N__35126\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__35129\,
            I => \N__35123\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__35126\,
            I => \N__35120\
        );

    \I__7168\ : Span4Mux_v
    port map (
            O => \N__35123\,
            I => \N__35114\
        );

    \I__7167\ : Span4Mux_h
    port map (
            O => \N__35120\,
            I => \N__35114\
        );

    \I__7166\ : InMux
    port map (
            O => \N__35119\,
            I => \N__35111\
        );

    \I__7165\ : Odrv4
    port map (
            O => \N__35114\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__35111\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__7163\ : InMux
    port map (
            O => \N__35106\,
            I => \N__35103\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__35103\,
            I => \N__35098\
        );

    \I__7161\ : InMux
    port map (
            O => \N__35102\,
            I => \N__35095\
        );

    \I__7160\ : InMux
    port map (
            O => \N__35101\,
            I => \N__35092\
        );

    \I__7159\ : Span4Mux_v
    port map (
            O => \N__35098\,
            I => \N__35089\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__35095\,
            I => \N__35084\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__35092\,
            I => \N__35084\
        );

    \I__7156\ : Span4Mux_h
    port map (
            O => \N__35089\,
            I => \N__35081\
        );

    \I__7155\ : Span4Mux_v
    port map (
            O => \N__35084\,
            I => \N__35078\
        );

    \I__7154\ : Odrv4
    port map (
            O => \N__35081\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__7153\ : Odrv4
    port map (
            O => \N__35078\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__7152\ : InMux
    port map (
            O => \N__35073\,
            I => \N__35069\
        );

    \I__7151\ : InMux
    port map (
            O => \N__35072\,
            I => \N__35066\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__35069\,
            I => \N__35060\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__35066\,
            I => \N__35060\
        );

    \I__7148\ : InMux
    port map (
            O => \N__35065\,
            I => \N__35056\
        );

    \I__7147\ : Span4Mux_s3_v
    port map (
            O => \N__35060\,
            I => \N__35051\
        );

    \I__7146\ : CascadeMux
    port map (
            O => \N__35059\,
            I => \N__35048\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__35056\,
            I => \N__35044\
        );

    \I__7144\ : InMux
    port map (
            O => \N__35055\,
            I => \N__35041\
        );

    \I__7143\ : InMux
    port map (
            O => \N__35054\,
            I => \N__35038\
        );

    \I__7142\ : Span4Mux_h
    port map (
            O => \N__35051\,
            I => \N__35034\
        );

    \I__7141\ : InMux
    port map (
            O => \N__35048\,
            I => \N__35031\
        );

    \I__7140\ : InMux
    port map (
            O => \N__35047\,
            I => \N__35028\
        );

    \I__7139\ : Span4Mux_v
    port map (
            O => \N__35044\,
            I => \N__35023\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__35041\,
            I => \N__35023\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__35038\,
            I => \N__35020\
        );

    \I__7136\ : InMux
    port map (
            O => \N__35037\,
            I => \N__35017\
        );

    \I__7135\ : Sp12to4
    port map (
            O => \N__35034\,
            I => \N__35014\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__35031\,
            I => \N__35009\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__35028\,
            I => \N__35009\
        );

    \I__7132\ : Span4Mux_v
    port map (
            O => \N__35023\,
            I => \N__35002\
        );

    \I__7131\ : Span4Mux_v
    port map (
            O => \N__35020\,
            I => \N__35002\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__35017\,
            I => \N__35002\
        );

    \I__7129\ : Span12Mux_v
    port map (
            O => \N__35014\,
            I => \N__34999\
        );

    \I__7128\ : Span4Mux_v
    port map (
            O => \N__35009\,
            I => \N__34996\
        );

    \I__7127\ : Span4Mux_v
    port map (
            O => \N__35002\,
            I => \N__34993\
        );

    \I__7126\ : Span12Mux_v
    port map (
            O => \N__34999\,
            I => \N__34988\
        );

    \I__7125\ : Sp12to4
    port map (
            O => \N__34996\,
            I => \N__34988\
        );

    \I__7124\ : Span4Mux_h
    port map (
            O => \N__34993\,
            I => \N__34985\
        );

    \I__7123\ : Span12Mux_h
    port map (
            O => \N__34988\,
            I => \N__34982\
        );

    \I__7122\ : Span4Mux_v
    port map (
            O => \N__34985\,
            I => \N__34979\
        );

    \I__7121\ : Odrv12
    port map (
            O => \N__34982\,
            I => start_stop_c
        );

    \I__7120\ : Odrv4
    port map (
            O => \N__34979\,
            I => start_stop_c
        );

    \I__7119\ : InMux
    port map (
            O => \N__34974\,
            I => \N__34964\
        );

    \I__7118\ : InMux
    port map (
            O => \N__34973\,
            I => \N__34964\
        );

    \I__7117\ : InMux
    port map (
            O => \N__34972\,
            I => \N__34964\
        );

    \I__7116\ : InMux
    port map (
            O => \N__34971\,
            I => \N__34961\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__34964\,
            I => \N__34958\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__34961\,
            I => \N__34955\
        );

    \I__7113\ : Span4Mux_v
    port map (
            O => \N__34958\,
            I => \N__34952\
        );

    \I__7112\ : Span4Mux_h
    port map (
            O => \N__34955\,
            I => \N__34949\
        );

    \I__7111\ : Odrv4
    port map (
            O => \N__34952\,
            I => shift_flag_start
        );

    \I__7110\ : Odrv4
    port map (
            O => \N__34949\,
            I => shift_flag_start
        );

    \I__7109\ : InMux
    port map (
            O => \N__34944\,
            I => \N__34938\
        );

    \I__7108\ : InMux
    port map (
            O => \N__34943\,
            I => \N__34935\
        );

    \I__7107\ : InMux
    port map (
            O => \N__34942\,
            I => \N__34930\
        );

    \I__7106\ : InMux
    port map (
            O => \N__34941\,
            I => \N__34930\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__34938\,
            I => \N__34927\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__34935\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__34930\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__7102\ : Odrv4
    port map (
            O => \N__34927\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__7101\ : InMux
    port map (
            O => \N__34920\,
            I => \N__34917\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__34917\,
            I => \phase_controller_slave.N_213\
        );

    \I__7099\ : InMux
    port map (
            O => \N__34914\,
            I => \N__34911\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__34911\,
            I => \phase_controller_slave.start_timer_hc_0_sqmuxa\
        );

    \I__7097\ : InMux
    port map (
            O => \N__34908\,
            I => \N__34905\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__34905\,
            I => \phase_controller_slave.N_214\
        );

    \I__7095\ : IoInMux
    port map (
            O => \N__34902\,
            I => \N__34899\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__34899\,
            I => \N__34896\
        );

    \I__7093\ : Span12Mux_s4_v
    port map (
            O => \N__34896\,
            I => \N__34892\
        );

    \I__7092\ : CascadeMux
    port map (
            O => \N__34895\,
            I => \N__34889\
        );

    \I__7091\ : Span12Mux_v
    port map (
            O => \N__34892\,
            I => \N__34886\
        );

    \I__7090\ : InMux
    port map (
            O => \N__34889\,
            I => \N__34883\
        );

    \I__7089\ : Odrv12
    port map (
            O => \N__34886\,
            I => s4_phy_c
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__34883\,
            I => s4_phy_c
        );

    \I__7087\ : InMux
    port map (
            O => \N__34878\,
            I => \N__34873\
        );

    \I__7086\ : InMux
    port map (
            O => \N__34877\,
            I => \N__34870\
        );

    \I__7085\ : InMux
    port map (
            O => \N__34876\,
            I => \N__34867\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__34873\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__34870\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__34867\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__7081\ : InMux
    port map (
            O => \N__34860\,
            I => \N__34854\
        );

    \I__7080\ : InMux
    port map (
            O => \N__34859\,
            I => \N__34851\
        );

    \I__7079\ : InMux
    port map (
            O => \N__34858\,
            I => \N__34848\
        );

    \I__7078\ : InMux
    port map (
            O => \N__34857\,
            I => \N__34845\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__34854\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__34851\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__34848\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__34845\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__7073\ : IoInMux
    port map (
            O => \N__34836\,
            I => \N__34833\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__34833\,
            I => \N__34830\
        );

    \I__7071\ : Span4Mux_s0_v
    port map (
            O => \N__34830\,
            I => \N__34827\
        );

    \I__7070\ : Sp12to4
    port map (
            O => \N__34827\,
            I => \N__34824\
        );

    \I__7069\ : Span12Mux_h
    port map (
            O => \N__34824\,
            I => \N__34820\
        );

    \I__7068\ : CascadeMux
    port map (
            O => \N__34823\,
            I => \N__34816\
        );

    \I__7067\ : Span12Mux_v
    port map (
            O => \N__34820\,
            I => \N__34813\
        );

    \I__7066\ : InMux
    port map (
            O => \N__34819\,
            I => \N__34810\
        );

    \I__7065\ : InMux
    port map (
            O => \N__34816\,
            I => \N__34807\
        );

    \I__7064\ : Odrv12
    port map (
            O => \N__34813\,
            I => s3_phy_c
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__34810\,
            I => s3_phy_c
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__34807\,
            I => s3_phy_c
        );

    \I__7061\ : CascadeMux
    port map (
            O => \N__34800\,
            I => \phase_controller_slave.N_211_cascade_\
        );

    \I__7060\ : IoInMux
    port map (
            O => \N__34797\,
            I => \N__34794\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__34794\,
            I => \N__34790\
        );

    \I__7058\ : CEMux
    port map (
            O => \N__34793\,
            I => \N__34787\
        );

    \I__7057\ : IoSpan4Mux
    port map (
            O => \N__34790\,
            I => \N__34782\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__34787\,
            I => \N__34778\
        );

    \I__7055\ : CEMux
    port map (
            O => \N__34786\,
            I => \N__34775\
        );

    \I__7054\ : CEMux
    port map (
            O => \N__34785\,
            I => \N__34772\
        );

    \I__7053\ : Span4Mux_s3_v
    port map (
            O => \N__34782\,
            I => \N__34769\
        );

    \I__7052\ : CEMux
    port map (
            O => \N__34781\,
            I => \N__34766\
        );

    \I__7051\ : Span4Mux_v
    port map (
            O => \N__34778\,
            I => \N__34761\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__34775\,
            I => \N__34761\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__34772\,
            I => \N__34758\
        );

    \I__7048\ : Sp12to4
    port map (
            O => \N__34769\,
            I => \N__34755\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__34766\,
            I => \N__34752\
        );

    \I__7046\ : Span4Mux_v
    port map (
            O => \N__34761\,
            I => \N__34747\
        );

    \I__7045\ : Span4Mux_h
    port map (
            O => \N__34758\,
            I => \N__34747\
        );

    \I__7044\ : Span12Mux_s11_v
    port map (
            O => \N__34755\,
            I => \N__34742\
        );

    \I__7043\ : Sp12to4
    port map (
            O => \N__34752\,
            I => \N__34742\
        );

    \I__7042\ : Span4Mux_v
    port map (
            O => \N__34747\,
            I => \N__34739\
        );

    \I__7041\ : Odrv12
    port map (
            O => \N__34742\,
            I => red_c_i
        );

    \I__7040\ : Odrv4
    port map (
            O => \N__34739\,
            I => red_c_i
        );

    \I__7039\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34731\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__34731\,
            I => \N__34726\
        );

    \I__7037\ : CascadeMux
    port map (
            O => \N__34730\,
            I => \N__34722\
        );

    \I__7036\ : InMux
    port map (
            O => \N__34729\,
            I => \N__34719\
        );

    \I__7035\ : Sp12to4
    port map (
            O => \N__34726\,
            I => \N__34715\
        );

    \I__7034\ : CascadeMux
    port map (
            O => \N__34725\,
            I => \N__34712\
        );

    \I__7033\ : InMux
    port map (
            O => \N__34722\,
            I => \N__34709\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__34719\,
            I => \N__34706\
        );

    \I__7031\ : InMux
    port map (
            O => \N__34718\,
            I => \N__34703\
        );

    \I__7030\ : Span12Mux_v
    port map (
            O => \N__34715\,
            I => \N__34700\
        );

    \I__7029\ : InMux
    port map (
            O => \N__34712\,
            I => \N__34697\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__34709\,
            I => \N__34690\
        );

    \I__7027\ : Span4Mux_v
    port map (
            O => \N__34706\,
            I => \N__34690\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__34703\,
            I => \N__34690\
        );

    \I__7025\ : Odrv12
    port map (
            O => \N__34700\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__34697\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7023\ : Odrv4
    port map (
            O => \N__34690\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__7022\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34678\
        );

    \I__7021\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34675\
        );

    \I__7020\ : InMux
    port map (
            O => \N__34681\,
            I => \N__34672\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__34678\,
            I => \N__34667\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__34675\,
            I => \N__34667\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__34672\,
            I => \N__34664\
        );

    \I__7016\ : Span4Mux_v
    port map (
            O => \N__34667\,
            I => \N__34661\
        );

    \I__7015\ : Odrv12
    port map (
            O => \N__34664\,
            I => \il_min_comp1_D2\
        );

    \I__7014\ : Odrv4
    port map (
            O => \N__34661\,
            I => \il_min_comp1_D2\
        );

    \I__7013\ : InMux
    port map (
            O => \N__34656\,
            I => \N__34653\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__34653\,
            I => \phase_controller_inst1.N_232\
        );

    \I__7011\ : CascadeMux
    port map (
            O => \N__34650\,
            I => \N__34647\
        );

    \I__7010\ : InMux
    port map (
            O => \N__34647\,
            I => \N__34644\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__34644\,
            I => \N__34641\
        );

    \I__7008\ : Odrv4
    port map (
            O => \N__34641\,
            I => \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__7007\ : InMux
    port map (
            O => \N__34638\,
            I => \N__34635\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__34635\,
            I => \N__34631\
        );

    \I__7005\ : InMux
    port map (
            O => \N__34634\,
            I => \N__34628\
        );

    \I__7004\ : Span4Mux_v
    port map (
            O => \N__34631\,
            I => \N__34623\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__34628\,
            I => \N__34620\
        );

    \I__7002\ : InMux
    port map (
            O => \N__34627\,
            I => \N__34617\
        );

    \I__7001\ : InMux
    port map (
            O => \N__34626\,
            I => \N__34614\
        );

    \I__7000\ : Odrv4
    port map (
            O => \N__34623\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__6999\ : Odrv4
    port map (
            O => \N__34620\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__34617\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__34614\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__6996\ : CascadeMux
    port map (
            O => \N__34605\,
            I => \N__34602\
        );

    \I__6995\ : InMux
    port map (
            O => \N__34602\,
            I => \N__34599\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__34599\,
            I => \N__34596\
        );

    \I__6993\ : Span4Mux_h
    port map (
            O => \N__34596\,
            I => \N__34593\
        );

    \I__6992\ : Odrv4
    port map (
            O => \N__34593\,
            I => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__6991\ : InMux
    port map (
            O => \N__34590\,
            I => \N__34586\
        );

    \I__6990\ : InMux
    port map (
            O => \N__34589\,
            I => \N__34583\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__34586\,
            I => \N__34576\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__34583\,
            I => \N__34573\
        );

    \I__6987\ : InMux
    port map (
            O => \N__34582\,
            I => \N__34570\
        );

    \I__6986\ : InMux
    port map (
            O => \N__34581\,
            I => \N__34563\
        );

    \I__6985\ : InMux
    port map (
            O => \N__34580\,
            I => \N__34563\
        );

    \I__6984\ : InMux
    port map (
            O => \N__34579\,
            I => \N__34563\
        );

    \I__6983\ : Odrv4
    port map (
            O => \N__34576\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6982\ : Odrv4
    port map (
            O => \N__34573\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__34570\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__34563\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6979\ : InMux
    port map (
            O => \N__34554\,
            I => \N__34550\
        );

    \I__6978\ : InMux
    port map (
            O => \N__34553\,
            I => \N__34547\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__34550\,
            I => \N__34541\
        );

    \I__6976\ : LocalMux
    port map (
            O => \N__34547\,
            I => \N__34541\
        );

    \I__6975\ : InMux
    port map (
            O => \N__34546\,
            I => \N__34538\
        );

    \I__6974\ : Span4Mux_v
    port map (
            O => \N__34541\,
            I => \N__34533\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__34538\,
            I => \N__34533\
        );

    \I__6972\ : Span4Mux_v
    port map (
            O => \N__34533\,
            I => \N__34530\
        );

    \I__6971\ : Odrv4
    port map (
            O => \N__34530\,
            I => \il_max_comp1_D2\
        );

    \I__6970\ : InMux
    port map (
            O => \N__34527\,
            I => \N__34523\
        );

    \I__6969\ : CascadeMux
    port map (
            O => \N__34526\,
            I => \N__34518\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__34523\,
            I => \N__34515\
        );

    \I__6967\ : CascadeMux
    port map (
            O => \N__34522\,
            I => \N__34511\
        );

    \I__6966\ : CascadeMux
    port map (
            O => \N__34521\,
            I => \N__34508\
        );

    \I__6965\ : InMux
    port map (
            O => \N__34518\,
            I => \N__34505\
        );

    \I__6964\ : Span4Mux_v
    port map (
            O => \N__34515\,
            I => \N__34502\
        );

    \I__6963\ : InMux
    port map (
            O => \N__34514\,
            I => \N__34499\
        );

    \I__6962\ : InMux
    port map (
            O => \N__34511\,
            I => \N__34496\
        );

    \I__6961\ : InMux
    port map (
            O => \N__34508\,
            I => \N__34493\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34490\
        );

    \I__6959\ : Span4Mux_v
    port map (
            O => \N__34502\,
            I => \N__34487\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__34499\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__34496\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__34493\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__6955\ : Odrv12
    port map (
            O => \N__34490\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__6954\ : Odrv4
    port map (
            O => \N__34487\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__6953\ : InMux
    port map (
            O => \N__34476\,
            I => \N__34466\
        );

    \I__6952\ : InMux
    port map (
            O => \N__34475\,
            I => \N__34466\
        );

    \I__6951\ : InMux
    port map (
            O => \N__34474\,
            I => \N__34466\
        );

    \I__6950\ : InMux
    port map (
            O => \N__34473\,
            I => \N__34463\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__34466\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__34463\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6947\ : InMux
    port map (
            O => \N__34458\,
            I => \N__34455\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__34455\,
            I => \N__34452\
        );

    \I__6945\ : Span4Mux_v
    port map (
            O => \N__34452\,
            I => \N__34446\
        );

    \I__6944\ : InMux
    port map (
            O => \N__34451\,
            I => \N__34441\
        );

    \I__6943\ : InMux
    port map (
            O => \N__34450\,
            I => \N__34441\
        );

    \I__6942\ : InMux
    port map (
            O => \N__34449\,
            I => \N__34438\
        );

    \I__6941\ : Odrv4
    port map (
            O => \N__34446\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__34441\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__34438\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6938\ : CascadeMux
    port map (
            O => \N__34431\,
            I => \N__34427\
        );

    \I__6937\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34423\
        );

    \I__6936\ : InMux
    port map (
            O => \N__34427\,
            I => \N__34419\
        );

    \I__6935\ : CascadeMux
    port map (
            O => \N__34426\,
            I => \N__34416\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__34423\,
            I => \N__34412\
        );

    \I__6933\ : InMux
    port map (
            O => \N__34422\,
            I => \N__34409\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__34419\,
            I => \N__34406\
        );

    \I__6931\ : InMux
    port map (
            O => \N__34416\,
            I => \N__34403\
        );

    \I__6930\ : InMux
    port map (
            O => \N__34415\,
            I => \N__34400\
        );

    \I__6929\ : Span4Mux_h
    port map (
            O => \N__34412\,
            I => \N__34395\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__34409\,
            I => \N__34395\
        );

    \I__6927\ : Span4Mux_v
    port map (
            O => \N__34406\,
            I => \N__34392\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__34403\,
            I => measured_delay_hc_18
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__34400\,
            I => measured_delay_hc_18
        );

    \I__6924\ : Odrv4
    port map (
            O => \N__34395\,
            I => measured_delay_hc_18
        );

    \I__6923\ : Odrv4
    port map (
            O => \N__34392\,
            I => measured_delay_hc_18
        );

    \I__6922\ : InMux
    port map (
            O => \N__34383\,
            I => \N__34376\
        );

    \I__6921\ : InMux
    port map (
            O => \N__34382\,
            I => \N__34376\
        );

    \I__6920\ : InMux
    port map (
            O => \N__34381\,
            I => \N__34373\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__34376\,
            I => \N__34370\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__34373\,
            I => \N__34365\
        );

    \I__6917\ : Span4Mux_v
    port map (
            O => \N__34370\,
            I => \N__34362\
        );

    \I__6916\ : InMux
    port map (
            O => \N__34369\,
            I => \N__34357\
        );

    \I__6915\ : InMux
    port map (
            O => \N__34368\,
            I => \N__34357\
        );

    \I__6914\ : Span4Mux_v
    port map (
            O => \N__34365\,
            I => \N__34354\
        );

    \I__6913\ : Odrv4
    port map (
            O => \N__34362\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_2\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__34357\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_2\
        );

    \I__6911\ : Odrv4
    port map (
            O => \N__34354\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_2\
        );

    \I__6910\ : InMux
    port map (
            O => \N__34347\,
            I => \N__34343\
        );

    \I__6909\ : InMux
    port map (
            O => \N__34346\,
            I => \N__34340\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__34343\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__34340\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__6906\ : InMux
    port map (
            O => \N__34335\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__6905\ : InMux
    port map (
            O => \N__34332\,
            I => \N__34329\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__34329\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\
        );

    \I__6903\ : CascadeMux
    port map (
            O => \N__34326\,
            I => \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_2_cascade_\
        );

    \I__6902\ : InMux
    port map (
            O => \N__34323\,
            I => \N__34320\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__34320\,
            I => \N__34317\
        );

    \I__6900\ : Span4Mux_h
    port map (
            O => \N__34317\,
            I => \N__34314\
        );

    \I__6899\ : Odrv4
    port map (
            O => \N__34314\,
            I => \phase_controller_inst1.stoper_hc.un1_N_4\
        );

    \I__6898\ : InMux
    port map (
            O => \N__34311\,
            I => \N__34308\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__34308\,
            I => \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_3\
        );

    \I__6896\ : InMux
    port map (
            O => \N__34305\,
            I => \N__34302\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__34302\,
            I => \N__34299\
        );

    \I__6894\ : Span4Mux_h
    port map (
            O => \N__34299\,
            I => \N__34296\
        );

    \I__6893\ : Odrv4
    port map (
            O => \N__34296\,
            I => \phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_1\
        );

    \I__6892\ : InMux
    port map (
            O => \N__34293\,
            I => \N__34288\
        );

    \I__6891\ : InMux
    port map (
            O => \N__34292\,
            I => \N__34284\
        );

    \I__6890\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34281\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__34288\,
            I => \N__34278\
        );

    \I__6888\ : InMux
    port map (
            O => \N__34287\,
            I => \N__34275\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__34284\,
            I => \N__34270\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__34281\,
            I => \N__34270\
        );

    \I__6885\ : Span4Mux_h
    port map (
            O => \N__34278\,
            I => \N__34265\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__34275\,
            I => \N__34265\
        );

    \I__6883\ : Span4Mux_v
    port map (
            O => \N__34270\,
            I => \N__34262\
        );

    \I__6882\ : Span4Mux_v
    port map (
            O => \N__34265\,
            I => \N__34259\
        );

    \I__6881\ : Odrv4
    port map (
            O => \N__34262\,
            I => delay_hc_d2
        );

    \I__6880\ : Odrv4
    port map (
            O => \N__34259\,
            I => delay_hc_d2
        );

    \I__6879\ : InMux
    port map (
            O => \N__34254\,
            I => \N__34250\
        );

    \I__6878\ : InMux
    port map (
            O => \N__34253\,
            I => \N__34247\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__34250\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__34247\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__6875\ : CascadeMux
    port map (
            O => \N__34242\,
            I => \N__34239\
        );

    \I__6874\ : InMux
    port map (
            O => \N__34239\,
            I => \N__34236\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__34236\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\
        );

    \I__6872\ : InMux
    port map (
            O => \N__34233\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__6871\ : InMux
    port map (
            O => \N__34230\,
            I => \N__34226\
        );

    \I__6870\ : InMux
    port map (
            O => \N__34229\,
            I => \N__34223\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__34226\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__34223\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__6867\ : InMux
    port map (
            O => \N__34218\,
            I => \N__34215\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__34215\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\
        );

    \I__6865\ : InMux
    port map (
            O => \N__34212\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__6864\ : InMux
    port map (
            O => \N__34209\,
            I => \N__34205\
        );

    \I__6863\ : InMux
    port map (
            O => \N__34208\,
            I => \N__34202\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__34205\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__34202\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__6860\ : InMux
    port map (
            O => \N__34197\,
            I => \N__34194\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__34194\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\
        );

    \I__6858\ : InMux
    port map (
            O => \N__34191\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__6857\ : InMux
    port map (
            O => \N__34188\,
            I => \N__34184\
        );

    \I__6856\ : InMux
    port map (
            O => \N__34187\,
            I => \N__34181\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__34184\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__34181\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__6853\ : InMux
    port map (
            O => \N__34176\,
            I => \N__34173\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__34173\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\
        );

    \I__6851\ : InMux
    port map (
            O => \N__34170\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__6850\ : InMux
    port map (
            O => \N__34167\,
            I => \N__34163\
        );

    \I__6849\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34160\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__34163\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__34160\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__6846\ : CascadeMux
    port map (
            O => \N__34155\,
            I => \N__34152\
        );

    \I__6845\ : InMux
    port map (
            O => \N__34152\,
            I => \N__34149\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__34149\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\
        );

    \I__6843\ : InMux
    port map (
            O => \N__34146\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__6842\ : InMux
    port map (
            O => \N__34143\,
            I => \N__34139\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34142\,
            I => \N__34136\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__34139\,
            I => \N__34133\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__34136\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__6838\ : Odrv4
    port map (
            O => \N__34133\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__6837\ : CascadeMux
    port map (
            O => \N__34128\,
            I => \N__34125\
        );

    \I__6836\ : InMux
    port map (
            O => \N__34125\,
            I => \N__34122\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__34122\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\
        );

    \I__6834\ : InMux
    port map (
            O => \N__34119\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__6833\ : InMux
    port map (
            O => \N__34116\,
            I => \N__34112\
        );

    \I__6832\ : InMux
    port map (
            O => \N__34115\,
            I => \N__34109\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__34112\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__34109\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__6829\ : InMux
    port map (
            O => \N__34104\,
            I => \N__34101\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__34101\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\
        );

    \I__6827\ : InMux
    port map (
            O => \N__34098\,
            I => \bfn_14_7_0_\
        );

    \I__6826\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34091\
        );

    \I__6825\ : InMux
    port map (
            O => \N__34094\,
            I => \N__34088\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__34091\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__34088\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__6822\ : InMux
    port map (
            O => \N__34083\,
            I => \N__34080\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__34080\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\
        );

    \I__6820\ : InMux
    port map (
            O => \N__34077\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__6819\ : InMux
    port map (
            O => \N__34074\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__6818\ : InMux
    port map (
            O => \N__34071\,
            I => \N__34067\
        );

    \I__6817\ : InMux
    port map (
            O => \N__34070\,
            I => \N__34064\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__34067\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__34064\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__6814\ : InMux
    port map (
            O => \N__34059\,
            I => \N__34056\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__34056\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\
        );

    \I__6812\ : InMux
    port map (
            O => \N__34053\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__6811\ : InMux
    port map (
            O => \N__34050\,
            I => \N__34046\
        );

    \I__6810\ : InMux
    port map (
            O => \N__34049\,
            I => \N__34043\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__34046\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__34043\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__6807\ : InMux
    port map (
            O => \N__34038\,
            I => \N__34035\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__34035\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\
        );

    \I__6805\ : InMux
    port map (
            O => \N__34032\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__6804\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34025\
        );

    \I__6803\ : InMux
    port map (
            O => \N__34028\,
            I => \N__34022\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__34025\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__34022\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__6800\ : CascadeMux
    port map (
            O => \N__34017\,
            I => \N__34014\
        );

    \I__6799\ : InMux
    port map (
            O => \N__34014\,
            I => \N__34011\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__34011\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\
        );

    \I__6797\ : InMux
    port map (
            O => \N__34008\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__6796\ : InMux
    port map (
            O => \N__34005\,
            I => \N__34001\
        );

    \I__6795\ : InMux
    port map (
            O => \N__34004\,
            I => \N__33998\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__34001\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__33998\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__6792\ : InMux
    port map (
            O => \N__33993\,
            I => \N__33990\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__33990\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\
        );

    \I__6790\ : InMux
    port map (
            O => \N__33987\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__6789\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33981\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__33981\,
            I => \N__33977\
        );

    \I__6787\ : InMux
    port map (
            O => \N__33980\,
            I => \N__33974\
        );

    \I__6786\ : Odrv4
    port map (
            O => \N__33977\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__33974\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__6784\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33966\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__33966\,
            I => \N__33963\
        );

    \I__6782\ : Span4Mux_h
    port map (
            O => \N__33963\,
            I => \N__33960\
        );

    \I__6781\ : Odrv4
    port map (
            O => \N__33960\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\
        );

    \I__6780\ : InMux
    port map (
            O => \N__33957\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__6779\ : InMux
    port map (
            O => \N__33954\,
            I => \N__33950\
        );

    \I__6778\ : InMux
    port map (
            O => \N__33953\,
            I => \N__33947\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__33950\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__33947\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__6775\ : InMux
    port map (
            O => \N__33942\,
            I => \N__33939\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__33939\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\
        );

    \I__6773\ : InMux
    port map (
            O => \N__33936\,
            I => \bfn_14_6_0_\
        );

    \I__6772\ : InMux
    port map (
            O => \N__33933\,
            I => \N__33929\
        );

    \I__6771\ : InMux
    port map (
            O => \N__33932\,
            I => \N__33926\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__33929\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__33926\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__6768\ : CascadeMux
    port map (
            O => \N__33921\,
            I => \N__33918\
        );

    \I__6767\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33915\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__33915\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\
        );

    \I__6765\ : InMux
    port map (
            O => \N__33912\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__6764\ : InMux
    port map (
            O => \N__33909\,
            I => \N__33906\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__33906\,
            I => \N__33903\
        );

    \I__6762\ : Span4Mux_v
    port map (
            O => \N__33903\,
            I => \N__33897\
        );

    \I__6761\ : InMux
    port map (
            O => \N__33902\,
            I => \N__33894\
        );

    \I__6760\ : InMux
    port map (
            O => \N__33901\,
            I => \N__33889\
        );

    \I__6759\ : InMux
    port map (
            O => \N__33900\,
            I => \N__33889\
        );

    \I__6758\ : Odrv4
    port map (
            O => \N__33897\,
            I => \delay_measurement_inst.delay_tr_timer.N_296\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__33894\,
            I => \delay_measurement_inst.delay_tr_timer.N_296\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__33889\,
            I => \delay_measurement_inst.delay_tr_timer.N_296\
        );

    \I__6755\ : CascadeMux
    port map (
            O => \N__33882\,
            I => \delay_measurement_inst.delay_tr_timer.N_293_cascade_\
        );

    \I__6754\ : InMux
    port map (
            O => \N__33879\,
            I => \N__33876\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__33876\,
            I => \N__33873\
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__33873\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\
        );

    \I__6751\ : InMux
    port map (
            O => \N__33870\,
            I => \N__33867\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__33867\,
            I => \N__33864\
        );

    \I__6749\ : Odrv12
    port map (
            O => \N__33864\,
            I => \delay_measurement_inst.N_307\
        );

    \I__6748\ : IoInMux
    port map (
            O => \N__33861\,
            I => \N__33858\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__33858\,
            I => \N__33855\
        );

    \I__6746\ : Odrv4
    port map (
            O => \N__33855\,
            I => s2_phy_c
        );

    \I__6745\ : IoInMux
    port map (
            O => \N__33852\,
            I => \N__33849\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__33849\,
            I => \N__33846\
        );

    \I__6743\ : Span4Mux_s3_v
    port map (
            O => \N__33846\,
            I => \N__33843\
        );

    \I__6742\ : Odrv4
    port map (
            O => \N__33843\,
            I => \delay_measurement_inst.delay_hc_timer.N_335_i\
        );

    \I__6741\ : InMux
    port map (
            O => \N__33840\,
            I => \N__33837\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__33837\,
            I => \N__33834\
        );

    \I__6739\ : Span4Mux_h
    port map (
            O => \N__33834\,
            I => \N__33831\
        );

    \I__6738\ : Odrv4
    port map (
            O => \N__33831\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\
        );

    \I__6737\ : CascadeMux
    port map (
            O => \N__33828\,
            I => \N__33825\
        );

    \I__6736\ : InMux
    port map (
            O => \N__33825\,
            I => \N__33821\
        );

    \I__6735\ : InMux
    port map (
            O => \N__33824\,
            I => \N__33817\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__33821\,
            I => \N__33814\
        );

    \I__6733\ : InMux
    port map (
            O => \N__33820\,
            I => \N__33811\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__33817\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6731\ : Odrv4
    port map (
            O => \N__33814\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__33811\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6729\ : InMux
    port map (
            O => \N__33804\,
            I => \N__33800\
        );

    \I__6728\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33797\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__33800\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__33797\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__6725\ : InMux
    port map (
            O => \N__33792\,
            I => \N__33789\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__33789\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\
        );

    \I__6723\ : InMux
    port map (
            O => \N__33786\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__6722\ : InMux
    port map (
            O => \N__33783\,
            I => \N__33780\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__33780\,
            I => \N__33777\
        );

    \I__6720\ : Span4Mux_h
    port map (
            O => \N__33777\,
            I => \N__33774\
        );

    \I__6719\ : Odrv4
    port map (
            O => \N__33774\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\
        );

    \I__6718\ : CascadeMux
    port map (
            O => \N__33771\,
            I => \N__33768\
        );

    \I__6717\ : InMux
    port map (
            O => \N__33768\,
            I => \N__33764\
        );

    \I__6716\ : InMux
    port map (
            O => \N__33767\,
            I => \N__33761\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__33764\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__33761\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__6713\ : CascadeMux
    port map (
            O => \N__33756\,
            I => \N__33753\
        );

    \I__6712\ : InMux
    port map (
            O => \N__33753\,
            I => \N__33750\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__33750\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\
        );

    \I__6710\ : CascadeMux
    port map (
            O => \N__33747\,
            I => \delay_measurement_inst.N_358_cascade_\
        );

    \I__6709\ : InMux
    port map (
            O => \N__33744\,
            I => \N__33739\
        );

    \I__6708\ : InMux
    port map (
            O => \N__33743\,
            I => \N__33736\
        );

    \I__6707\ : InMux
    port map (
            O => \N__33742\,
            I => \N__33733\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__33739\,
            I => \N__33730\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__33736\,
            I => \N__33726\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__33733\,
            I => \N__33721\
        );

    \I__6703\ : Span12Mux_h
    port map (
            O => \N__33730\,
            I => \N__33721\
        );

    \I__6702\ : InMux
    port map (
            O => \N__33729\,
            I => \N__33718\
        );

    \I__6701\ : Span12Mux_v
    port map (
            O => \N__33726\,
            I => \N__33715\
        );

    \I__6700\ : Span12Mux_v
    port map (
            O => \N__33721\,
            I => \N__33712\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__33718\,
            I => \current_shift_inst.stop_timer_phaseZ0\
        );

    \I__6698\ : Odrv12
    port map (
            O => \N__33715\,
            I => \current_shift_inst.stop_timer_phaseZ0\
        );

    \I__6697\ : Odrv12
    port map (
            O => \N__33712\,
            I => \current_shift_inst.stop_timer_phaseZ0\
        );

    \I__6696\ : InMux
    port map (
            O => \N__33705\,
            I => \N__33702\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__33702\,
            I => \N__33698\
        );

    \I__6694\ : InMux
    port map (
            O => \N__33701\,
            I => \N__33695\
        );

    \I__6693\ : Span4Mux_h
    port map (
            O => \N__33698\,
            I => \N__33690\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__33695\,
            I => \N__33690\
        );

    \I__6691\ : Span4Mux_v
    port map (
            O => \N__33690\,
            I => \N__33686\
        );

    \I__6690\ : InMux
    port map (
            O => \N__33689\,
            I => \N__33683\
        );

    \I__6689\ : Span4Mux_v
    port map (
            O => \N__33686\,
            I => \N__33680\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__33683\,
            I => \current_shift_inst.start_timer_phaseZ0\
        );

    \I__6687\ : Odrv4
    port map (
            O => \N__33680\,
            I => \current_shift_inst.start_timer_phaseZ0\
        );

    \I__6686\ : InMux
    port map (
            O => \N__33675\,
            I => \N__33670\
        );

    \I__6685\ : InMux
    port map (
            O => \N__33674\,
            I => \N__33667\
        );

    \I__6684\ : InMux
    port map (
            O => \N__33673\,
            I => \N__33663\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__33670\,
            I => \N__33660\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__33667\,
            I => \N__33657\
        );

    \I__6681\ : InMux
    port map (
            O => \N__33666\,
            I => \N__33654\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__33663\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__6679\ : Odrv12
    port map (
            O => \N__33660\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__6678\ : Odrv4
    port map (
            O => \N__33657\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__33654\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__6676\ : CEMux
    port map (
            O => \N__33645\,
            I => \N__33642\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__33642\,
            I => \N__33636\
        );

    \I__6674\ : CEMux
    port map (
            O => \N__33641\,
            I => \N__33633\
        );

    \I__6673\ : CEMux
    port map (
            O => \N__33640\,
            I => \N__33630\
        );

    \I__6672\ : CEMux
    port map (
            O => \N__33639\,
            I => \N__33627\
        );

    \I__6671\ : Span4Mux_v
    port map (
            O => \N__33636\,
            I => \N__33624\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__33633\,
            I => \N__33619\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__33630\,
            I => \N__33619\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__33627\,
            I => \N__33616\
        );

    \I__6667\ : Span4Mux_h
    port map (
            O => \N__33624\,
            I => \N__33611\
        );

    \I__6666\ : Span4Mux_v
    port map (
            O => \N__33619\,
            I => \N__33611\
        );

    \I__6665\ : Span4Mux_h
    port map (
            O => \N__33616\,
            I => \N__33608\
        );

    \I__6664\ : Span4Mux_h
    port map (
            O => \N__33611\,
            I => \N__33605\
        );

    \I__6663\ : Span4Mux_h
    port map (
            O => \N__33608\,
            I => \N__33602\
        );

    \I__6662\ : Odrv4
    port map (
            O => \N__33605\,
            I => \current_shift_inst.timer_phase.N_192_i\
        );

    \I__6661\ : Odrv4
    port map (
            O => \N__33602\,
            I => \current_shift_inst.timer_phase.N_192_i\
        );

    \I__6660\ : InMux
    port map (
            O => \N__33597\,
            I => \N__33594\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__33594\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19\
        );

    \I__6658\ : InMux
    port map (
            O => \N__33591\,
            I => \N__33588\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__33588\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\
        );

    \I__6656\ : InMux
    port map (
            O => \N__33585\,
            I => \N__33579\
        );

    \I__6655\ : InMux
    port map (
            O => \N__33584\,
            I => \N__33579\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__33579\,
            I => \delay_measurement_inst.delay_tr_timer.N_320_4\
        );

    \I__6653\ : CascadeMux
    port map (
            O => \N__33576\,
            I => \delay_measurement_inst.N_305_1_cascade_\
        );

    \I__6652\ : CascadeMux
    port map (
            O => \N__33573\,
            I => \N__33568\
        );

    \I__6651\ : InMux
    port map (
            O => \N__33572\,
            I => \N__33558\
        );

    \I__6650\ : InMux
    port map (
            O => \N__33571\,
            I => \N__33558\
        );

    \I__6649\ : InMux
    port map (
            O => \N__33568\,
            I => \N__33558\
        );

    \I__6648\ : InMux
    port map (
            O => \N__33567\,
            I => \N__33558\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__33558\,
            I => \delay_measurement_inst.N_305_1\
        );

    \I__6646\ : InMux
    port map (
            O => \N__33555\,
            I => \N__33551\
        );

    \I__6645\ : InMux
    port map (
            O => \N__33554\,
            I => \N__33548\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__33551\,
            I => \N__33545\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__33548\,
            I => \delay_measurement_inst.delay_tr_timer.N_299\
        );

    \I__6642\ : Odrv12
    port map (
            O => \N__33545\,
            I => \delay_measurement_inst.delay_tr_timer.N_299\
        );

    \I__6641\ : CascadeMux
    port map (
            O => \N__33540\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5_cascade_\
        );

    \I__6640\ : CascadeMux
    port map (
            O => \N__33537\,
            I => \delay_measurement_inst.delay_tr_timer.N_321_cascade_\
        );

    \I__6639\ : CascadeMux
    port map (
            O => \N__33534\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6_cascade_\
        );

    \I__6638\ : InMux
    port map (
            O => \N__33531\,
            I => \N__33528\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__33528\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7\
        );

    \I__6636\ : InMux
    port map (
            O => \N__33525\,
            I => \N__33522\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__33522\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3\
        );

    \I__6634\ : CascadeMux
    port map (
            O => \N__33519\,
            I => \N__33516\
        );

    \I__6633\ : InMux
    port map (
            O => \N__33516\,
            I => \N__33513\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__33513\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3\
        );

    \I__6631\ : InMux
    port map (
            O => \N__33510\,
            I => \N__33507\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__33507\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_12\
        );

    \I__6629\ : InMux
    port map (
            O => \N__33504\,
            I => \N__33501\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__33501\,
            I => \N__33498\
        );

    \I__6627\ : Span4Mux_h
    port map (
            O => \N__33498\,
            I => \N__33495\
        );

    \I__6626\ : Odrv4
    port map (
            O => \N__33495\,
            I => \current_shift_inst.un4_control_input_axb_12\
        );

    \I__6625\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33489\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__33489\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_18\
        );

    \I__6623\ : InMux
    port map (
            O => \N__33486\,
            I => \N__33483\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__33483\,
            I => \N__33480\
        );

    \I__6621\ : Span4Mux_h
    port map (
            O => \N__33480\,
            I => \N__33477\
        );

    \I__6620\ : Odrv4
    port map (
            O => \N__33477\,
            I => \current_shift_inst.un4_control_input_axb_18\
        );

    \I__6619\ : InMux
    port map (
            O => \N__33474\,
            I => \N__33471\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__33471\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_13\
        );

    \I__6617\ : InMux
    port map (
            O => \N__33468\,
            I => \N__33465\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__33465\,
            I => \N__33462\
        );

    \I__6615\ : Span4Mux_v
    port map (
            O => \N__33462\,
            I => \N__33459\
        );

    \I__6614\ : Odrv4
    port map (
            O => \N__33459\,
            I => \current_shift_inst.un4_control_input_axb_13\
        );

    \I__6613\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33453\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__33453\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_14\
        );

    \I__6611\ : InMux
    port map (
            O => \N__33450\,
            I => \N__33447\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__33447\,
            I => \N__33444\
        );

    \I__6609\ : Span4Mux_h
    port map (
            O => \N__33444\,
            I => \N__33441\
        );

    \I__6608\ : Odrv4
    port map (
            O => \N__33441\,
            I => \current_shift_inst.un4_control_input_axb_14\
        );

    \I__6607\ : InMux
    port map (
            O => \N__33438\,
            I => \N__33435\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__33435\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_23\
        );

    \I__6605\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33429\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__33429\,
            I => \N__33426\
        );

    \I__6603\ : Span4Mux_h
    port map (
            O => \N__33426\,
            I => \N__33423\
        );

    \I__6602\ : Odrv4
    port map (
            O => \N__33423\,
            I => \current_shift_inst.un4_control_input_axb_23\
        );

    \I__6601\ : InMux
    port map (
            O => \N__33420\,
            I => \N__33417\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__33417\,
            I => \N__33414\
        );

    \I__6599\ : Span4Mux_v
    port map (
            O => \N__33414\,
            I => \N__33411\
        );

    \I__6598\ : Odrv4
    port map (
            O => \N__33411\,
            I => \current_shift_inst.un4_control_input_axb_15\
        );

    \I__6597\ : InMux
    port map (
            O => \N__33408\,
            I => \N__33405\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__33405\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_16\
        );

    \I__6595\ : InMux
    port map (
            O => \N__33402\,
            I => \N__33399\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__33399\,
            I => \N__33396\
        );

    \I__6593\ : Span4Mux_h
    port map (
            O => \N__33396\,
            I => \N__33393\
        );

    \I__6592\ : Odrv4
    port map (
            O => \N__33393\,
            I => \current_shift_inst.un4_control_input_axb_16\
        );

    \I__6591\ : InMux
    port map (
            O => \N__33390\,
            I => \N__33387\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__33387\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_17\
        );

    \I__6589\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33381\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__33381\,
            I => \N__33378\
        );

    \I__6587\ : Span4Mux_v
    port map (
            O => \N__33378\,
            I => \N__33375\
        );

    \I__6586\ : Odrv4
    port map (
            O => \N__33375\,
            I => \current_shift_inst.un4_control_input_axb_17\
        );

    \I__6585\ : InMux
    port map (
            O => \N__33372\,
            I => \N__33366\
        );

    \I__6584\ : InMux
    port map (
            O => \N__33371\,
            I => \N__33361\
        );

    \I__6583\ : InMux
    port map (
            O => \N__33370\,
            I => \N__33361\
        );

    \I__6582\ : InMux
    port map (
            O => \N__33369\,
            I => \N__33358\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__33366\,
            I => \N__33355\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__33361\,
            I => \N__33352\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__33358\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6578\ : Odrv12
    port map (
            O => \N__33355\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6577\ : Odrv4
    port map (
            O => \N__33352\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6576\ : InMux
    port map (
            O => \N__33345\,
            I => \N__33323\
        );

    \I__6575\ : InMux
    port map (
            O => \N__33344\,
            I => \N__33323\
        );

    \I__6574\ : InMux
    port map (
            O => \N__33343\,
            I => \N__33323\
        );

    \I__6573\ : InMux
    port map (
            O => \N__33342\,
            I => \N__33323\
        );

    \I__6572\ : InMux
    port map (
            O => \N__33341\,
            I => \N__33302\
        );

    \I__6571\ : InMux
    port map (
            O => \N__33340\,
            I => \N__33302\
        );

    \I__6570\ : InMux
    port map (
            O => \N__33339\,
            I => \N__33293\
        );

    \I__6569\ : InMux
    port map (
            O => \N__33338\,
            I => \N__33293\
        );

    \I__6568\ : InMux
    port map (
            O => \N__33337\,
            I => \N__33293\
        );

    \I__6567\ : InMux
    port map (
            O => \N__33336\,
            I => \N__33293\
        );

    \I__6566\ : InMux
    port map (
            O => \N__33335\,
            I => \N__33284\
        );

    \I__6565\ : InMux
    port map (
            O => \N__33334\,
            I => \N__33284\
        );

    \I__6564\ : InMux
    port map (
            O => \N__33333\,
            I => \N__33284\
        );

    \I__6563\ : InMux
    port map (
            O => \N__33332\,
            I => \N__33284\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__33323\,
            I => \N__33281\
        );

    \I__6561\ : InMux
    port map (
            O => \N__33322\,
            I => \N__33272\
        );

    \I__6560\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33272\
        );

    \I__6559\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33272\
        );

    \I__6558\ : InMux
    port map (
            O => \N__33319\,
            I => \N__33272\
        );

    \I__6557\ : InMux
    port map (
            O => \N__33318\,
            I => \N__33263\
        );

    \I__6556\ : InMux
    port map (
            O => \N__33317\,
            I => \N__33263\
        );

    \I__6555\ : InMux
    port map (
            O => \N__33316\,
            I => \N__33263\
        );

    \I__6554\ : InMux
    port map (
            O => \N__33315\,
            I => \N__33263\
        );

    \I__6553\ : InMux
    port map (
            O => \N__33314\,
            I => \N__33254\
        );

    \I__6552\ : InMux
    port map (
            O => \N__33313\,
            I => \N__33254\
        );

    \I__6551\ : InMux
    port map (
            O => \N__33312\,
            I => \N__33254\
        );

    \I__6550\ : InMux
    port map (
            O => \N__33311\,
            I => \N__33254\
        );

    \I__6549\ : InMux
    port map (
            O => \N__33310\,
            I => \N__33245\
        );

    \I__6548\ : InMux
    port map (
            O => \N__33309\,
            I => \N__33245\
        );

    \I__6547\ : InMux
    port map (
            O => \N__33308\,
            I => \N__33245\
        );

    \I__6546\ : InMux
    port map (
            O => \N__33307\,
            I => \N__33245\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__33302\,
            I => \N__33242\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__33293\,
            I => \N__33239\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__33284\,
            I => \N__33236\
        );

    \I__6542\ : Span4Mux_h
    port map (
            O => \N__33281\,
            I => \N__33221\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__33272\,
            I => \N__33221\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__33263\,
            I => \N__33221\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__33254\,
            I => \N__33221\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__33245\,
            I => \N__33221\
        );

    \I__6537\ : Span4Mux_v
    port map (
            O => \N__33242\,
            I => \N__33221\
        );

    \I__6536\ : Span4Mux_v
    port map (
            O => \N__33239\,
            I => \N__33221\
        );

    \I__6535\ : Span4Mux_v
    port map (
            O => \N__33236\,
            I => \N__33216\
        );

    \I__6534\ : Span4Mux_v
    port map (
            O => \N__33221\,
            I => \N__33216\
        );

    \I__6533\ : Odrv4
    port map (
            O => \N__33216\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__6532\ : InMux
    port map (
            O => \N__33213\,
            I => \N__33210\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__33210\,
            I => \N__33207\
        );

    \I__6530\ : Odrv4
    port map (
            O => \N__33207\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_21\
        );

    \I__6529\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33201\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__33201\,
            I => \N__33198\
        );

    \I__6527\ : Span4Mux_v
    port map (
            O => \N__33198\,
            I => \N__33195\
        );

    \I__6526\ : Odrv4
    port map (
            O => \N__33195\,
            I => \current_shift_inst.un4_control_input_axb_21\
        );

    \I__6525\ : InMux
    port map (
            O => \N__33192\,
            I => \N__33189\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__33189\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_10\
        );

    \I__6523\ : InMux
    port map (
            O => \N__33186\,
            I => \N__33183\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__33183\,
            I => \N__33180\
        );

    \I__6521\ : Span4Mux_v
    port map (
            O => \N__33180\,
            I => \N__33177\
        );

    \I__6520\ : Odrv4
    port map (
            O => \N__33177\,
            I => \current_shift_inst.un4_control_input_axb_10\
        );

    \I__6519\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33171\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__33171\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_11\
        );

    \I__6517\ : InMux
    port map (
            O => \N__33168\,
            I => \N__33165\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__33165\,
            I => \N__33162\
        );

    \I__6515\ : Span4Mux_v
    port map (
            O => \N__33162\,
            I => \N__33159\
        );

    \I__6514\ : Odrv4
    port map (
            O => \N__33159\,
            I => \current_shift_inst.un4_control_input_axb_11\
        );

    \I__6513\ : CascadeMux
    port map (
            O => \N__33156\,
            I => \N__33151\
        );

    \I__6512\ : CascadeMux
    port map (
            O => \N__33155\,
            I => \N__33148\
        );

    \I__6511\ : InMux
    port map (
            O => \N__33154\,
            I => \N__33145\
        );

    \I__6510\ : InMux
    port map (
            O => \N__33151\,
            I => \N__33142\
        );

    \I__6509\ : InMux
    port map (
            O => \N__33148\,
            I => \N__33137\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__33145\,
            I => \N__33134\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__33142\,
            I => \N__33131\
        );

    \I__6506\ : InMux
    port map (
            O => \N__33141\,
            I => \N__33126\
        );

    \I__6505\ : InMux
    port map (
            O => \N__33140\,
            I => \N__33126\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__33137\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6503\ : Odrv4
    port map (
            O => \N__33134\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6502\ : Odrv4
    port map (
            O => \N__33131\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__33126\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6500\ : InMux
    port map (
            O => \N__33117\,
            I => \N__33111\
        );

    \I__6499\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33108\
        );

    \I__6498\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33103\
        );

    \I__6497\ : InMux
    port map (
            O => \N__33114\,
            I => \N__33103\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__33111\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__33108\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__33103\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6493\ : InMux
    port map (
            O => \N__33096\,
            I => \N__33092\
        );

    \I__6492\ : InMux
    port map (
            O => \N__33095\,
            I => \N__33089\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__33092\,
            I => \N__33085\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__33089\,
            I => \N__33082\
        );

    \I__6489\ : InMux
    port map (
            O => \N__33088\,
            I => \N__33079\
        );

    \I__6488\ : Odrv4
    port map (
            O => \N__33085\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__33082\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__33079\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__6485\ : InMux
    port map (
            O => \N__33072\,
            I => \N__33069\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__33069\,
            I => \N__33065\
        );

    \I__6483\ : InMux
    port map (
            O => \N__33068\,
            I => \N__33062\
        );

    \I__6482\ : Span4Mux_h
    port map (
            O => \N__33065\,
            I => \N__33058\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__33062\,
            I => \N__33055\
        );

    \I__6480\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33052\
        );

    \I__6479\ : Odrv4
    port map (
            O => \N__33058\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__6478\ : Odrv4
    port map (
            O => \N__33055\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__33052\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__6476\ : InMux
    port map (
            O => \N__33045\,
            I => \N__33041\
        );

    \I__6475\ : InMux
    port map (
            O => \N__33044\,
            I => \N__33037\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__33041\,
            I => \N__33034\
        );

    \I__6473\ : InMux
    port map (
            O => \N__33040\,
            I => \N__33031\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__33037\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6471\ : Odrv4
    port map (
            O => \N__33034\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__33031\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6469\ : CEMux
    port map (
            O => \N__33024\,
            I => \N__33021\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__33021\,
            I => \N__33018\
        );

    \I__6467\ : Sp12to4
    port map (
            O => \N__33018\,
            I => \N__33015\
        );

    \I__6466\ : Odrv12
    port map (
            O => \N__33015\,
            I => \phase_controller_inst1.N_221_0\
        );

    \I__6465\ : InMux
    port map (
            O => \N__33012\,
            I => \N__33006\
        );

    \I__6464\ : InMux
    port map (
            O => \N__33011\,
            I => \N__33006\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__33006\,
            I => \N__33003\
        );

    \I__6462\ : Odrv4
    port map (
            O => \N__33003\,
            I => \current_shift_inst.S3_syncZ0Z1\
        );

    \I__6461\ : InMux
    port map (
            O => \N__33000\,
            I => \N__32997\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__32997\,
            I => \current_shift_inst.S3_syncZ0Z0\
        );

    \I__6459\ : InMux
    port map (
            O => \N__32994\,
            I => \N__32991\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__32991\,
            I => \N__32988\
        );

    \I__6457\ : Odrv4
    port map (
            O => \N__32988\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_24\
        );

    \I__6456\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32982\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__32982\,
            I => \N__32979\
        );

    \I__6454\ : Span4Mux_v
    port map (
            O => \N__32979\,
            I => \N__32976\
        );

    \I__6453\ : Odrv4
    port map (
            O => \N__32976\,
            I => \current_shift_inst.un4_control_input_axb_24\
        );

    \I__6452\ : InMux
    port map (
            O => \N__32973\,
            I => \N__32970\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__32970\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_15\
        );

    \I__6450\ : CascadeMux
    port map (
            O => \N__32967\,
            I => \N__32963\
        );

    \I__6449\ : InMux
    port map (
            O => \N__32966\,
            I => \N__32960\
        );

    \I__6448\ : InMux
    port map (
            O => \N__32963\,
            I => \N__32957\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__32960\,
            I => \N__32954\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__32957\,
            I => measured_delay_hc_26
        );

    \I__6445\ : Odrv4
    port map (
            O => \N__32954\,
            I => measured_delay_hc_26
        );

    \I__6444\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32945\
        );

    \I__6443\ : InMux
    port map (
            O => \N__32948\,
            I => \N__32942\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__32945\,
            I => \N__32939\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__32942\,
            I => measured_delay_hc_24
        );

    \I__6440\ : Odrv4
    port map (
            O => \N__32939\,
            I => measured_delay_hc_24
        );

    \I__6439\ : IoInMux
    port map (
            O => \N__32934\,
            I => \N__32931\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__32931\,
            I => \N__32928\
        );

    \I__6437\ : IoSpan4Mux
    port map (
            O => \N__32928\,
            I => \N__32925\
        );

    \I__6436\ : Span4Mux_s1_v
    port map (
            O => \N__32925\,
            I => \N__32921\
        );

    \I__6435\ : InMux
    port map (
            O => \N__32924\,
            I => \N__32918\
        );

    \I__6434\ : Sp12to4
    port map (
            O => \N__32921\,
            I => \N__32915\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__32918\,
            I => \N__32912\
        );

    \I__6432\ : Span12Mux_s8_v
    port map (
            O => \N__32915\,
            I => \N__32909\
        );

    \I__6431\ : Span4Mux_v
    port map (
            O => \N__32912\,
            I => \N__32906\
        );

    \I__6430\ : Odrv12
    port map (
            O => \N__32909\,
            I => s1_phy_c
        );

    \I__6429\ : Odrv4
    port map (
            O => \N__32906\,
            I => s1_phy_c
        );

    \I__6428\ : InMux
    port map (
            O => \N__32901\,
            I => \N__32898\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__32898\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__6426\ : InMux
    port map (
            O => \N__32895\,
            I => \N__32891\
        );

    \I__6425\ : CascadeMux
    port map (
            O => \N__32894\,
            I => \N__32888\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__32891\,
            I => \N__32885\
        );

    \I__6423\ : InMux
    port map (
            O => \N__32888\,
            I => \N__32882\
        );

    \I__6422\ : Span4Mux_h
    port map (
            O => \N__32885\,
            I => \N__32879\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__32882\,
            I => measured_delay_hc_25
        );

    \I__6420\ : Odrv4
    port map (
            O => \N__32879\,
            I => measured_delay_hc_25
        );

    \I__6419\ : InMux
    port map (
            O => \N__32874\,
            I => \N__32840\
        );

    \I__6418\ : InMux
    port map (
            O => \N__32873\,
            I => \N__32840\
        );

    \I__6417\ : InMux
    port map (
            O => \N__32872\,
            I => \N__32840\
        );

    \I__6416\ : InMux
    port map (
            O => \N__32871\,
            I => \N__32840\
        );

    \I__6415\ : InMux
    port map (
            O => \N__32870\,
            I => \N__32840\
        );

    \I__6414\ : InMux
    port map (
            O => \N__32869\,
            I => \N__32840\
        );

    \I__6413\ : InMux
    port map (
            O => \N__32868\,
            I => \N__32840\
        );

    \I__6412\ : InMux
    port map (
            O => \N__32867\,
            I => \N__32825\
        );

    \I__6411\ : InMux
    port map (
            O => \N__32866\,
            I => \N__32825\
        );

    \I__6410\ : InMux
    port map (
            O => \N__32865\,
            I => \N__32825\
        );

    \I__6409\ : InMux
    port map (
            O => \N__32864\,
            I => \N__32825\
        );

    \I__6408\ : InMux
    port map (
            O => \N__32863\,
            I => \N__32825\
        );

    \I__6407\ : InMux
    port map (
            O => \N__32862\,
            I => \N__32825\
        );

    \I__6406\ : InMux
    port map (
            O => \N__32861\,
            I => \N__32825\
        );

    \I__6405\ : InMux
    port map (
            O => \N__32860\,
            I => \N__32814\
        );

    \I__6404\ : InMux
    port map (
            O => \N__32859\,
            I => \N__32814\
        );

    \I__6403\ : InMux
    port map (
            O => \N__32858\,
            I => \N__32814\
        );

    \I__6402\ : InMux
    port map (
            O => \N__32857\,
            I => \N__32814\
        );

    \I__6401\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32814\
        );

    \I__6400\ : InMux
    port map (
            O => \N__32855\,
            I => \N__32809\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__32840\,
            I => \N__32804\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__32825\,
            I => \N__32804\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__32814\,
            I => \N__32800\
        );

    \I__6396\ : InMux
    port map (
            O => \N__32813\,
            I => \N__32797\
        );

    \I__6395\ : InMux
    port map (
            O => \N__32812\,
            I => \N__32793\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__32809\,
            I => \N__32790\
        );

    \I__6393\ : Span4Mux_v
    port map (
            O => \N__32804\,
            I => \N__32787\
        );

    \I__6392\ : InMux
    port map (
            O => \N__32803\,
            I => \N__32784\
        );

    \I__6391\ : Span4Mux_h
    port map (
            O => \N__32800\,
            I => \N__32779\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__32797\,
            I => \N__32779\
        );

    \I__6389\ : InMux
    port map (
            O => \N__32796\,
            I => \N__32776\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__32793\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__6387\ : Odrv4
    port map (
            O => \N__32790\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__6386\ : Odrv4
    port map (
            O => \N__32787\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__32784\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__6384\ : Odrv4
    port map (
            O => \N__32779\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__32776\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__6382\ : CascadeMux
    port map (
            O => \N__32763\,
            I => \N__32757\
        );

    \I__6381\ : CascadeMux
    port map (
            O => \N__32762\,
            I => \N__32754\
        );

    \I__6380\ : CascadeMux
    port map (
            O => \N__32761\,
            I => \N__32751\
        );

    \I__6379\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32732\
        );

    \I__6378\ : InMux
    port map (
            O => \N__32757\,
            I => \N__32722\
        );

    \I__6377\ : InMux
    port map (
            O => \N__32754\,
            I => \N__32722\
        );

    \I__6376\ : InMux
    port map (
            O => \N__32751\,
            I => \N__32722\
        );

    \I__6375\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32719\
        );

    \I__6374\ : InMux
    port map (
            O => \N__32749\,
            I => \N__32704\
        );

    \I__6373\ : InMux
    port map (
            O => \N__32748\,
            I => \N__32704\
        );

    \I__6372\ : InMux
    port map (
            O => \N__32747\,
            I => \N__32704\
        );

    \I__6371\ : InMux
    port map (
            O => \N__32746\,
            I => \N__32704\
        );

    \I__6370\ : InMux
    port map (
            O => \N__32745\,
            I => \N__32704\
        );

    \I__6369\ : InMux
    port map (
            O => \N__32744\,
            I => \N__32704\
        );

    \I__6368\ : InMux
    port map (
            O => \N__32743\,
            I => \N__32704\
        );

    \I__6367\ : InMux
    port map (
            O => \N__32742\,
            I => \N__32689\
        );

    \I__6366\ : InMux
    port map (
            O => \N__32741\,
            I => \N__32689\
        );

    \I__6365\ : InMux
    port map (
            O => \N__32740\,
            I => \N__32689\
        );

    \I__6364\ : InMux
    port map (
            O => \N__32739\,
            I => \N__32689\
        );

    \I__6363\ : InMux
    port map (
            O => \N__32738\,
            I => \N__32689\
        );

    \I__6362\ : InMux
    port map (
            O => \N__32737\,
            I => \N__32689\
        );

    \I__6361\ : InMux
    port map (
            O => \N__32736\,
            I => \N__32689\
        );

    \I__6360\ : InMux
    port map (
            O => \N__32735\,
            I => \N__32686\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__32732\,
            I => \N__32683\
        );

    \I__6358\ : InMux
    port map (
            O => \N__32731\,
            I => \N__32679\
        );

    \I__6357\ : InMux
    port map (
            O => \N__32730\,
            I => \N__32674\
        );

    \I__6356\ : InMux
    port map (
            O => \N__32729\,
            I => \N__32674\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__32722\,
            I => \N__32669\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__32719\,
            I => \N__32669\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__32704\,
            I => \N__32666\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__32689\,
            I => \N__32663\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__32686\,
            I => \N__32658\
        );

    \I__6350\ : Span4Mux_v
    port map (
            O => \N__32683\,
            I => \N__32658\
        );

    \I__6349\ : InMux
    port map (
            O => \N__32682\,
            I => \N__32655\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__32679\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__32674\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__6346\ : Odrv4
    port map (
            O => \N__32669\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__6345\ : Odrv4
    port map (
            O => \N__32666\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__6344\ : Odrv4
    port map (
            O => \N__32663\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__6343\ : Odrv4
    port map (
            O => \N__32658\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__32655\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__6341\ : InMux
    port map (
            O => \N__32640\,
            I => \N__32637\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__32637\,
            I => \N__32634\
        );

    \I__6339\ : Glb2LocalMux
    port map (
            O => \N__32634\,
            I => \N__32631\
        );

    \I__6338\ : GlobalMux
    port map (
            O => \N__32631\,
            I => clk_12mhz
        );

    \I__6337\ : IoInMux
    port map (
            O => \N__32628\,
            I => \N__32625\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__32625\,
            I => \N__32622\
        );

    \I__6335\ : Span4Mux_s0_v
    port map (
            O => \N__32622\,
            I => \N__32619\
        );

    \I__6334\ : Odrv4
    port map (
            O => \N__32619\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__6333\ : InMux
    port map (
            O => \N__32616\,
            I => \N__32613\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__32613\,
            I => \N__32610\
        );

    \I__6331\ : Span4Mux_v
    port map (
            O => \N__32610\,
            I => \N__32607\
        );

    \I__6330\ : Span4Mux_h
    port map (
            O => \N__32607\,
            I => \N__32604\
        );

    \I__6329\ : Span4Mux_h
    port map (
            O => \N__32604\,
            I => \N__32601\
        );

    \I__6328\ : Odrv4
    port map (
            O => \N__32601\,
            I => il_max_comp2_c
        );

    \I__6327\ : InMux
    port map (
            O => \N__32598\,
            I => \N__32595\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__32595\,
            I => \il_max_comp2_D1\
        );

    \I__6325\ : CascadeMux
    port map (
            O => \N__32592\,
            I => \N__32588\
        );

    \I__6324\ : CascadeMux
    port map (
            O => \N__32591\,
            I => \N__32585\
        );

    \I__6323\ : InMux
    port map (
            O => \N__32588\,
            I => \N__32580\
        );

    \I__6322\ : InMux
    port map (
            O => \N__32585\,
            I => \N__32580\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__32580\,
            I => \N__32576\
        );

    \I__6320\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32573\
        );

    \I__6319\ : Span4Mux_v
    port map (
            O => \N__32576\,
            I => \N__32570\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__32573\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__6317\ : Odrv4
    port map (
            O => \N__32570\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__6316\ : InMux
    port map (
            O => \N__32565\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__6315\ : InMux
    port map (
            O => \N__32562\,
            I => \N__32558\
        );

    \I__6314\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32555\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__32558\,
            I => \N__32549\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__32555\,
            I => \N__32549\
        );

    \I__6311\ : InMux
    port map (
            O => \N__32554\,
            I => \N__32546\
        );

    \I__6310\ : Span4Mux_v
    port map (
            O => \N__32549\,
            I => \N__32543\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__32546\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__6308\ : Odrv4
    port map (
            O => \N__32543\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__6307\ : InMux
    port map (
            O => \N__32538\,
            I => \bfn_12_22_0_\
        );

    \I__6306\ : CascadeMux
    port map (
            O => \N__32535\,
            I => \N__32532\
        );

    \I__6305\ : InMux
    port map (
            O => \N__32532\,
            I => \N__32528\
        );

    \I__6304\ : InMux
    port map (
            O => \N__32531\,
            I => \N__32525\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__32528\,
            I => \N__32519\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__32525\,
            I => \N__32519\
        );

    \I__6301\ : InMux
    port map (
            O => \N__32524\,
            I => \N__32516\
        );

    \I__6300\ : Span4Mux_v
    port map (
            O => \N__32519\,
            I => \N__32513\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__32516\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__6298\ : Odrv4
    port map (
            O => \N__32513\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__6297\ : InMux
    port map (
            O => \N__32508\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__6296\ : CascadeMux
    port map (
            O => \N__32505\,
            I => \N__32501\
        );

    \I__6295\ : CascadeMux
    port map (
            O => \N__32504\,
            I => \N__32498\
        );

    \I__6294\ : InMux
    port map (
            O => \N__32501\,
            I => \N__32493\
        );

    \I__6293\ : InMux
    port map (
            O => \N__32498\,
            I => \N__32493\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__32493\,
            I => \N__32489\
        );

    \I__6291\ : InMux
    port map (
            O => \N__32492\,
            I => \N__32486\
        );

    \I__6290\ : Span4Mux_v
    port map (
            O => \N__32489\,
            I => \N__32483\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__32486\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__6288\ : Odrv4
    port map (
            O => \N__32483\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__6287\ : InMux
    port map (
            O => \N__32478\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__6286\ : InMux
    port map (
            O => \N__32475\,
            I => \N__32468\
        );

    \I__6285\ : InMux
    port map (
            O => \N__32474\,
            I => \N__32468\
        );

    \I__6284\ : InMux
    port map (
            O => \N__32473\,
            I => \N__32465\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__32468\,
            I => \N__32462\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__32465\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__6281\ : Odrv12
    port map (
            O => \N__32462\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__6280\ : InMux
    port map (
            O => \N__32457\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__6279\ : InMux
    port map (
            O => \N__32454\,
            I => \N__32451\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__32451\,
            I => \N__32447\
        );

    \I__6277\ : InMux
    port map (
            O => \N__32450\,
            I => \N__32444\
        );

    \I__6276\ : Span4Mux_v
    port map (
            O => \N__32447\,
            I => \N__32441\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__32444\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__6274\ : Odrv4
    port map (
            O => \N__32441\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__6273\ : InMux
    port map (
            O => \N__32436\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__6272\ : InMux
    port map (
            O => \N__32433\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__6271\ : CascadeMux
    port map (
            O => \N__32430\,
            I => \N__32427\
        );

    \I__6270\ : InMux
    port map (
            O => \N__32427\,
            I => \N__32423\
        );

    \I__6269\ : InMux
    port map (
            O => \N__32426\,
            I => \N__32420\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__32423\,
            I => \N__32417\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__32420\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__6266\ : Odrv12
    port map (
            O => \N__32417\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__6265\ : CEMux
    port map (
            O => \N__32412\,
            I => \N__32408\
        );

    \I__6264\ : CEMux
    port map (
            O => \N__32411\,
            I => \N__32405\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__32408\,
            I => \N__32398\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__32405\,
            I => \N__32398\
        );

    \I__6261\ : CEMux
    port map (
            O => \N__32404\,
            I => \N__32395\
        );

    \I__6260\ : CEMux
    port map (
            O => \N__32403\,
            I => \N__32392\
        );

    \I__6259\ : Span4Mux_v
    port map (
            O => \N__32398\,
            I => \N__32389\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__32395\,
            I => \N__32384\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__32392\,
            I => \N__32384\
        );

    \I__6256\ : Span4Mux_h
    port map (
            O => \N__32389\,
            I => \N__32379\
        );

    \I__6255\ : Span4Mux_v
    port map (
            O => \N__32384\,
            I => \N__32379\
        );

    \I__6254\ : Span4Mux_v
    port map (
            O => \N__32379\,
            I => \N__32376\
        );

    \I__6253\ : Odrv4
    port map (
            O => \N__32376\,
            I => \current_shift_inst.timer_s1.N_191_i\
        );

    \I__6252\ : IoInMux
    port map (
            O => \N__32373\,
            I => \N__32370\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__32370\,
            I => \N__32367\
        );

    \I__6250\ : Span4Mux_s0_v
    port map (
            O => \N__32367\,
            I => \N__32364\
        );

    \I__6249\ : Span4Mux_v
    port map (
            O => \N__32364\,
            I => \N__32361\
        );

    \I__6248\ : Odrv4
    port map (
            O => \N__32361\,
            I => \current_shift_inst.timer_phase.N_188_i\
        );

    \I__6247\ : CascadeMux
    port map (
            O => \N__32358\,
            I => \N__32354\
        );

    \I__6246\ : CascadeMux
    port map (
            O => \N__32357\,
            I => \N__32351\
        );

    \I__6245\ : InMux
    port map (
            O => \N__32354\,
            I => \N__32346\
        );

    \I__6244\ : InMux
    port map (
            O => \N__32351\,
            I => \N__32346\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__32346\,
            I => \N__32342\
        );

    \I__6242\ : InMux
    port map (
            O => \N__32345\,
            I => \N__32339\
        );

    \I__6241\ : Span4Mux_v
    port map (
            O => \N__32342\,
            I => \N__32336\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__32339\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__6239\ : Odrv4
    port map (
            O => \N__32336\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__6238\ : InMux
    port map (
            O => \N__32331\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__6237\ : CascadeMux
    port map (
            O => \N__32328\,
            I => \N__32324\
        );

    \I__6236\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32321\
        );

    \I__6235\ : InMux
    port map (
            O => \N__32324\,
            I => \N__32318\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__32321\,
            I => \N__32312\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__32318\,
            I => \N__32312\
        );

    \I__6232\ : InMux
    port map (
            O => \N__32317\,
            I => \N__32309\
        );

    \I__6231\ : Span4Mux_v
    port map (
            O => \N__32312\,
            I => \N__32306\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__32309\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__6229\ : Odrv4
    port map (
            O => \N__32306\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__6228\ : InMux
    port map (
            O => \N__32301\,
            I => \bfn_12_21_0_\
        );

    \I__6227\ : InMux
    port map (
            O => \N__32298\,
            I => \N__32294\
        );

    \I__6226\ : InMux
    port map (
            O => \N__32297\,
            I => \N__32291\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__32294\,
            I => \N__32285\
        );

    \I__6224\ : LocalMux
    port map (
            O => \N__32291\,
            I => \N__32285\
        );

    \I__6223\ : InMux
    port map (
            O => \N__32290\,
            I => \N__32282\
        );

    \I__6222\ : Span4Mux_v
    port map (
            O => \N__32285\,
            I => \N__32279\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__32282\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__6220\ : Odrv4
    port map (
            O => \N__32279\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__6219\ : InMux
    port map (
            O => \N__32274\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__6218\ : CascadeMux
    port map (
            O => \N__32271\,
            I => \N__32267\
        );

    \I__6217\ : CascadeMux
    port map (
            O => \N__32270\,
            I => \N__32264\
        );

    \I__6216\ : InMux
    port map (
            O => \N__32267\,
            I => \N__32259\
        );

    \I__6215\ : InMux
    port map (
            O => \N__32264\,
            I => \N__32259\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__32259\,
            I => \N__32255\
        );

    \I__6213\ : InMux
    port map (
            O => \N__32258\,
            I => \N__32252\
        );

    \I__6212\ : Span4Mux_v
    port map (
            O => \N__32255\,
            I => \N__32249\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__32252\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__6210\ : Odrv4
    port map (
            O => \N__32249\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__6209\ : InMux
    port map (
            O => \N__32244\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__6208\ : CascadeMux
    port map (
            O => \N__32241\,
            I => \N__32237\
        );

    \I__6207\ : CascadeMux
    port map (
            O => \N__32240\,
            I => \N__32234\
        );

    \I__6206\ : InMux
    port map (
            O => \N__32237\,
            I => \N__32229\
        );

    \I__6205\ : InMux
    port map (
            O => \N__32234\,
            I => \N__32229\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__32229\,
            I => \N__32225\
        );

    \I__6203\ : InMux
    port map (
            O => \N__32228\,
            I => \N__32222\
        );

    \I__6202\ : Span4Mux_v
    port map (
            O => \N__32225\,
            I => \N__32219\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__32222\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__6200\ : Odrv4
    port map (
            O => \N__32219\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__6199\ : InMux
    port map (
            O => \N__32214\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__6198\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32205\
        );

    \I__6197\ : InMux
    port map (
            O => \N__32210\,
            I => \N__32205\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__32205\,
            I => \N__32201\
        );

    \I__6195\ : InMux
    port map (
            O => \N__32204\,
            I => \N__32198\
        );

    \I__6194\ : Span4Mux_v
    port map (
            O => \N__32201\,
            I => \N__32195\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__32198\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__6192\ : Odrv4
    port map (
            O => \N__32195\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__6191\ : InMux
    port map (
            O => \N__32190\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__6190\ : InMux
    port map (
            O => \N__32187\,
            I => \N__32180\
        );

    \I__6189\ : InMux
    port map (
            O => \N__32186\,
            I => \N__32180\
        );

    \I__6188\ : InMux
    port map (
            O => \N__32185\,
            I => \N__32177\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__32180\,
            I => \N__32174\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__32177\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__6185\ : Odrv12
    port map (
            O => \N__32174\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__6184\ : InMux
    port map (
            O => \N__32169\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__6183\ : CascadeMux
    port map (
            O => \N__32166\,
            I => \N__32162\
        );

    \I__6182\ : CascadeMux
    port map (
            O => \N__32165\,
            I => \N__32159\
        );

    \I__6181\ : InMux
    port map (
            O => \N__32162\,
            I => \N__32153\
        );

    \I__6180\ : InMux
    port map (
            O => \N__32159\,
            I => \N__32153\
        );

    \I__6179\ : InMux
    port map (
            O => \N__32158\,
            I => \N__32150\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__32153\,
            I => \N__32147\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__32150\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__6176\ : Odrv12
    port map (
            O => \N__32147\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__6175\ : InMux
    port map (
            O => \N__32142\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__6174\ : CascadeMux
    port map (
            O => \N__32139\,
            I => \N__32135\
        );

    \I__6173\ : CascadeMux
    port map (
            O => \N__32138\,
            I => \N__32132\
        );

    \I__6172\ : InMux
    port map (
            O => \N__32135\,
            I => \N__32126\
        );

    \I__6171\ : InMux
    port map (
            O => \N__32132\,
            I => \N__32126\
        );

    \I__6170\ : InMux
    port map (
            O => \N__32131\,
            I => \N__32123\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__32126\,
            I => \N__32120\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__32123\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__6167\ : Odrv12
    port map (
            O => \N__32120\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__6166\ : InMux
    port map (
            O => \N__32115\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__6165\ : CascadeMux
    port map (
            O => \N__32112\,
            I => \N__32108\
        );

    \I__6164\ : CascadeMux
    port map (
            O => \N__32111\,
            I => \N__32105\
        );

    \I__6163\ : InMux
    port map (
            O => \N__32108\,
            I => \N__32100\
        );

    \I__6162\ : InMux
    port map (
            O => \N__32105\,
            I => \N__32100\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__32100\,
            I => \N__32096\
        );

    \I__6160\ : InMux
    port map (
            O => \N__32099\,
            I => \N__32093\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__32096\,
            I => \N__32090\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__32093\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__6157\ : Odrv4
    port map (
            O => \N__32090\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__6156\ : InMux
    port map (
            O => \N__32085\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__6155\ : InMux
    port map (
            O => \N__32082\,
            I => \N__32078\
        );

    \I__6154\ : InMux
    port map (
            O => \N__32081\,
            I => \N__32075\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__32078\,
            I => \N__32069\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__32075\,
            I => \N__32069\
        );

    \I__6151\ : InMux
    port map (
            O => \N__32074\,
            I => \N__32066\
        );

    \I__6150\ : Span4Mux_v
    port map (
            O => \N__32069\,
            I => \N__32063\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__32066\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__6148\ : Odrv4
    port map (
            O => \N__32063\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__6147\ : InMux
    port map (
            O => \N__32058\,
            I => \bfn_12_20_0_\
        );

    \I__6146\ : InMux
    port map (
            O => \N__32055\,
            I => \N__32050\
        );

    \I__6145\ : InMux
    port map (
            O => \N__32054\,
            I => \N__32047\
        );

    \I__6144\ : InMux
    port map (
            O => \N__32053\,
            I => \N__32044\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__32050\,
            I => \N__32039\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__32047\,
            I => \N__32039\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__32044\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__6140\ : Odrv12
    port map (
            O => \N__32039\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__6139\ : InMux
    port map (
            O => \N__32034\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__6138\ : CascadeMux
    port map (
            O => \N__32031\,
            I => \N__32027\
        );

    \I__6137\ : CascadeMux
    port map (
            O => \N__32030\,
            I => \N__32024\
        );

    \I__6136\ : InMux
    port map (
            O => \N__32027\,
            I => \N__32018\
        );

    \I__6135\ : InMux
    port map (
            O => \N__32024\,
            I => \N__32018\
        );

    \I__6134\ : InMux
    port map (
            O => \N__32023\,
            I => \N__32015\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__32018\,
            I => \N__32012\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__32015\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__6131\ : Odrv12
    port map (
            O => \N__32012\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__6130\ : InMux
    port map (
            O => \N__32007\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__6129\ : CascadeMux
    port map (
            O => \N__32004\,
            I => \N__32000\
        );

    \I__6128\ : CascadeMux
    port map (
            O => \N__32003\,
            I => \N__31997\
        );

    \I__6127\ : InMux
    port map (
            O => \N__32000\,
            I => \N__31991\
        );

    \I__6126\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31991\
        );

    \I__6125\ : InMux
    port map (
            O => \N__31996\,
            I => \N__31988\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__31991\,
            I => \N__31985\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__31988\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__6122\ : Odrv12
    port map (
            O => \N__31985\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__6121\ : InMux
    port map (
            O => \N__31980\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__6120\ : InMux
    port map (
            O => \N__31977\,
            I => \N__31970\
        );

    \I__6119\ : InMux
    port map (
            O => \N__31976\,
            I => \N__31970\
        );

    \I__6118\ : InMux
    port map (
            O => \N__31975\,
            I => \N__31967\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__31970\,
            I => \N__31964\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__31967\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__6115\ : Odrv12
    port map (
            O => \N__31964\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__6114\ : InMux
    port map (
            O => \N__31959\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__6113\ : InMux
    port map (
            O => \N__31956\,
            I => \N__31950\
        );

    \I__6112\ : InMux
    port map (
            O => \N__31955\,
            I => \N__31950\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__31950\,
            I => \N__31946\
        );

    \I__6110\ : InMux
    port map (
            O => \N__31949\,
            I => \N__31943\
        );

    \I__6109\ : Span4Mux_v
    port map (
            O => \N__31946\,
            I => \N__31940\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__31943\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__6107\ : Odrv4
    port map (
            O => \N__31940\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__6106\ : InMux
    port map (
            O => \N__31935\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__6105\ : CascadeMux
    port map (
            O => \N__31932\,
            I => \N__31929\
        );

    \I__6104\ : InMux
    port map (
            O => \N__31929\,
            I => \N__31925\
        );

    \I__6103\ : InMux
    port map (
            O => \N__31928\,
            I => \N__31921\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__31925\,
            I => \N__31918\
        );

    \I__6101\ : InMux
    port map (
            O => \N__31924\,
            I => \N__31915\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__31921\,
            I => \N__31912\
        );

    \I__6099\ : Span4Mux_v
    port map (
            O => \N__31918\,
            I => \N__31909\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__31915\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__6097\ : Odrv12
    port map (
            O => \N__31912\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__6096\ : Odrv4
    port map (
            O => \N__31909\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__6095\ : InMux
    port map (
            O => \N__31902\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__6094\ : InMux
    port map (
            O => \N__31899\,
            I => \N__31896\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__31896\,
            I => \N__31893\
        );

    \I__6092\ : Odrv4
    port map (
            O => \N__31893\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_25\
        );

    \I__6091\ : InMux
    port map (
            O => \N__31890\,
            I => \N__31887\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__31887\,
            I => \current_shift_inst.un4_control_input_axb_25\
        );

    \I__6089\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31881\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__31881\,
            I => \N__31878\
        );

    \I__6087\ : Odrv4
    port map (
            O => \N__31878\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_22\
        );

    \I__6086\ : InMux
    port map (
            O => \N__31875\,
            I => \N__31872\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__31872\,
            I => \current_shift_inst.un4_control_input_axb_22\
        );

    \I__6084\ : InMux
    port map (
            O => \N__31869\,
            I => \N__31865\
        );

    \I__6083\ : CascadeMux
    port map (
            O => \N__31868\,
            I => \N__31862\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__31865\,
            I => \N__31859\
        );

    \I__6081\ : InMux
    port map (
            O => \N__31862\,
            I => \N__31855\
        );

    \I__6080\ : Span4Mux_h
    port map (
            O => \N__31859\,
            I => \N__31852\
        );

    \I__6079\ : InMux
    port map (
            O => \N__31858\,
            I => \N__31849\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__31855\,
            I => \N__31846\
        );

    \I__6077\ : Odrv4
    port map (
            O => \N__31852\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__31849\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__6075\ : Odrv12
    port map (
            O => \N__31846\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__6074\ : InMux
    port map (
            O => \N__31839\,
            I => \bfn_12_19_0_\
        );

    \I__6073\ : InMux
    port map (
            O => \N__31836\,
            I => \N__31832\
        );

    \I__6072\ : CascadeMux
    port map (
            O => \N__31835\,
            I => \N__31829\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__31832\,
            I => \N__31826\
        );

    \I__6070\ : InMux
    port map (
            O => \N__31829\,
            I => \N__31822\
        );

    \I__6069\ : Span4Mux_h
    port map (
            O => \N__31826\,
            I => \N__31819\
        );

    \I__6068\ : InMux
    port map (
            O => \N__31825\,
            I => \N__31816\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__31822\,
            I => \N__31813\
        );

    \I__6066\ : Odrv4
    port map (
            O => \N__31819\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__31816\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__6064\ : Odrv12
    port map (
            O => \N__31813\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__6063\ : InMux
    port map (
            O => \N__31806\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__6062\ : InMux
    port map (
            O => \N__31803\,
            I => \N__31796\
        );

    \I__6061\ : InMux
    port map (
            O => \N__31802\,
            I => \N__31796\
        );

    \I__6060\ : InMux
    port map (
            O => \N__31801\,
            I => \N__31793\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__31796\,
            I => \N__31790\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__31793\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__6057\ : Odrv12
    port map (
            O => \N__31790\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__6056\ : InMux
    port map (
            O => \N__31785\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__6055\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31775\
        );

    \I__6054\ : InMux
    port map (
            O => \N__31781\,
            I => \N__31775\
        );

    \I__6053\ : InMux
    port map (
            O => \N__31780\,
            I => \N__31772\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__31775\,
            I => \N__31769\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__31772\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__6050\ : Odrv12
    port map (
            O => \N__31769\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__6049\ : InMux
    port map (
            O => \N__31764\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__6048\ : CascadeMux
    port map (
            O => \N__31761\,
            I => \N__31758\
        );

    \I__6047\ : InMux
    port map (
            O => \N__31758\,
            I => \N__31754\
        );

    \I__6046\ : InMux
    port map (
            O => \N__31757\,
            I => \N__31750\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__31754\,
            I => \N__31747\
        );

    \I__6044\ : InMux
    port map (
            O => \N__31753\,
            I => \N__31744\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__31750\,
            I => \N__31739\
        );

    \I__6042\ : Sp12to4
    port map (
            O => \N__31747\,
            I => \N__31739\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__31744\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__6040\ : Odrv12
    port map (
            O => \N__31739\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__6039\ : InMux
    port map (
            O => \N__31734\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__6038\ : CascadeMux
    port map (
            O => \N__31731\,
            I => \N__31728\
        );

    \I__6037\ : InMux
    port map (
            O => \N__31728\,
            I => \N__31724\
        );

    \I__6036\ : InMux
    port map (
            O => \N__31727\,
            I => \N__31720\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__31724\,
            I => \N__31717\
        );

    \I__6034\ : InMux
    port map (
            O => \N__31723\,
            I => \N__31714\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__31720\,
            I => \N__31709\
        );

    \I__6032\ : Sp12to4
    port map (
            O => \N__31717\,
            I => \N__31709\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__31714\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__6030\ : Odrv12
    port map (
            O => \N__31709\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__6029\ : InMux
    port map (
            O => \N__31704\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__6028\ : InMux
    port map (
            O => \N__31701\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__6027\ : CEMux
    port map (
            O => \N__31698\,
            I => \N__31683\
        );

    \I__6026\ : CEMux
    port map (
            O => \N__31697\,
            I => \N__31683\
        );

    \I__6025\ : CEMux
    port map (
            O => \N__31696\,
            I => \N__31683\
        );

    \I__6024\ : CEMux
    port map (
            O => \N__31695\,
            I => \N__31683\
        );

    \I__6023\ : CEMux
    port map (
            O => \N__31694\,
            I => \N__31683\
        );

    \I__6022\ : GlobalMux
    port map (
            O => \N__31683\,
            I => \N__31680\
        );

    \I__6021\ : gio2CtrlBuf
    port map (
            O => \N__31680\,
            I => \current_shift_inst.timer_s1.N_187_i_g\
        );

    \I__6020\ : InMux
    port map (
            O => \N__31677\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__6019\ : InMux
    port map (
            O => \N__31674\,
            I => \N__31668\
        );

    \I__6018\ : InMux
    port map (
            O => \N__31673\,
            I => \N__31668\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__31668\,
            I => \N__31665\
        );

    \I__6016\ : Span4Mux_h
    port map (
            O => \N__31665\,
            I => \N__31662\
        );

    \I__6015\ : Odrv4
    port map (
            O => \N__31662\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__6014\ : InMux
    port map (
            O => \N__31659\,
            I => \N__31656\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__31656\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_29\
        );

    \I__6012\ : InMux
    port map (
            O => \N__31653\,
            I => \N__31650\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__31650\,
            I => \N__31647\
        );

    \I__6010\ : Odrv4
    port map (
            O => \N__31647\,
            I => \current_shift_inst.un4_control_input_axb_29\
        );

    \I__6009\ : InMux
    port map (
            O => \N__31644\,
            I => \N__31641\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__31641\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_28\
        );

    \I__6007\ : InMux
    port map (
            O => \N__31638\,
            I => \N__31635\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__31635\,
            I => \current_shift_inst.un4_control_input_axb_28\
        );

    \I__6005\ : InMux
    port map (
            O => \N__31632\,
            I => \N__31629\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__31629\,
            I => \N__31626\
        );

    \I__6003\ : Odrv4
    port map (
            O => \N__31626\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_20\
        );

    \I__6002\ : InMux
    port map (
            O => \N__31623\,
            I => \N__31620\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__31620\,
            I => \current_shift_inst.un4_control_input_axb_20\
        );

    \I__6000\ : InMux
    port map (
            O => \N__31617\,
            I => \N__31614\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__31614\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_30\
        );

    \I__5998\ : CascadeMux
    port map (
            O => \N__31611\,
            I => \N__31608\
        );

    \I__5997\ : InMux
    port map (
            O => \N__31608\,
            I => \N__31605\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__31605\,
            I => \current_shift_inst.un4_control_input_axb_30\
        );

    \I__5995\ : InMux
    port map (
            O => \N__31602\,
            I => \N__31599\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__31599\,
            I => \N__31596\
        );

    \I__5993\ : Odrv4
    port map (
            O => \N__31596\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_19\
        );

    \I__5992\ : CascadeMux
    port map (
            O => \N__31593\,
            I => \N__31590\
        );

    \I__5991\ : InMux
    port map (
            O => \N__31590\,
            I => \N__31587\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__31587\,
            I => \current_shift_inst.un4_control_input_axb_19\
        );

    \I__5989\ : InMux
    port map (
            O => \N__31584\,
            I => \N__31581\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__31581\,
            I => \N__31578\
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__31578\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_26\
        );

    \I__5986\ : InMux
    port map (
            O => \N__31575\,
            I => \N__31572\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__31572\,
            I => \current_shift_inst.un4_control_input_axb_26\
        );

    \I__5984\ : InMux
    port map (
            O => \N__31569\,
            I => \N__31566\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__31566\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_27\
        );

    \I__5982\ : InMux
    port map (
            O => \N__31563\,
            I => \N__31560\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__31560\,
            I => \current_shift_inst.un4_control_input_axb_27\
        );

    \I__5980\ : InMux
    port map (
            O => \N__31557\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__5979\ : InMux
    port map (
            O => \N__31554\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__5978\ : InMux
    port map (
            O => \N__31551\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__5977\ : InMux
    port map (
            O => \N__31548\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__5976\ : InMux
    port map (
            O => \N__31545\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__5975\ : InMux
    port map (
            O => \N__31542\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__5974\ : InMux
    port map (
            O => \N__31539\,
            I => \bfn_12_17_0_\
        );

    \I__5973\ : InMux
    port map (
            O => \N__31536\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__5972\ : InMux
    port map (
            O => \N__31533\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__5971\ : InMux
    port map (
            O => \N__31530\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__5970\ : InMux
    port map (
            O => \N__31527\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__5969\ : InMux
    port map (
            O => \N__31524\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__5968\ : InMux
    port map (
            O => \N__31521\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__5967\ : InMux
    port map (
            O => \N__31518\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__5966\ : InMux
    port map (
            O => \N__31515\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__5965\ : InMux
    port map (
            O => \N__31512\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__5964\ : InMux
    port map (
            O => \N__31509\,
            I => \bfn_12_16_0_\
        );

    \I__5963\ : InMux
    port map (
            O => \N__31506\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__5962\ : InMux
    port map (
            O => \N__31503\,
            I => \N__31500\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__31500\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_4\
        );

    \I__5960\ : InMux
    port map (
            O => \N__31497\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__5959\ : InMux
    port map (
            O => \N__31494\,
            I => \N__31491\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__31491\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_5\
        );

    \I__5957\ : InMux
    port map (
            O => \N__31488\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__5956\ : InMux
    port map (
            O => \N__31485\,
            I => \N__31482\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__31482\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_6\
        );

    \I__5954\ : InMux
    port map (
            O => \N__31479\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__5953\ : InMux
    port map (
            O => \N__31476\,
            I => \N__31473\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__31473\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_7\
        );

    \I__5951\ : InMux
    port map (
            O => \N__31470\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__5950\ : InMux
    port map (
            O => \N__31467\,
            I => \N__31464\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__31464\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_8\
        );

    \I__5948\ : InMux
    port map (
            O => \N__31461\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__5947\ : InMux
    port map (
            O => \N__31458\,
            I => \N__31455\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__31455\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_9\
        );

    \I__5945\ : InMux
    port map (
            O => \N__31452\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__5944\ : InMux
    port map (
            O => \N__31449\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__5943\ : InMux
    port map (
            O => \N__31446\,
            I => \bfn_12_15_0_\
        );

    \I__5942\ : InMux
    port map (
            O => \N__31443\,
            I => \N__31439\
        );

    \I__5941\ : InMux
    port map (
            O => \N__31442\,
            I => \N__31436\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__31439\,
            I => \N__31433\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__31436\,
            I => \N__31430\
        );

    \I__5938\ : Odrv4
    port map (
            O => \N__31433\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt15\
        );

    \I__5937\ : Odrv12
    port map (
            O => \N__31430\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt15\
        );

    \I__5936\ : InMux
    port map (
            O => \N__31425\,
            I => \N__31422\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__31422\,
            I => \N__31417\
        );

    \I__5934\ : CascadeMux
    port map (
            O => \N__31421\,
            I => \N__31414\
        );

    \I__5933\ : CascadeMux
    port map (
            O => \N__31420\,
            I => \N__31411\
        );

    \I__5932\ : Span4Mux_v
    port map (
            O => \N__31417\,
            I => \N__31408\
        );

    \I__5931\ : InMux
    port map (
            O => \N__31414\,
            I => \N__31405\
        );

    \I__5930\ : InMux
    port map (
            O => \N__31411\,
            I => \N__31402\
        );

    \I__5929\ : Odrv4
    port map (
            O => \N__31408\,
            I => \current_shift_inst.S3_riseZ0\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__31405\,
            I => \current_shift_inst.S3_riseZ0\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__31402\,
            I => \current_shift_inst.S3_riseZ0\
        );

    \I__5926\ : InMux
    port map (
            O => \N__31395\,
            I => \N__31389\
        );

    \I__5925\ : InMux
    port map (
            O => \N__31394\,
            I => \N__31386\
        );

    \I__5924\ : InMux
    port map (
            O => \N__31393\,
            I => \N__31381\
        );

    \I__5923\ : InMux
    port map (
            O => \N__31392\,
            I => \N__31381\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__31389\,
            I => \N__31374\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__31386\,
            I => \N__31374\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__31381\,
            I => \N__31374\
        );

    \I__5919\ : Span4Mux_h
    port map (
            O => \N__31374\,
            I => \N__31368\
        );

    \I__5918\ : InMux
    port map (
            O => \N__31373\,
            I => \N__31363\
        );

    \I__5917\ : InMux
    port map (
            O => \N__31372\,
            I => \N__31363\
        );

    \I__5916\ : InMux
    port map (
            O => \N__31371\,
            I => \N__31360\
        );

    \I__5915\ : Odrv4
    port map (
            O => \N__31368\,
            I => \current_shift_inst.S1_riseZ0\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__31363\,
            I => \current_shift_inst.S1_riseZ0\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__31360\,
            I => \current_shift_inst.S1_riseZ0\
        );

    \I__5912\ : InMux
    port map (
            O => \N__31353\,
            I => \N__31350\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__31350\,
            I => \N__31347\
        );

    \I__5910\ : Odrv4
    port map (
            O => \N__31347\,
            I => \current_shift_inst.N_199\
        );

    \I__5909\ : CascadeMux
    port map (
            O => \N__31344\,
            I => \N__31339\
        );

    \I__5908\ : CascadeMux
    port map (
            O => \N__31343\,
            I => \N__31336\
        );

    \I__5907\ : InMux
    port map (
            O => \N__31342\,
            I => \N__31328\
        );

    \I__5906\ : InMux
    port map (
            O => \N__31339\,
            I => \N__31328\
        );

    \I__5905\ : InMux
    port map (
            O => \N__31336\,
            I => \N__31323\
        );

    \I__5904\ : InMux
    port map (
            O => \N__31335\,
            I => \N__31323\
        );

    \I__5903\ : InMux
    port map (
            O => \N__31334\,
            I => \N__31317\
        );

    \I__5902\ : InMux
    port map (
            O => \N__31333\,
            I => \N__31317\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__31328\,
            I => \N__31312\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__31323\,
            I => \N__31312\
        );

    \I__5899\ : InMux
    port map (
            O => \N__31322\,
            I => \N__31309\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__31317\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__5897\ : Odrv4
    port map (
            O => \N__31312\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__31309\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__5895\ : InMux
    port map (
            O => \N__31302\,
            I => \N__31298\
        );

    \I__5894\ : InMux
    port map (
            O => \N__31301\,
            I => \N__31295\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__31298\,
            I => measured_delay_hc_28
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__31295\,
            I => measured_delay_hc_28
        );

    \I__5891\ : CascadeMux
    port map (
            O => \N__31290\,
            I => \N__31287\
        );

    \I__5890\ : InMux
    port map (
            O => \N__31287\,
            I => \N__31283\
        );

    \I__5889\ : InMux
    port map (
            O => \N__31286\,
            I => \N__31280\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__31283\,
            I => measured_delay_hc_29
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__31280\,
            I => measured_delay_hc_29
        );

    \I__5886\ : CascadeMux
    port map (
            O => \N__31275\,
            I => \N__31271\
        );

    \I__5885\ : InMux
    port map (
            O => \N__31274\,
            I => \N__31268\
        );

    \I__5884\ : InMux
    port map (
            O => \N__31271\,
            I => \N__31265\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__31268\,
            I => measured_delay_hc_30
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__31265\,
            I => measured_delay_hc_30
        );

    \I__5881\ : InMux
    port map (
            O => \N__31260\,
            I => \N__31257\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__31257\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_3\
        );

    \I__5879\ : CascadeMux
    port map (
            O => \N__31254\,
            I => \N__31251\
        );

    \I__5878\ : InMux
    port map (
            O => \N__31251\,
            I => \N__31248\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__31248\,
            I => \N__31245\
        );

    \I__5876\ : Odrv12
    port map (
            O => \N__31245\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__5875\ : InMux
    port map (
            O => \N__31242\,
            I => \N__31239\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__31239\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\
        );

    \I__5873\ : CascadeMux
    port map (
            O => \N__31236\,
            I => \N__31233\
        );

    \I__5872\ : InMux
    port map (
            O => \N__31233\,
            I => \N__31230\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__31230\,
            I => \N__31227\
        );

    \I__5870\ : Span4Mux_v
    port map (
            O => \N__31227\,
            I => \N__31224\
        );

    \I__5869\ : Odrv4
    port map (
            O => \N__31224\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__5868\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31218\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__31218\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\
        );

    \I__5866\ : InMux
    port map (
            O => \N__31215\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__5865\ : InMux
    port map (
            O => \N__31212\,
            I => \N__31209\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__31209\,
            I => \N__31206\
        );

    \I__5863\ : Odrv4
    port map (
            O => \N__31206\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10\
        );

    \I__5862\ : InMux
    port map (
            O => \N__31203\,
            I => \N__31200\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__31200\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\
        );

    \I__5860\ : InMux
    port map (
            O => \N__31197\,
            I => \N__31194\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__31194\,
            I => \current_shift_inst.S3_sync_prevZ0\
        );

    \I__5858\ : InMux
    port map (
            O => \N__31191\,
            I => \N__31187\
        );

    \I__5857\ : CascadeMux
    port map (
            O => \N__31190\,
            I => \N__31184\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__31187\,
            I => \N__31181\
        );

    \I__5855\ : InMux
    port map (
            O => \N__31184\,
            I => \N__31178\
        );

    \I__5854\ : Odrv4
    port map (
            O => \N__31181\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__31178\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\
        );

    \I__5852\ : CascadeMux
    port map (
            O => \N__31173\,
            I => \N__31170\
        );

    \I__5851\ : InMux
    port map (
            O => \N__31170\,
            I => \N__31167\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__31167\,
            I => \N__31164\
        );

    \I__5849\ : Odrv4
    port map (
            O => \N__31164\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__5848\ : InMux
    port map (
            O => \N__31161\,
            I => \N__31158\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__31158\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__5846\ : CascadeMux
    port map (
            O => \N__31155\,
            I => \N__31152\
        );

    \I__5845\ : InMux
    port map (
            O => \N__31152\,
            I => \N__31149\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__31149\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__5843\ : InMux
    port map (
            O => \N__31146\,
            I => \N__31143\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__31143\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__5841\ : CascadeMux
    port map (
            O => \N__31140\,
            I => \N__31137\
        );

    \I__5840\ : InMux
    port map (
            O => \N__31137\,
            I => \N__31134\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__31134\,
            I => \N__31131\
        );

    \I__5838\ : Odrv4
    port map (
            O => \N__31131\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__5837\ : InMux
    port map (
            O => \N__31128\,
            I => \N__31125\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__31125\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__5835\ : CascadeMux
    port map (
            O => \N__31122\,
            I => \N__31119\
        );

    \I__5834\ : InMux
    port map (
            O => \N__31119\,
            I => \N__31116\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__31116\,
            I => \N__31113\
        );

    \I__5832\ : Span4Mux_h
    port map (
            O => \N__31113\,
            I => \N__31110\
        );

    \I__5831\ : Odrv4
    port map (
            O => \N__31110\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__5830\ : InMux
    port map (
            O => \N__31107\,
            I => \N__31104\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__31104\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__5828\ : CascadeMux
    port map (
            O => \N__31101\,
            I => \N__31098\
        );

    \I__5827\ : InMux
    port map (
            O => \N__31098\,
            I => \N__31095\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__31095\,
            I => \N__31092\
        );

    \I__5825\ : Odrv4
    port map (
            O => \N__31092\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__5824\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31086\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__31086\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__31083\,
            I => \N__31080\
        );

    \I__5821\ : InMux
    port map (
            O => \N__31080\,
            I => \N__31077\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__31077\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__5819\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31071\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__31071\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\
        );

    \I__5817\ : CascadeMux
    port map (
            O => \N__31068\,
            I => \N__31065\
        );

    \I__5816\ : InMux
    port map (
            O => \N__31065\,
            I => \N__31062\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__31062\,
            I => \N__31059\
        );

    \I__5814\ : Odrv4
    port map (
            O => \N__31059\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__5813\ : InMux
    port map (
            O => \N__31056\,
            I => \N__31053\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__31053\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\
        );

    \I__5811\ : CascadeMux
    port map (
            O => \N__31050\,
            I => \N__31047\
        );

    \I__5810\ : InMux
    port map (
            O => \N__31047\,
            I => \N__31044\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__31044\,
            I => \N__31041\
        );

    \I__5808\ : Odrv4
    port map (
            O => \N__31041\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__5807\ : InMux
    port map (
            O => \N__31038\,
            I => \N__31035\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__31035\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__31032\,
            I => \N__31029\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31029\,
            I => \N__31026\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__31026\,
            I => \N__31023\
        );

    \I__5802\ : Odrv4
    port map (
            O => \N__31023\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__5801\ : InMux
    port map (
            O => \N__31020\,
            I => \N__31017\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__31017\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__5799\ : CascadeMux
    port map (
            O => \N__31014\,
            I => \N__31011\
        );

    \I__5798\ : InMux
    port map (
            O => \N__31011\,
            I => \N__31008\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__31008\,
            I => \N__31005\
        );

    \I__5796\ : Span4Mux_h
    port map (
            O => \N__31005\,
            I => \N__31002\
        );

    \I__5795\ : Odrv4
    port map (
            O => \N__31002\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__5794\ : InMux
    port map (
            O => \N__30999\,
            I => \N__30996\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__30996\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__5792\ : CascadeMux
    port map (
            O => \N__30993\,
            I => \N__30990\
        );

    \I__5791\ : InMux
    port map (
            O => \N__30990\,
            I => \N__30987\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__30987\,
            I => \N__30984\
        );

    \I__5789\ : Span4Mux_v
    port map (
            O => \N__30984\,
            I => \N__30981\
        );

    \I__5788\ : Odrv4
    port map (
            O => \N__30981\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\
        );

    \I__5787\ : InMux
    port map (
            O => \N__30978\,
            I => \N__30975\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__30975\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__5785\ : CascadeMux
    port map (
            O => \N__30972\,
            I => \N__30969\
        );

    \I__5784\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30966\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__30966\,
            I => \N__30963\
        );

    \I__5782\ : Odrv4
    port map (
            O => \N__30963\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__5781\ : InMux
    port map (
            O => \N__30960\,
            I => \N__30957\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__30957\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__30954\,
            I => \N__30951\
        );

    \I__5778\ : InMux
    port map (
            O => \N__30951\,
            I => \N__30948\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__30948\,
            I => \N__30945\
        );

    \I__5776\ : Span4Mux_v
    port map (
            O => \N__30945\,
            I => \N__30942\
        );

    \I__5775\ : Odrv4
    port map (
            O => \N__30942\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__5774\ : InMux
    port map (
            O => \N__30939\,
            I => \N__30936\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__30936\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__5772\ : CascadeMux
    port map (
            O => \N__30933\,
            I => \N__30930\
        );

    \I__5771\ : InMux
    port map (
            O => \N__30930\,
            I => \N__30927\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__30927\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__5769\ : InMux
    port map (
            O => \N__30924\,
            I => \N__30921\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__30921\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__5767\ : CascadeMux
    port map (
            O => \N__30918\,
            I => \N__30915\
        );

    \I__5766\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30912\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__30912\,
            I => \N__30909\
        );

    \I__5764\ : Odrv4
    port map (
            O => \N__30909\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__5763\ : InMux
    port map (
            O => \N__30906\,
            I => \N__30903\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__30903\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__5761\ : InMux
    port map (
            O => \N__30900\,
            I => \N__30897\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__30897\,
            I => \N__30894\
        );

    \I__5759\ : Odrv12
    port map (
            O => \N__30894\,
            I => \il_max_comp1_D1\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__30891\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto9_cZ0_cascade_\
        );

    \I__5757\ : CEMux
    port map (
            O => \N__30888\,
            I => \N__30878\
        );

    \I__5756\ : CEMux
    port map (
            O => \N__30887\,
            I => \N__30875\
        );

    \I__5755\ : CEMux
    port map (
            O => \N__30886\,
            I => \N__30872\
        );

    \I__5754\ : CEMux
    port map (
            O => \N__30885\,
            I => \N__30869\
        );

    \I__5753\ : CEMux
    port map (
            O => \N__30884\,
            I => \N__30866\
        );

    \I__5752\ : CEMux
    port map (
            O => \N__30883\,
            I => \N__30863\
        );

    \I__5751\ : CEMux
    port map (
            O => \N__30882\,
            I => \N__30860\
        );

    \I__5750\ : CEMux
    port map (
            O => \N__30881\,
            I => \N__30857\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__30878\,
            I => \N__30853\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__30875\,
            I => \N__30850\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__30872\,
            I => \N__30847\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__30869\,
            I => \N__30844\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__30866\,
            I => \N__30841\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__30863\,
            I => \N__30838\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__30860\,
            I => \N__30835\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__30857\,
            I => \N__30832\
        );

    \I__5741\ : CEMux
    port map (
            O => \N__30856\,
            I => \N__30829\
        );

    \I__5740\ : Span12Mux_s10_h
    port map (
            O => \N__30853\,
            I => \N__30826\
        );

    \I__5739\ : Span4Mux_v
    port map (
            O => \N__30850\,
            I => \N__30823\
        );

    \I__5738\ : Span4Mux_v
    port map (
            O => \N__30847\,
            I => \N__30818\
        );

    \I__5737\ : Span4Mux_v
    port map (
            O => \N__30844\,
            I => \N__30818\
        );

    \I__5736\ : Span4Mux_v
    port map (
            O => \N__30841\,
            I => \N__30811\
        );

    \I__5735\ : Span4Mux_h
    port map (
            O => \N__30838\,
            I => \N__30811\
        );

    \I__5734\ : Span4Mux_v
    port map (
            O => \N__30835\,
            I => \N__30811\
        );

    \I__5733\ : Span4Mux_v
    port map (
            O => \N__30832\,
            I => \N__30806\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__30829\,
            I => \N__30806\
        );

    \I__5731\ : Odrv12
    port map (
            O => \N__30826\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5730\ : Odrv4
    port map (
            O => \N__30823\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5729\ : Odrv4
    port map (
            O => \N__30818\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5728\ : Odrv4
    port map (
            O => \N__30811\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5727\ : Odrv4
    port map (
            O => \N__30806\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5726\ : InMux
    port map (
            O => \N__30795\,
            I => \N__30792\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__30792\,
            I => \N__30789\
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__30789\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\
        );

    \I__5723\ : CascadeMux
    port map (
            O => \N__30786\,
            I => \N__30783\
        );

    \I__5722\ : InMux
    port map (
            O => \N__30783\,
            I => \N__30780\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__30780\,
            I => \N__30777\
        );

    \I__5720\ : Odrv4
    port map (
            O => \N__30777\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__5719\ : InMux
    port map (
            O => \N__30774\,
            I => \N__30771\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__30771\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__5717\ : CascadeMux
    port map (
            O => \N__30768\,
            I => \N__30765\
        );

    \I__5716\ : InMux
    port map (
            O => \N__30765\,
            I => \N__30762\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__30762\,
            I => \N__30759\
        );

    \I__5714\ : Span4Mux_v
    port map (
            O => \N__30759\,
            I => \N__30756\
        );

    \I__5713\ : Sp12to4
    port map (
            O => \N__30756\,
            I => \N__30753\
        );

    \I__5712\ : Odrv12
    port map (
            O => \N__30753\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__5711\ : InMux
    port map (
            O => \N__30750\,
            I => \N__30747\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__30747\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__5709\ : CascadeMux
    port map (
            O => \N__30744\,
            I => \N__30741\
        );

    \I__5708\ : InMux
    port map (
            O => \N__30741\,
            I => \N__30738\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__30738\,
            I => \N__30735\
        );

    \I__5706\ : Span4Mux_h
    port map (
            O => \N__30735\,
            I => \N__30732\
        );

    \I__5705\ : Odrv4
    port map (
            O => \N__30732\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24\
        );

    \I__5704\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30726\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__30726\,
            I => \N__30723\
        );

    \I__5702\ : Span4Mux_h
    port map (
            O => \N__30723\,
            I => \N__30719\
        );

    \I__5701\ : InMux
    port map (
            O => \N__30722\,
            I => \N__30716\
        );

    \I__5700\ : Span4Mux_v
    port map (
            O => \N__30719\,
            I => \N__30713\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__30716\,
            I => \current_shift_inst.z_31\
        );

    \I__5698\ : Odrv4
    port map (
            O => \N__30713\,
            I => \current_shift_inst.z_31\
        );

    \I__5697\ : CascadeMux
    port map (
            O => \N__30708\,
            I => \N__30704\
        );

    \I__5696\ : InMux
    port map (
            O => \N__30707\,
            I => \N__30701\
        );

    \I__5695\ : InMux
    port map (
            O => \N__30704\,
            I => \N__30698\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__30701\,
            I => \N__30693\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__30698\,
            I => \N__30693\
        );

    \I__5692\ : Span4Mux_h
    port map (
            O => \N__30693\,
            I => \N__30690\
        );

    \I__5691\ : Span4Mux_v
    port map (
            O => \N__30690\,
            I => \N__30687\
        );

    \I__5690\ : Odrv4
    port map (
            O => \N__30687\,
            I => \current_shift_inst.z_i_31\
        );

    \I__5689\ : CascadeMux
    port map (
            O => \N__30684\,
            I => \N__30680\
        );

    \I__5688\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30676\
        );

    \I__5687\ : InMux
    port map (
            O => \N__30680\,
            I => \N__30671\
        );

    \I__5686\ : InMux
    port map (
            O => \N__30679\,
            I => \N__30671\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__30676\,
            I => \N__30668\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__30671\,
            I => \N__30665\
        );

    \I__5683\ : Span12Mux_s11_v
    port map (
            O => \N__30668\,
            I => \N__30661\
        );

    \I__5682\ : Span4Mux_v
    port map (
            O => \N__30665\,
            I => \N__30658\
        );

    \I__5681\ : InMux
    port map (
            O => \N__30664\,
            I => \N__30655\
        );

    \I__5680\ : Odrv12
    port map (
            O => \N__30661\,
            I => \current_shift_inst.elapsed_time_ns_phase_24\
        );

    \I__5679\ : Odrv4
    port map (
            O => \N__30658\,
            I => \current_shift_inst.elapsed_time_ns_phase_24\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__30655\,
            I => \current_shift_inst.elapsed_time_ns_phase_24\
        );

    \I__5677\ : CascadeMux
    port map (
            O => \N__30648\,
            I => \N__30642\
        );

    \I__5676\ : CascadeMux
    port map (
            O => \N__30647\,
            I => \N__30639\
        );

    \I__5675\ : InMux
    port map (
            O => \N__30646\,
            I => \N__30636\
        );

    \I__5674\ : InMux
    port map (
            O => \N__30645\,
            I => \N__30631\
        );

    \I__5673\ : InMux
    port map (
            O => \N__30642\,
            I => \N__30631\
        );

    \I__5672\ : InMux
    port map (
            O => \N__30639\,
            I => \N__30628\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__30636\,
            I => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__30631\,
            I => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__30628\,
            I => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\
        );

    \I__5668\ : InMux
    port map (
            O => \N__30621\,
            I => \N__30618\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__30618\,
            I => \N__30615\
        );

    \I__5666\ : Span4Mux_h
    port map (
            O => \N__30615\,
            I => \N__30612\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__30612\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23\
        );

    \I__5664\ : CascadeMux
    port map (
            O => \N__30609\,
            I => \N__30606\
        );

    \I__5663\ : InMux
    port map (
            O => \N__30606\,
            I => \N__30603\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__30603\,
            I => \N__30600\
        );

    \I__5661\ : Span4Mux_h
    port map (
            O => \N__30600\,
            I => \N__30597\
        );

    \I__5660\ : Odrv4
    port map (
            O => \N__30597\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIU73K_23\
        );

    \I__5659\ : InMux
    port map (
            O => \N__30594\,
            I => \N__30589\
        );

    \I__5658\ : InMux
    port map (
            O => \N__30593\,
            I => \N__30586\
        );

    \I__5657\ : CascadeMux
    port map (
            O => \N__30592\,
            I => \N__30582\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__30589\,
            I => \N__30574\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__30586\,
            I => \N__30574\
        );

    \I__5654\ : InMux
    port map (
            O => \N__30585\,
            I => \N__30571\
        );

    \I__5653\ : InMux
    port map (
            O => \N__30582\,
            I => \N__30568\
        );

    \I__5652\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30565\
        );

    \I__5651\ : CascadeMux
    port map (
            O => \N__30580\,
            I => \N__30561\
        );

    \I__5650\ : CascadeMux
    port map (
            O => \N__30579\,
            I => \N__30557\
        );

    \I__5649\ : Span4Mux_v
    port map (
            O => \N__30574\,
            I => \N__30552\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__30571\,
            I => \N__30552\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__30568\,
            I => \N__30549\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__30565\,
            I => \N__30546\
        );

    \I__5645\ : InMux
    port map (
            O => \N__30564\,
            I => \N__30537\
        );

    \I__5644\ : InMux
    port map (
            O => \N__30561\,
            I => \N__30537\
        );

    \I__5643\ : InMux
    port map (
            O => \N__30560\,
            I => \N__30537\
        );

    \I__5642\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30537\
        );

    \I__5641\ : Span4Mux_v
    port map (
            O => \N__30552\,
            I => \N__30534\
        );

    \I__5640\ : Odrv4
    port map (
            O => \N__30549\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5639\ : Odrv4
    port map (
            O => \N__30546\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__30537\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5637\ : Odrv4
    port map (
            O => \N__30534\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5636\ : InMux
    port map (
            O => \N__30525\,
            I => \N__30521\
        );

    \I__5635\ : InMux
    port map (
            O => \N__30524\,
            I => \N__30518\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__30521\,
            I => \N__30514\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__30518\,
            I => \N__30511\
        );

    \I__5632\ : InMux
    port map (
            O => \N__30517\,
            I => \N__30508\
        );

    \I__5631\ : Odrv4
    port map (
            O => \N__30514\,
            I => \current_shift_inst.elapsed_time_ns_phase_30\
        );

    \I__5630\ : Odrv4
    port map (
            O => \N__30511\,
            I => \current_shift_inst.elapsed_time_ns_phase_30\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__30508\,
            I => \current_shift_inst.elapsed_time_ns_phase_30\
        );

    \I__5628\ : CascadeMux
    port map (
            O => \N__30501\,
            I => \N__30497\
        );

    \I__5627\ : CascadeMux
    port map (
            O => \N__30500\,
            I => \N__30494\
        );

    \I__5626\ : InMux
    port map (
            O => \N__30497\,
            I => \N__30491\
        );

    \I__5625\ : InMux
    port map (
            O => \N__30494\,
            I => \N__30488\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__30491\,
            I => \N__30483\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__30488\,
            I => \N__30483\
        );

    \I__5622\ : Span4Mux_h
    port map (
            O => \N__30483\,
            I => \N__30480\
        );

    \I__5621\ : Odrv4
    port map (
            O => \N__30480\,
            I => \current_shift_inst.elapsed_time_ns_phase_31\
        );

    \I__5620\ : InMux
    port map (
            O => \N__30477\,
            I => \N__30474\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__30474\,
            I => \N__30470\
        );

    \I__5618\ : InMux
    port map (
            O => \N__30473\,
            I => \N__30466\
        );

    \I__5617\ : Span4Mux_h
    port map (
            O => \N__30470\,
            I => \N__30463\
        );

    \I__5616\ : InMux
    port map (
            O => \N__30469\,
            I => \N__30460\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__30466\,
            I => \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\
        );

    \I__5614\ : Odrv4
    port map (
            O => \N__30463\,
            I => \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__30460\,
            I => \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\
        );

    \I__5612\ : InMux
    port map (
            O => \N__30453\,
            I => \N__30450\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__30450\,
            I => \N__30447\
        );

    \I__5610\ : Span4Mux_v
    port map (
            O => \N__30447\,
            I => \N__30444\
        );

    \I__5609\ : Odrv4
    port map (
            O => \N__30444\,
            I => \current_shift_inst.un38_control_input_0_axb_31\
        );

    \I__5608\ : InMux
    port map (
            O => \N__30441\,
            I => \N__30436\
        );

    \I__5607\ : InMux
    port map (
            O => \N__30440\,
            I => \N__30433\
        );

    \I__5606\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30429\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__30436\,
            I => \N__30426\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__30433\,
            I => \N__30423\
        );

    \I__5603\ : InMux
    port map (
            O => \N__30432\,
            I => \N__30420\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__30429\,
            I => \N__30417\
        );

    \I__5601\ : Span4Mux_h
    port map (
            O => \N__30426\,
            I => \N__30412\
        );

    \I__5600\ : Span4Mux_h
    port map (
            O => \N__30423\,
            I => \N__30412\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__30420\,
            I => \N__30409\
        );

    \I__5598\ : Odrv12
    port map (
            O => \N__30417\,
            I => \current_shift_inst.elapsed_time_ns_phase_26\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__30412\,
            I => \current_shift_inst.elapsed_time_ns_phase_26\
        );

    \I__5596\ : Odrv4
    port map (
            O => \N__30409\,
            I => \current_shift_inst.elapsed_time_ns_phase_26\
        );

    \I__5595\ : InMux
    port map (
            O => \N__30402\,
            I => \N__30399\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__30399\,
            I => \N__30395\
        );

    \I__5593\ : CascadeMux
    port map (
            O => \N__30398\,
            I => \N__30390\
        );

    \I__5592\ : Span4Mux_h
    port map (
            O => \N__30395\,
            I => \N__30387\
        );

    \I__5591\ : InMux
    port map (
            O => \N__30394\,
            I => \N__30384\
        );

    \I__5590\ : InMux
    port map (
            O => \N__30393\,
            I => \N__30381\
        );

    \I__5589\ : InMux
    port map (
            O => \N__30390\,
            I => \N__30378\
        );

    \I__5588\ : Odrv4
    port map (
            O => \N__30387\,
            I => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__30384\,
            I => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__30381\,
            I => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__30378\,
            I => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\
        );

    \I__5584\ : CascadeMux
    port map (
            O => \N__30369\,
            I => \N__30366\
        );

    \I__5583\ : InMux
    port map (
            O => \N__30366\,
            I => \N__30363\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__30363\,
            I => \N__30360\
        );

    \I__5581\ : Span4Mux_h
    port map (
            O => \N__30360\,
            I => \N__30357\
        );

    \I__5580\ : Span4Mux_v
    port map (
            O => \N__30357\,
            I => \N__30354\
        );

    \I__5579\ : Odrv4
    port map (
            O => \N__30354\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26\
        );

    \I__5578\ : CascadeMux
    port map (
            O => \N__30351\,
            I => \N__30347\
        );

    \I__5577\ : InMux
    port map (
            O => \N__30350\,
            I => \N__30343\
        );

    \I__5576\ : InMux
    port map (
            O => \N__30347\,
            I => \N__30338\
        );

    \I__5575\ : InMux
    port map (
            O => \N__30346\,
            I => \N__30338\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__30343\,
            I => \N__30335\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__30338\,
            I => \N__30332\
        );

    \I__5572\ : Span4Mux_v
    port map (
            O => \N__30335\,
            I => \N__30328\
        );

    \I__5571\ : Span4Mux_h
    port map (
            O => \N__30332\,
            I => \N__30325\
        );

    \I__5570\ : InMux
    port map (
            O => \N__30331\,
            I => \N__30322\
        );

    \I__5569\ : Odrv4
    port map (
            O => \N__30328\,
            I => \current_shift_inst.elapsed_time_ns_phase_22\
        );

    \I__5568\ : Odrv4
    port map (
            O => \N__30325\,
            I => \current_shift_inst.elapsed_time_ns_phase_22\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__30322\,
            I => \current_shift_inst.elapsed_time_ns_phase_22\
        );

    \I__5566\ : InMux
    port map (
            O => \N__30315\,
            I => \N__30305\
        );

    \I__5565\ : InMux
    port map (
            O => \N__30314\,
            I => \N__30305\
        );

    \I__5564\ : InMux
    port map (
            O => \N__30313\,
            I => \N__30305\
        );

    \I__5563\ : CascadeMux
    port map (
            O => \N__30312\,
            I => \N__30302\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__30305\,
            I => \N__30299\
        );

    \I__5561\ : InMux
    port map (
            O => \N__30302\,
            I => \N__30296\
        );

    \I__5560\ : Odrv4
    port map (
            O => \N__30299\,
            I => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__30296\,
            I => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\
        );

    \I__5558\ : CascadeMux
    port map (
            O => \N__30291\,
            I => \N__30286\
        );

    \I__5557\ : InMux
    port map (
            O => \N__30290\,
            I => \N__30281\
        );

    \I__5556\ : InMux
    port map (
            O => \N__30289\,
            I => \N__30281\
        );

    \I__5555\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30277\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__30281\,
            I => \N__30274\
        );

    \I__5553\ : CascadeMux
    port map (
            O => \N__30280\,
            I => \N__30271\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__30277\,
            I => \N__30268\
        );

    \I__5551\ : Span4Mux_h
    port map (
            O => \N__30274\,
            I => \N__30265\
        );

    \I__5550\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30262\
        );

    \I__5549\ : Odrv4
    port map (
            O => \N__30268\,
            I => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__30265\,
            I => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__30262\,
            I => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\
        );

    \I__5546\ : CascadeMux
    port map (
            O => \N__30255\,
            I => \N__30251\
        );

    \I__5545\ : InMux
    port map (
            O => \N__30254\,
            I => \N__30243\
        );

    \I__5544\ : InMux
    port map (
            O => \N__30251\,
            I => \N__30243\
        );

    \I__5543\ : InMux
    port map (
            O => \N__30250\,
            I => \N__30243\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__30243\,
            I => \N__30240\
        );

    \I__5541\ : Span4Mux_v
    port map (
            O => \N__30240\,
            I => \N__30236\
        );

    \I__5540\ : InMux
    port map (
            O => \N__30239\,
            I => \N__30233\
        );

    \I__5539\ : Odrv4
    port map (
            O => \N__30236\,
            I => \current_shift_inst.elapsed_time_ns_phase_23\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__30233\,
            I => \current_shift_inst.elapsed_time_ns_phase_23\
        );

    \I__5537\ : InMux
    port map (
            O => \N__30228\,
            I => \N__30225\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__30225\,
            I => \N__30222\
        );

    \I__5535\ : Span4Mux_h
    port map (
            O => \N__30222\,
            I => \N__30219\
        );

    \I__5534\ : Span4Mux_v
    port map (
            O => \N__30219\,
            I => \N__30216\
        );

    \I__5533\ : Odrv4
    port map (
            O => \N__30216\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPB581_22\
        );

    \I__5532\ : InMux
    port map (
            O => \N__30213\,
            I => \bfn_11_19_0_\
        );

    \I__5531\ : InMux
    port map (
            O => \N__30210\,
            I => \current_shift_inst.un4_control_input_cry_25\
        );

    \I__5530\ : InMux
    port map (
            O => \N__30207\,
            I => \current_shift_inst.un4_control_input_cry_26\
        );

    \I__5529\ : CascadeMux
    port map (
            O => \N__30204\,
            I => \N__30200\
        );

    \I__5528\ : CascadeMux
    port map (
            O => \N__30203\,
            I => \N__30197\
        );

    \I__5527\ : InMux
    port map (
            O => \N__30200\,
            I => \N__30189\
        );

    \I__5526\ : InMux
    port map (
            O => \N__30197\,
            I => \N__30189\
        );

    \I__5525\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30189\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__30189\,
            I => \N__30185\
        );

    \I__5523\ : CascadeMux
    port map (
            O => \N__30188\,
            I => \N__30182\
        );

    \I__5522\ : Span4Mux_h
    port map (
            O => \N__30185\,
            I => \N__30179\
        );

    \I__5521\ : InMux
    port map (
            O => \N__30182\,
            I => \N__30176\
        );

    \I__5520\ : Odrv4
    port map (
            O => \N__30179\,
            I => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__30176\,
            I => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\
        );

    \I__5518\ : InMux
    port map (
            O => \N__30171\,
            I => \current_shift_inst.un4_control_input_cry_27\
        );

    \I__5517\ : InMux
    port map (
            O => \N__30168\,
            I => \N__30159\
        );

    \I__5516\ : InMux
    port map (
            O => \N__30167\,
            I => \N__30159\
        );

    \I__5515\ : InMux
    port map (
            O => \N__30166\,
            I => \N__30159\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__30159\,
            I => \N__30155\
        );

    \I__5513\ : CascadeMux
    port map (
            O => \N__30158\,
            I => \N__30152\
        );

    \I__5512\ : Span4Mux_v
    port map (
            O => \N__30155\,
            I => \N__30149\
        );

    \I__5511\ : InMux
    port map (
            O => \N__30152\,
            I => \N__30146\
        );

    \I__5510\ : Odrv4
    port map (
            O => \N__30149\,
            I => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__30146\,
            I => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\
        );

    \I__5508\ : InMux
    port map (
            O => \N__30141\,
            I => \current_shift_inst.un4_control_input_cry_28\
        );

    \I__5507\ : InMux
    port map (
            O => \N__30138\,
            I => \N__30132\
        );

    \I__5506\ : InMux
    port map (
            O => \N__30137\,
            I => \N__30132\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__30132\,
            I => \N__30129\
        );

    \I__5504\ : Span4Mux_v
    port map (
            O => \N__30129\,
            I => \N__30125\
        );

    \I__5503\ : InMux
    port map (
            O => \N__30128\,
            I => \N__30122\
        );

    \I__5502\ : Odrv4
    port map (
            O => \N__30125\,
            I => \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__30122\,
            I => \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\
        );

    \I__5500\ : InMux
    port map (
            O => \N__30117\,
            I => \current_shift_inst.un4_control_input_cry_29\
        );

    \I__5499\ : InMux
    port map (
            O => \N__30114\,
            I => \current_shift_inst.un4_control_input_cry_30\
        );

    \I__5498\ : InMux
    port map (
            O => \N__30111\,
            I => \N__30108\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__30108\,
            I => \N__30105\
        );

    \I__5496\ : Span4Mux_h
    port map (
            O => \N__30105\,
            I => \N__30102\
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__30102\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25\
        );

    \I__5494\ : InMux
    port map (
            O => \N__30099\,
            I => \N__30095\
        );

    \I__5493\ : InMux
    port map (
            O => \N__30098\,
            I => \N__30090\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__30095\,
            I => \N__30087\
        );

    \I__5491\ : InMux
    port map (
            O => \N__30094\,
            I => \N__30084\
        );

    \I__5490\ : InMux
    port map (
            O => \N__30093\,
            I => \N__30081\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__30090\,
            I => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\
        );

    \I__5488\ : Odrv12
    port map (
            O => \N__30087\,
            I => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__30084\,
            I => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__30081\,
            I => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\
        );

    \I__5485\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30067\
        );

    \I__5484\ : CascadeMux
    port map (
            O => \N__30071\,
            I => \N__30064\
        );

    \I__5483\ : InMux
    port map (
            O => \N__30070\,
            I => \N__30061\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__30067\,
            I => \N__30058\
        );

    \I__5481\ : InMux
    port map (
            O => \N__30064\,
            I => \N__30054\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__30061\,
            I => \N__30051\
        );

    \I__5479\ : Span4Mux_h
    port map (
            O => \N__30058\,
            I => \N__30048\
        );

    \I__5478\ : InMux
    port map (
            O => \N__30057\,
            I => \N__30045\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__30054\,
            I => \N__30042\
        );

    \I__5476\ : Span4Mux_h
    port map (
            O => \N__30051\,
            I => \N__30037\
        );

    \I__5475\ : Span4Mux_v
    port map (
            O => \N__30048\,
            I => \N__30037\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__30045\,
            I => \N__30034\
        );

    \I__5473\ : Odrv12
    port map (
            O => \N__30042\,
            I => \current_shift_inst.elapsed_time_ns_phase_25\
        );

    \I__5472\ : Odrv4
    port map (
            O => \N__30037\,
            I => \current_shift_inst.elapsed_time_ns_phase_25\
        );

    \I__5471\ : Odrv4
    port map (
            O => \N__30034\,
            I => \current_shift_inst.elapsed_time_ns_phase_25\
        );

    \I__5470\ : InMux
    port map (
            O => \N__30027\,
            I => \N__30024\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__30024\,
            I => \N__30021\
        );

    \I__5468\ : Span4Mux_h
    port map (
            O => \N__30021\,
            I => \N__30018\
        );

    \I__5467\ : Odrv4
    port map (
            O => \N__30018\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5S981_24\
        );

    \I__5466\ : CascadeMux
    port map (
            O => \N__30015\,
            I => \N__30012\
        );

    \I__5465\ : InMux
    port map (
            O => \N__30012\,
            I => \N__30003\
        );

    \I__5464\ : InMux
    port map (
            O => \N__30011\,
            I => \N__30003\
        );

    \I__5463\ : InMux
    port map (
            O => \N__30010\,
            I => \N__30003\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__30003\,
            I => \N__29999\
        );

    \I__5461\ : CascadeMux
    port map (
            O => \N__30002\,
            I => \N__29996\
        );

    \I__5460\ : Span4Mux_h
    port map (
            O => \N__29999\,
            I => \N__29993\
        );

    \I__5459\ : InMux
    port map (
            O => \N__29996\,
            I => \N__29990\
        );

    \I__5458\ : Odrv4
    port map (
            O => \N__29993\,
            I => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__29990\,
            I => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\
        );

    \I__5456\ : InMux
    port map (
            O => \N__29985\,
            I => \current_shift_inst.un4_control_input_cry_15\
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__29982\,
            I => \N__29979\
        );

    \I__5454\ : InMux
    port map (
            O => \N__29979\,
            I => \N__29970\
        );

    \I__5453\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29970\
        );

    \I__5452\ : InMux
    port map (
            O => \N__29977\,
            I => \N__29970\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__29970\,
            I => \N__29966\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__29969\,
            I => \N__29963\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__29966\,
            I => \N__29960\
        );

    \I__5448\ : InMux
    port map (
            O => \N__29963\,
            I => \N__29957\
        );

    \I__5447\ : Odrv4
    port map (
            O => \N__29960\,
            I => \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__29957\,
            I => \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\
        );

    \I__5445\ : InMux
    port map (
            O => \N__29952\,
            I => \bfn_11_18_0_\
        );

    \I__5444\ : CascadeMux
    port map (
            O => \N__29949\,
            I => \N__29946\
        );

    \I__5443\ : InMux
    port map (
            O => \N__29946\,
            I => \N__29943\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__29943\,
            I => \N__29938\
        );

    \I__5441\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29935\
        );

    \I__5440\ : InMux
    port map (
            O => \N__29941\,
            I => \N__29932\
        );

    \I__5439\ : Span4Mux_v
    port map (
            O => \N__29938\,
            I => \N__29924\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__29935\,
            I => \N__29924\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__29932\,
            I => \N__29924\
        );

    \I__5436\ : CascadeMux
    port map (
            O => \N__29931\,
            I => \N__29921\
        );

    \I__5435\ : Span4Mux_h
    port map (
            O => \N__29924\,
            I => \N__29918\
        );

    \I__5434\ : InMux
    port map (
            O => \N__29921\,
            I => \N__29915\
        );

    \I__5433\ : Odrv4
    port map (
            O => \N__29918\,
            I => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__29915\,
            I => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\
        );

    \I__5431\ : InMux
    port map (
            O => \N__29910\,
            I => \current_shift_inst.un4_control_input_cry_17\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__29907\,
            I => \N__29904\
        );

    \I__5429\ : InMux
    port map (
            O => \N__29904\,
            I => \N__29899\
        );

    \I__5428\ : InMux
    port map (
            O => \N__29903\,
            I => \N__29894\
        );

    \I__5427\ : InMux
    port map (
            O => \N__29902\,
            I => \N__29894\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__29899\,
            I => \N__29890\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__29894\,
            I => \N__29887\
        );

    \I__5424\ : CascadeMux
    port map (
            O => \N__29893\,
            I => \N__29884\
        );

    \I__5423\ : Span4Mux_h
    port map (
            O => \N__29890\,
            I => \N__29881\
        );

    \I__5422\ : Span4Mux_v
    port map (
            O => \N__29887\,
            I => \N__29878\
        );

    \I__5421\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29875\
        );

    \I__5420\ : Odrv4
    port map (
            O => \N__29881\,
            I => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\
        );

    \I__5419\ : Odrv4
    port map (
            O => \N__29878\,
            I => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__29875\,
            I => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\
        );

    \I__5417\ : InMux
    port map (
            O => \N__29868\,
            I => \current_shift_inst.un4_control_input_cry_18\
        );

    \I__5416\ : CascadeMux
    port map (
            O => \N__29865\,
            I => \N__29862\
        );

    \I__5415\ : InMux
    port map (
            O => \N__29862\,
            I => \N__29853\
        );

    \I__5414\ : InMux
    port map (
            O => \N__29861\,
            I => \N__29853\
        );

    \I__5413\ : InMux
    port map (
            O => \N__29860\,
            I => \N__29853\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__29853\,
            I => \N__29849\
        );

    \I__5411\ : CascadeMux
    port map (
            O => \N__29852\,
            I => \N__29846\
        );

    \I__5410\ : Span4Mux_h
    port map (
            O => \N__29849\,
            I => \N__29843\
        );

    \I__5409\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29840\
        );

    \I__5408\ : Odrv4
    port map (
            O => \N__29843\,
            I => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__29840\,
            I => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\
        );

    \I__5406\ : InMux
    port map (
            O => \N__29835\,
            I => \current_shift_inst.un4_control_input_cry_19\
        );

    \I__5405\ : InMux
    port map (
            O => \N__29832\,
            I => \N__29823\
        );

    \I__5404\ : InMux
    port map (
            O => \N__29831\,
            I => \N__29823\
        );

    \I__5403\ : InMux
    port map (
            O => \N__29830\,
            I => \N__29823\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__29823\,
            I => \N__29820\
        );

    \I__5401\ : Span4Mux_v
    port map (
            O => \N__29820\,
            I => \N__29816\
        );

    \I__5400\ : InMux
    port map (
            O => \N__29819\,
            I => \N__29813\
        );

    \I__5399\ : Odrv4
    port map (
            O => \N__29816\,
            I => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__29813\,
            I => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\
        );

    \I__5397\ : InMux
    port map (
            O => \N__29808\,
            I => \current_shift_inst.un4_control_input_cry_20\
        );

    \I__5396\ : CascadeMux
    port map (
            O => \N__29805\,
            I => \N__29802\
        );

    \I__5395\ : InMux
    port map (
            O => \N__29802\,
            I => \N__29793\
        );

    \I__5394\ : InMux
    port map (
            O => \N__29801\,
            I => \N__29793\
        );

    \I__5393\ : InMux
    port map (
            O => \N__29800\,
            I => \N__29793\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__29793\,
            I => \N__29789\
        );

    \I__5391\ : CascadeMux
    port map (
            O => \N__29792\,
            I => \N__29786\
        );

    \I__5390\ : Span4Mux_v
    port map (
            O => \N__29789\,
            I => \N__29783\
        );

    \I__5389\ : InMux
    port map (
            O => \N__29786\,
            I => \N__29780\
        );

    \I__5388\ : Odrv4
    port map (
            O => \N__29783\,
            I => \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__29780\,
            I => \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\
        );

    \I__5386\ : InMux
    port map (
            O => \N__29775\,
            I => \current_shift_inst.un4_control_input_cry_21\
        );

    \I__5385\ : InMux
    port map (
            O => \N__29772\,
            I => \current_shift_inst.un4_control_input_cry_22\
        );

    \I__5384\ : InMux
    port map (
            O => \N__29769\,
            I => \current_shift_inst.un4_control_input_cry_23\
        );

    \I__5383\ : InMux
    port map (
            O => \N__29766\,
            I => \N__29763\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__29763\,
            I => \current_shift_inst.un4_control_input_axb_8\
        );

    \I__5381\ : InMux
    port map (
            O => \N__29760\,
            I => \N__29755\
        );

    \I__5380\ : InMux
    port map (
            O => \N__29759\,
            I => \N__29750\
        );

    \I__5379\ : InMux
    port map (
            O => \N__29758\,
            I => \N__29750\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__29755\,
            I => \N__29744\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__29750\,
            I => \N__29744\
        );

    \I__5376\ : CascadeMux
    port map (
            O => \N__29749\,
            I => \N__29741\
        );

    \I__5375\ : Span4Mux_h
    port map (
            O => \N__29744\,
            I => \N__29738\
        );

    \I__5374\ : InMux
    port map (
            O => \N__29741\,
            I => \N__29735\
        );

    \I__5373\ : Odrv4
    port map (
            O => \N__29738\,
            I => \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__29735\,
            I => \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\
        );

    \I__5371\ : InMux
    port map (
            O => \N__29730\,
            I => \current_shift_inst.un4_control_input_cry_7\
        );

    \I__5370\ : InMux
    port map (
            O => \N__29727\,
            I => \N__29724\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__29724\,
            I => \N__29721\
        );

    \I__5368\ : Odrv4
    port map (
            O => \N__29721\,
            I => \current_shift_inst.un4_control_input_axb_9\
        );

    \I__5367\ : CascadeMux
    port map (
            O => \N__29718\,
            I => \N__29714\
        );

    \I__5366\ : CascadeMux
    port map (
            O => \N__29717\,
            I => \N__29711\
        );

    \I__5365\ : InMux
    port map (
            O => \N__29714\,
            I => \N__29707\
        );

    \I__5364\ : InMux
    port map (
            O => \N__29711\,
            I => \N__29702\
        );

    \I__5363\ : InMux
    port map (
            O => \N__29710\,
            I => \N__29702\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__29707\,
            I => \N__29698\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__29702\,
            I => \N__29695\
        );

    \I__5360\ : CascadeMux
    port map (
            O => \N__29701\,
            I => \N__29692\
        );

    \I__5359\ : Span4Mux_h
    port map (
            O => \N__29698\,
            I => \N__29689\
        );

    \I__5358\ : Span4Mux_h
    port map (
            O => \N__29695\,
            I => \N__29686\
        );

    \I__5357\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29683\
        );

    \I__5356\ : Odrv4
    port map (
            O => \N__29689\,
            I => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\
        );

    \I__5355\ : Odrv4
    port map (
            O => \N__29686\,
            I => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\
        );

    \I__5354\ : LocalMux
    port map (
            O => \N__29683\,
            I => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\
        );

    \I__5353\ : InMux
    port map (
            O => \N__29676\,
            I => \bfn_11_17_0_\
        );

    \I__5352\ : CascadeMux
    port map (
            O => \N__29673\,
            I => \N__29669\
        );

    \I__5351\ : InMux
    port map (
            O => \N__29672\,
            I => \N__29665\
        );

    \I__5350\ : InMux
    port map (
            O => \N__29669\,
            I => \N__29660\
        );

    \I__5349\ : InMux
    port map (
            O => \N__29668\,
            I => \N__29660\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__29665\,
            I => \N__29654\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__29660\,
            I => \N__29654\
        );

    \I__5346\ : CascadeMux
    port map (
            O => \N__29659\,
            I => \N__29651\
        );

    \I__5345\ : Span4Mux_h
    port map (
            O => \N__29654\,
            I => \N__29648\
        );

    \I__5344\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29645\
        );

    \I__5343\ : Odrv4
    port map (
            O => \N__29648\,
            I => \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__29645\,
            I => \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\
        );

    \I__5341\ : InMux
    port map (
            O => \N__29640\,
            I => \current_shift_inst.un4_control_input_cry_9\
        );

    \I__5340\ : InMux
    port map (
            O => \N__29637\,
            I => \N__29628\
        );

    \I__5339\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29628\
        );

    \I__5338\ : InMux
    port map (
            O => \N__29635\,
            I => \N__29628\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__29628\,
            I => \N__29624\
        );

    \I__5336\ : CascadeMux
    port map (
            O => \N__29627\,
            I => \N__29621\
        );

    \I__5335\ : Span4Mux_h
    port map (
            O => \N__29624\,
            I => \N__29618\
        );

    \I__5334\ : InMux
    port map (
            O => \N__29621\,
            I => \N__29615\
        );

    \I__5333\ : Odrv4
    port map (
            O => \N__29618\,
            I => \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__29615\,
            I => \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\
        );

    \I__5331\ : InMux
    port map (
            O => \N__29610\,
            I => \current_shift_inst.un4_control_input_cry_10\
        );

    \I__5330\ : CascadeMux
    port map (
            O => \N__29607\,
            I => \N__29602\
        );

    \I__5329\ : InMux
    port map (
            O => \N__29606\,
            I => \N__29599\
        );

    \I__5328\ : InMux
    port map (
            O => \N__29605\,
            I => \N__29594\
        );

    \I__5327\ : InMux
    port map (
            O => \N__29602\,
            I => \N__29594\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__29599\,
            I => \N__29588\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__29594\,
            I => \N__29588\
        );

    \I__5324\ : CascadeMux
    port map (
            O => \N__29593\,
            I => \N__29585\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__29588\,
            I => \N__29582\
        );

    \I__5322\ : InMux
    port map (
            O => \N__29585\,
            I => \N__29579\
        );

    \I__5321\ : Odrv4
    port map (
            O => \N__29582\,
            I => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__29579\,
            I => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\
        );

    \I__5319\ : InMux
    port map (
            O => \N__29574\,
            I => \current_shift_inst.un4_control_input_cry_11\
        );

    \I__5318\ : CascadeMux
    port map (
            O => \N__29571\,
            I => \N__29568\
        );

    \I__5317\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29564\
        );

    \I__5316\ : InMux
    port map (
            O => \N__29567\,
            I => \N__29560\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__29564\,
            I => \N__29556\
        );

    \I__5314\ : InMux
    port map (
            O => \N__29563\,
            I => \N__29553\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__29560\,
            I => \N__29550\
        );

    \I__5312\ : CascadeMux
    port map (
            O => \N__29559\,
            I => \N__29547\
        );

    \I__5311\ : Span4Mux_v
    port map (
            O => \N__29556\,
            I => \N__29540\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__29553\,
            I => \N__29540\
        );

    \I__5309\ : Span4Mux_h
    port map (
            O => \N__29550\,
            I => \N__29540\
        );

    \I__5308\ : InMux
    port map (
            O => \N__29547\,
            I => \N__29537\
        );

    \I__5307\ : Odrv4
    port map (
            O => \N__29540\,
            I => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__29537\,
            I => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\
        );

    \I__5305\ : InMux
    port map (
            O => \N__29532\,
            I => \current_shift_inst.un4_control_input_cry_12\
        );

    \I__5304\ : CascadeMux
    port map (
            O => \N__29529\,
            I => \N__29526\
        );

    \I__5303\ : InMux
    port map (
            O => \N__29526\,
            I => \N__29523\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__29523\,
            I => \N__29518\
        );

    \I__5301\ : InMux
    port map (
            O => \N__29522\,
            I => \N__29513\
        );

    \I__5300\ : InMux
    port map (
            O => \N__29521\,
            I => \N__29513\
        );

    \I__5299\ : Span4Mux_v
    port map (
            O => \N__29518\,
            I => \N__29509\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__29513\,
            I => \N__29506\
        );

    \I__5297\ : CascadeMux
    port map (
            O => \N__29512\,
            I => \N__29503\
        );

    \I__5296\ : Span4Mux_h
    port map (
            O => \N__29509\,
            I => \N__29498\
        );

    \I__5295\ : Span4Mux_v
    port map (
            O => \N__29506\,
            I => \N__29498\
        );

    \I__5294\ : InMux
    port map (
            O => \N__29503\,
            I => \N__29495\
        );

    \I__5293\ : Odrv4
    port map (
            O => \N__29498\,
            I => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__29495\,
            I => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\
        );

    \I__5291\ : InMux
    port map (
            O => \N__29490\,
            I => \current_shift_inst.un4_control_input_cry_13\
        );

    \I__5290\ : CascadeMux
    port map (
            O => \N__29487\,
            I => \N__29484\
        );

    \I__5289\ : InMux
    port map (
            O => \N__29484\,
            I => \N__29477\
        );

    \I__5288\ : InMux
    port map (
            O => \N__29483\,
            I => \N__29477\
        );

    \I__5287\ : InMux
    port map (
            O => \N__29482\,
            I => \N__29474\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__29477\,
            I => \N__29468\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__29474\,
            I => \N__29468\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__29473\,
            I => \N__29465\
        );

    \I__5283\ : Span4Mux_h
    port map (
            O => \N__29468\,
            I => \N__29462\
        );

    \I__5282\ : InMux
    port map (
            O => \N__29465\,
            I => \N__29459\
        );

    \I__5281\ : Odrv4
    port map (
            O => \N__29462\,
            I => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__29459\,
            I => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\
        );

    \I__5279\ : InMux
    port map (
            O => \N__29454\,
            I => \current_shift_inst.un4_control_input_cry_14\
        );

    \I__5278\ : InMux
    port map (
            O => \N__29451\,
            I => \N__29448\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__29448\,
            I => \N__29445\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__29445\,
            I => \current_shift_inst.un4_control_input_axb_1\
        );

    \I__5275\ : InMux
    port map (
            O => \N__29442\,
            I => \N__29437\
        );

    \I__5274\ : CascadeMux
    port map (
            O => \N__29441\,
            I => \N__29434\
        );

    \I__5273\ : InMux
    port map (
            O => \N__29440\,
            I => \N__29431\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__29437\,
            I => \N__29428\
        );

    \I__5271\ : InMux
    port map (
            O => \N__29434\,
            I => \N__29425\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__29431\,
            I => \current_shift_inst.elapsed_time_ns_1_fast_31\
        );

    \I__5269\ : Odrv4
    port map (
            O => \N__29428\,
            I => \current_shift_inst.elapsed_time_ns_1_fast_31\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__29425\,
            I => \current_shift_inst.elapsed_time_ns_1_fast_31\
        );

    \I__5267\ : CascadeMux
    port map (
            O => \N__29418\,
            I => \N__29415\
        );

    \I__5266\ : InMux
    port map (
            O => \N__29415\,
            I => \N__29412\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__29412\,
            I => \N__29409\
        );

    \I__5264\ : Span4Mux_h
    port map (
            O => \N__29409\,
            I => \N__29405\
        );

    \I__5263\ : InMux
    port map (
            O => \N__29408\,
            I => \N__29402\
        );

    \I__5262\ : Odrv4
    port map (
            O => \N__29405\,
            I => \current_shift_inst.un38_control_input_0\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__29402\,
            I => \current_shift_inst.un38_control_input_0\
        );

    \I__5260\ : InMux
    port map (
            O => \N__29397\,
            I => \N__29394\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__29394\,
            I => \N__29391\
        );

    \I__5258\ : Odrv4
    port map (
            O => \N__29391\,
            I => \current_shift_inst.un4_control_input_axb_2\
        );

    \I__5257\ : InMux
    port map (
            O => \N__29388\,
            I => \N__29385\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__29385\,
            I => \N__29381\
        );

    \I__5255\ : InMux
    port map (
            O => \N__29384\,
            I => \N__29377\
        );

    \I__5254\ : Span4Mux_h
    port map (
            O => \N__29381\,
            I => \N__29374\
        );

    \I__5253\ : InMux
    port map (
            O => \N__29380\,
            I => \N__29371\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__29377\,
            I => \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\
        );

    \I__5251\ : Odrv4
    port map (
            O => \N__29374\,
            I => \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__29371\,
            I => \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\
        );

    \I__5249\ : InMux
    port map (
            O => \N__29364\,
            I => \current_shift_inst.un4_control_input_cry_1\
        );

    \I__5248\ : InMux
    port map (
            O => \N__29361\,
            I => \N__29358\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__29358\,
            I => \N__29355\
        );

    \I__5246\ : Odrv4
    port map (
            O => \N__29355\,
            I => \current_shift_inst.un4_control_input_axb_3\
        );

    \I__5245\ : InMux
    port map (
            O => \N__29352\,
            I => \N__29349\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__29349\,
            I => \N__29345\
        );

    \I__5243\ : InMux
    port map (
            O => \N__29348\,
            I => \N__29341\
        );

    \I__5242\ : Span4Mux_h
    port map (
            O => \N__29345\,
            I => \N__29338\
        );

    \I__5241\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29335\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__29341\,
            I => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__29338\,
            I => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__29335\,
            I => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\
        );

    \I__5237\ : InMux
    port map (
            O => \N__29328\,
            I => \current_shift_inst.un4_control_input_cry_2\
        );

    \I__5236\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29322\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__29322\,
            I => \current_shift_inst.un4_control_input_axb_4\
        );

    \I__5234\ : InMux
    port map (
            O => \N__29319\,
            I => \N__29316\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__29316\,
            I => \N__29313\
        );

    \I__5232\ : Span4Mux_h
    port map (
            O => \N__29313\,
            I => \N__29309\
        );

    \I__5231\ : InMux
    port map (
            O => \N__29312\,
            I => \N__29306\
        );

    \I__5230\ : Odrv4
    port map (
            O => \N__29309\,
            I => \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__29306\,
            I => \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\
        );

    \I__5228\ : InMux
    port map (
            O => \N__29301\,
            I => \current_shift_inst.un4_control_input_cry_3\
        );

    \I__5227\ : InMux
    port map (
            O => \N__29298\,
            I => \N__29295\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__29295\,
            I => \current_shift_inst.un4_control_input_axb_5\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__29292\,
            I => \N__29289\
        );

    \I__5224\ : InMux
    port map (
            O => \N__29289\,
            I => \N__29286\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__29286\,
            I => \N__29282\
        );

    \I__5222\ : CascadeMux
    port map (
            O => \N__29285\,
            I => \N__29277\
        );

    \I__5221\ : Span4Mux_v
    port map (
            O => \N__29282\,
            I => \N__29274\
        );

    \I__5220\ : InMux
    port map (
            O => \N__29281\,
            I => \N__29269\
        );

    \I__5219\ : InMux
    port map (
            O => \N__29280\,
            I => \N__29269\
        );

    \I__5218\ : InMux
    port map (
            O => \N__29277\,
            I => \N__29266\
        );

    \I__5217\ : Odrv4
    port map (
            O => \N__29274\,
            I => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__29269\,
            I => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__29266\,
            I => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\
        );

    \I__5214\ : InMux
    port map (
            O => \N__29259\,
            I => \current_shift_inst.un4_control_input_cry_4\
        );

    \I__5213\ : InMux
    port map (
            O => \N__29256\,
            I => \N__29253\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__29253\,
            I => \current_shift_inst.un4_control_input_axb_6\
        );

    \I__5211\ : InMux
    port map (
            O => \N__29250\,
            I => \N__29245\
        );

    \I__5210\ : InMux
    port map (
            O => \N__29249\,
            I => \N__29240\
        );

    \I__5209\ : InMux
    port map (
            O => \N__29248\,
            I => \N__29240\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__29245\,
            I => \N__29234\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__29240\,
            I => \N__29234\
        );

    \I__5206\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29231\
        );

    \I__5205\ : Odrv4
    port map (
            O => \N__29234\,
            I => \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__29231\,
            I => \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\
        );

    \I__5203\ : InMux
    port map (
            O => \N__29226\,
            I => \current_shift_inst.un4_control_input_cry_5\
        );

    \I__5202\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29220\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__29220\,
            I => \current_shift_inst.un4_control_input_axb_7\
        );

    \I__5200\ : InMux
    port map (
            O => \N__29217\,
            I => \N__29211\
        );

    \I__5199\ : InMux
    port map (
            O => \N__29216\,
            I => \N__29211\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__29211\,
            I => \N__29207\
        );

    \I__5197\ : InMux
    port map (
            O => \N__29210\,
            I => \N__29204\
        );

    \I__5196\ : Span4Mux_h
    port map (
            O => \N__29207\,
            I => \N__29200\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__29204\,
            I => \N__29197\
        );

    \I__5194\ : InMux
    port map (
            O => \N__29203\,
            I => \N__29194\
        );

    \I__5193\ : Odrv4
    port map (
            O => \N__29200\,
            I => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\
        );

    \I__5192\ : Odrv12
    port map (
            O => \N__29197\,
            I => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__29194\,
            I => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\
        );

    \I__5190\ : InMux
    port map (
            O => \N__29187\,
            I => \current_shift_inst.un4_control_input_cry_6\
        );

    \I__5189\ : InMux
    port map (
            O => \N__29184\,
            I => \N__29181\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__29181\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_1\
        );

    \I__5187\ : InMux
    port map (
            O => \N__29178\,
            I => \N__29175\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__29175\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_2\
        );

    \I__5185\ : InMux
    port map (
            O => \N__29172\,
            I => \N__29168\
        );

    \I__5184\ : InMux
    port map (
            O => \N__29171\,
            I => \N__29165\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__29168\,
            I => measured_delay_hc_27
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__29165\,
            I => measured_delay_hc_27
        );

    \I__5181\ : InMux
    port map (
            O => \N__29160\,
            I => \N__29157\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__29157\,
            I => \N__29154\
        );

    \I__5179\ : Odrv4
    port map (
            O => \N__29154\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4\
        );

    \I__5178\ : CascadeMux
    port map (
            O => \N__29151\,
            I => \N__29148\
        );

    \I__5177\ : InMux
    port map (
            O => \N__29148\,
            I => \N__29145\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__29145\,
            I => \N__29142\
        );

    \I__5175\ : Span4Mux_v
    port map (
            O => \N__29142\,
            I => \N__29139\
        );

    \I__5174\ : Odrv4
    port map (
            O => \N__29139\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25\
        );

    \I__5173\ : CascadeMux
    port map (
            O => \N__29136\,
            I => \N__29133\
        );

    \I__5172\ : InMux
    port map (
            O => \N__29133\,
            I => \N__29126\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29132\,
            I => \N__29126\
        );

    \I__5170\ : InMux
    port map (
            O => \N__29131\,
            I => \N__29123\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__29126\,
            I => \N__29118\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__29123\,
            I => \N__29118\
        );

    \I__5167\ : Span4Mux_h
    port map (
            O => \N__29118\,
            I => \N__29114\
        );

    \I__5166\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29111\
        );

    \I__5165\ : Odrv4
    port map (
            O => \N__29114\,
            I => \current_shift_inst.elapsed_time_ns_phase_6\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__29111\,
            I => \current_shift_inst.elapsed_time_ns_phase_6\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__29106\,
            I => \N__29103\
        );

    \I__5162\ : InMux
    port map (
            O => \N__29103\,
            I => \N__29098\
        );

    \I__5161\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29093\
        );

    \I__5160\ : InMux
    port map (
            O => \N__29101\,
            I => \N__29093\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__29098\,
            I => \N__29088\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__29093\,
            I => \N__29088\
        );

    \I__5157\ : Span4Mux_h
    port map (
            O => \N__29088\,
            I => \N__29084\
        );

    \I__5156\ : InMux
    port map (
            O => \N__29087\,
            I => \N__29081\
        );

    \I__5155\ : Odrv4
    port map (
            O => \N__29084\,
            I => \current_shift_inst.elapsed_time_ns_phase_5\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__29081\,
            I => \current_shift_inst.elapsed_time_ns_phase_5\
        );

    \I__5153\ : InMux
    port map (
            O => \N__29076\,
            I => \N__29073\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__29073\,
            I => \N__29070\
        );

    \I__5151\ : Odrv12
    port map (
            O => \N__29070\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5\
        );

    \I__5150\ : InMux
    port map (
            O => \N__29067\,
            I => \N__29063\
        );

    \I__5149\ : InMux
    port map (
            O => \N__29066\,
            I => \N__29060\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__29063\,
            I => measured_delay_hc_23
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__29060\,
            I => measured_delay_hc_23
        );

    \I__5146\ : CascadeMux
    port map (
            O => \N__29055\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_3_cascade_\
        );

    \I__5145\ : InMux
    port map (
            O => \N__29052\,
            I => \N__29046\
        );

    \I__5144\ : InMux
    port map (
            O => \N__29051\,
            I => \N__29046\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__29046\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_14\
        );

    \I__5142\ : InMux
    port map (
            O => \N__29043\,
            I => \N__29040\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__29040\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\
        );

    \I__5140\ : CascadeMux
    port map (
            O => \N__29037\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt30_0_cascade_\
        );

    \I__5139\ : InMux
    port map (
            O => \N__29034\,
            I => \N__29031\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__29031\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6\
        );

    \I__5137\ : InMux
    port map (
            O => \N__29028\,
            I => \N__29025\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__29025\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_6\
        );

    \I__5135\ : IoInMux
    port map (
            O => \N__29022\,
            I => \N__29019\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__29019\,
            I => \N__29016\
        );

    \I__5133\ : IoSpan4Mux
    port map (
            O => \N__29016\,
            I => \N__29013\
        );

    \I__5132\ : IoSpan4Mux
    port map (
            O => \N__29013\,
            I => \N__29010\
        );

    \I__5131\ : Span4Mux_s1_v
    port map (
            O => \N__29010\,
            I => \N__29007\
        );

    \I__5130\ : Sp12to4
    port map (
            O => \N__29007\,
            I => \N__29004\
        );

    \I__5129\ : Span12Mux_s9_v
    port map (
            O => \N__29004\,
            I => \N__29001\
        );

    \I__5128\ : Odrv12
    port map (
            O => \N__29001\,
            I => \current_shift_inst.timer_s1.N_187_i\
        );

    \I__5127\ : InMux
    port map (
            O => \N__28998\,
            I => \N__28995\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__28995\,
            I => \N__28991\
        );

    \I__5125\ : CascadeMux
    port map (
            O => \N__28994\,
            I => \N__28988\
        );

    \I__5124\ : Span4Mux_v
    port map (
            O => \N__28991\,
            I => \N__28983\
        );

    \I__5123\ : InMux
    port map (
            O => \N__28988\,
            I => \N__28977\
        );

    \I__5122\ : InMux
    port map (
            O => \N__28987\,
            I => \N__28977\
        );

    \I__5121\ : InMux
    port map (
            O => \N__28986\,
            I => \N__28974\
        );

    \I__5120\ : Span4Mux_h
    port map (
            O => \N__28983\,
            I => \N__28971\
        );

    \I__5119\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28968\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__28977\,
            I => \current_shift_inst.phase_validZ0\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__28974\,
            I => \current_shift_inst.phase_validZ0\
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__28971\,
            I => \current_shift_inst.phase_validZ0\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__28968\,
            I => \current_shift_inst.phase_validZ0\
        );

    \I__5114\ : CascadeMux
    port map (
            O => \N__28959\,
            I => \N__28955\
        );

    \I__5113\ : InMux
    port map (
            O => \N__28958\,
            I => \N__28951\
        );

    \I__5112\ : InMux
    port map (
            O => \N__28955\,
            I => \N__28948\
        );

    \I__5111\ : InMux
    port map (
            O => \N__28954\,
            I => \N__28945\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__28951\,
            I => measured_delay_hc_20
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__28948\,
            I => measured_delay_hc_20
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__28945\,
            I => measured_delay_hc_20
        );

    \I__5107\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28935\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__28935\,
            I => \current_shift_inst.z_5_27\
        );

    \I__5105\ : InMux
    port map (
            O => \N__28932\,
            I => \N__28929\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__28929\,
            I => \current_shift_inst.z_5_28\
        );

    \I__5103\ : CascadeMux
    port map (
            O => \N__28926\,
            I => \N__28923\
        );

    \I__5102\ : InMux
    port map (
            O => \N__28923\,
            I => \N__28920\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__28920\,
            I => \current_shift_inst.z_5_29\
        );

    \I__5100\ : CascadeMux
    port map (
            O => \N__28917\,
            I => \N__28914\
        );

    \I__5099\ : InMux
    port map (
            O => \N__28914\,
            I => \N__28911\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__28911\,
            I => \current_shift_inst.z_5_30\
        );

    \I__5097\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28905\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__28905\,
            I => \current_shift_inst.z_5_cry_30_THRU_CO\
        );

    \I__5095\ : InMux
    port map (
            O => \N__28902\,
            I => \current_shift_inst.z_cry_30\
        );

    \I__5094\ : CascadeMux
    port map (
            O => \N__28899\,
            I => \N__28894\
        );

    \I__5093\ : InMux
    port map (
            O => \N__28898\,
            I => \N__28889\
        );

    \I__5092\ : InMux
    port map (
            O => \N__28897\,
            I => \N__28889\
        );

    \I__5091\ : InMux
    port map (
            O => \N__28894\,
            I => \N__28886\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__28889\,
            I => \N__28883\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__28886\,
            I => measured_delay_hc_21
        );

    \I__5088\ : Odrv4
    port map (
            O => \N__28883\,
            I => measured_delay_hc_21
        );

    \I__5087\ : CascadeMux
    port map (
            O => \N__28878\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0_cascade_\
        );

    \I__5086\ : InMux
    port map (
            O => \N__28875\,
            I => \N__28872\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__28872\,
            I => \current_shift_inst.z_5_19\
        );

    \I__5084\ : CascadeMux
    port map (
            O => \N__28869\,
            I => \N__28866\
        );

    \I__5083\ : InMux
    port map (
            O => \N__28866\,
            I => \N__28863\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__28863\,
            I => \current_shift_inst.z_5_20\
        );

    \I__5081\ : InMux
    port map (
            O => \N__28860\,
            I => \N__28857\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__28857\,
            I => \current_shift_inst.z_5_21\
        );

    \I__5079\ : InMux
    port map (
            O => \N__28854\,
            I => \N__28851\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__28851\,
            I => \current_shift_inst.z_5_22\
        );

    \I__5077\ : InMux
    port map (
            O => \N__28848\,
            I => \N__28845\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__28845\,
            I => \current_shift_inst.z_5_23\
        );

    \I__5075\ : InMux
    port map (
            O => \N__28842\,
            I => \N__28839\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__28839\,
            I => \current_shift_inst.z_5_24\
        );

    \I__5073\ : CascadeMux
    port map (
            O => \N__28836\,
            I => \N__28833\
        );

    \I__5072\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28830\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__28830\,
            I => \current_shift_inst.z_5_25\
        );

    \I__5070\ : InMux
    port map (
            O => \N__28827\,
            I => \N__28824\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__28824\,
            I => \current_shift_inst.z_5_26\
        );

    \I__5068\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28818\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__28818\,
            I => \current_shift_inst.z_5_10\
        );

    \I__5066\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28812\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__28812\,
            I => \current_shift_inst.z_5_11\
        );

    \I__5064\ : InMux
    port map (
            O => \N__28809\,
            I => \N__28806\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__28806\,
            I => \current_shift_inst.z_5_12\
        );

    \I__5062\ : InMux
    port map (
            O => \N__28803\,
            I => \N__28800\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__28800\,
            I => \current_shift_inst.z_5_13\
        );

    \I__5060\ : InMux
    port map (
            O => \N__28797\,
            I => \N__28794\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__28794\,
            I => \current_shift_inst.z_5_14\
        );

    \I__5058\ : InMux
    port map (
            O => \N__28791\,
            I => \N__28788\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__28788\,
            I => \current_shift_inst.z_5_15\
        );

    \I__5056\ : InMux
    port map (
            O => \N__28785\,
            I => \N__28782\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__28782\,
            I => \N__28779\
        );

    \I__5054\ : Odrv4
    port map (
            O => \N__28779\,
            I => \current_shift_inst.z_5_16\
        );

    \I__5053\ : InMux
    port map (
            O => \N__28776\,
            I => \N__28773\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__28773\,
            I => \current_shift_inst.z_5_17\
        );

    \I__5051\ : InMux
    port map (
            O => \N__28770\,
            I => \N__28767\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__28767\,
            I => \current_shift_inst.z_5_18\
        );

    \I__5049\ : CascadeMux
    port map (
            O => \N__28764\,
            I => \N__28761\
        );

    \I__5048\ : InMux
    port map (
            O => \N__28761\,
            I => \N__28758\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__28758\,
            I => \current_shift_inst.z_5_2\
        );

    \I__5046\ : CascadeMux
    port map (
            O => \N__28755\,
            I => \N__28752\
        );

    \I__5045\ : InMux
    port map (
            O => \N__28752\,
            I => \N__28749\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__28749\,
            I => \current_shift_inst.z_5_3\
        );

    \I__5043\ : InMux
    port map (
            O => \N__28746\,
            I => \N__28743\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__28743\,
            I => \current_shift_inst.z_5_4\
        );

    \I__5041\ : CascadeMux
    port map (
            O => \N__28740\,
            I => \N__28737\
        );

    \I__5040\ : InMux
    port map (
            O => \N__28737\,
            I => \N__28734\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__28734\,
            I => \current_shift_inst.z_5_5\
        );

    \I__5038\ : CascadeMux
    port map (
            O => \N__28731\,
            I => \N__28728\
        );

    \I__5037\ : InMux
    port map (
            O => \N__28728\,
            I => \N__28725\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__28725\,
            I => \current_shift_inst.z_5_6\
        );

    \I__5035\ : InMux
    port map (
            O => \N__28722\,
            I => \N__28719\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__28719\,
            I => \current_shift_inst.z_5_7\
        );

    \I__5033\ : InMux
    port map (
            O => \N__28716\,
            I => \N__28713\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__28713\,
            I => \N__28710\
        );

    \I__5031\ : Odrv4
    port map (
            O => \N__28710\,
            I => \current_shift_inst.z_5_8\
        );

    \I__5030\ : InMux
    port map (
            O => \N__28707\,
            I => \N__28704\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__28704\,
            I => \current_shift_inst.z_5_9\
        );

    \I__5028\ : InMux
    port map (
            O => \N__28701\,
            I => \N__28697\
        );

    \I__5027\ : InMux
    port map (
            O => \N__28700\,
            I => \N__28694\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__28697\,
            I => \N__28691\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__28694\,
            I => \N__28688\
        );

    \I__5024\ : Span4Mux_h
    port map (
            O => \N__28691\,
            I => \N__28684\
        );

    \I__5023\ : Span4Mux_h
    port map (
            O => \N__28688\,
            I => \N__28681\
        );

    \I__5022\ : InMux
    port map (
            O => \N__28687\,
            I => \N__28678\
        );

    \I__5021\ : Odrv4
    port map (
            O => \N__28684\,
            I => \current_shift_inst.timer_phase.counterZ0Z_1\
        );

    \I__5020\ : Odrv4
    port map (
            O => \N__28681\,
            I => \current_shift_inst.timer_phase.counterZ0Z_1\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__28678\,
            I => \current_shift_inst.timer_phase.counterZ0Z_1\
        );

    \I__5018\ : InMux
    port map (
            O => \N__28671\,
            I => \N__28668\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__28668\,
            I => \N__28665\
        );

    \I__5016\ : Span4Mux_v
    port map (
            O => \N__28665\,
            I => \N__28662\
        );

    \I__5015\ : Odrv4
    port map (
            O => \N__28662\,
            I => \current_shift_inst.N_1633_i\
        );

    \I__5014\ : InMux
    port map (
            O => \N__28659\,
            I => \N__28656\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__28656\,
            I => \N__28652\
        );

    \I__5012\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28649\
        );

    \I__5011\ : Span4Mux_h
    port map (
            O => \N__28652\,
            I => \N__28645\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__28649\,
            I => \N__28642\
        );

    \I__5009\ : InMux
    port map (
            O => \N__28648\,
            I => \N__28639\
        );

    \I__5008\ : Odrv4
    port map (
            O => \N__28645\,
            I => \current_shift_inst.timer_phase.counterZ0Z_0\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__28642\,
            I => \current_shift_inst.timer_phase.counterZ0Z_0\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__28639\,
            I => \current_shift_inst.timer_phase.counterZ0Z_0\
        );

    \I__5005\ : CEMux
    port map (
            O => \N__28632\,
            I => \N__28617\
        );

    \I__5004\ : CEMux
    port map (
            O => \N__28631\,
            I => \N__28617\
        );

    \I__5003\ : CEMux
    port map (
            O => \N__28630\,
            I => \N__28617\
        );

    \I__5002\ : CEMux
    port map (
            O => \N__28629\,
            I => \N__28617\
        );

    \I__5001\ : CEMux
    port map (
            O => \N__28628\,
            I => \N__28617\
        );

    \I__5000\ : GlobalMux
    port map (
            O => \N__28617\,
            I => \N__28614\
        );

    \I__4999\ : gio2CtrlBuf
    port map (
            O => \N__28614\,
            I => \current_shift_inst.timer_phase.N_188_i_g\
        );

    \I__4998\ : CascadeMux
    port map (
            O => \N__28611\,
            I => \N__28608\
        );

    \I__4997\ : InMux
    port map (
            O => \N__28608\,
            I => \N__28605\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__28605\,
            I => \N__28602\
        );

    \I__4995\ : Span4Mux_v
    port map (
            O => \N__28602\,
            I => \N__28599\
        );

    \I__4994\ : Odrv4
    port map (
            O => \N__28599\,
            I => \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0\
        );

    \I__4993\ : InMux
    port map (
            O => \N__28596\,
            I => \N__28590\
        );

    \I__4992\ : InMux
    port map (
            O => \N__28595\,
            I => \N__28590\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__28590\,
            I => \N__28586\
        );

    \I__4990\ : CascadeMux
    port map (
            O => \N__28589\,
            I => \N__28583\
        );

    \I__4989\ : Span4Mux_v
    port map (
            O => \N__28586\,
            I => \N__28580\
        );

    \I__4988\ : InMux
    port map (
            O => \N__28583\,
            I => \N__28577\
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__28580\,
            I => \current_shift_inst.elapsed_time_ns_phase_3\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__28577\,
            I => \current_shift_inst.elapsed_time_ns_phase_3\
        );

    \I__4985\ : CascadeMux
    port map (
            O => \N__28572\,
            I => \N__28567\
        );

    \I__4984\ : InMux
    port map (
            O => \N__28571\,
            I => \N__28563\
        );

    \I__4983\ : InMux
    port map (
            O => \N__28570\,
            I => \N__28560\
        );

    \I__4982\ : InMux
    port map (
            O => \N__28567\,
            I => \N__28555\
        );

    \I__4981\ : InMux
    port map (
            O => \N__28566\,
            I => \N__28555\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__28563\,
            I => \N__28552\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__28560\,
            I => \current_shift_inst.elapsed_time_ns_phase_2\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__28555\,
            I => \current_shift_inst.elapsed_time_ns_phase_2\
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__28552\,
            I => \current_shift_inst.elapsed_time_ns_phase_2\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__28545\,
            I => \N__28542\
        );

    \I__4975\ : InMux
    port map (
            O => \N__28542\,
            I => \N__28539\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__28539\,
            I => \N__28536\
        );

    \I__4973\ : Span4Mux_v
    port map (
            O => \N__28536\,
            I => \N__28533\
        );

    \I__4972\ : Odrv4
    port map (
            O => \N__28533\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3\
        );

    \I__4971\ : CascadeMux
    port map (
            O => \N__28530\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3_cascade_\
        );

    \I__4970\ : InMux
    port map (
            O => \N__28527\,
            I => \N__28524\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__28524\,
            I => \N__28521\
        );

    \I__4968\ : Span4Mux_h
    port map (
            O => \N__28521\,
            I => \N__28518\
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__28518\,
            I => \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0\
        );

    \I__4966\ : InMux
    port map (
            O => \N__28515\,
            I => \N__28511\
        );

    \I__4965\ : CascadeMux
    port map (
            O => \N__28514\,
            I => \N__28508\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__28511\,
            I => \N__28504\
        );

    \I__4963\ : InMux
    port map (
            O => \N__28508\,
            I => \N__28499\
        );

    \I__4962\ : InMux
    port map (
            O => \N__28507\,
            I => \N__28499\
        );

    \I__4961\ : Span4Mux_h
    port map (
            O => \N__28504\,
            I => \N__28494\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__28499\,
            I => \N__28494\
        );

    \I__4959\ : Span4Mux_v
    port map (
            O => \N__28494\,
            I => \N__28490\
        );

    \I__4958\ : InMux
    port map (
            O => \N__28493\,
            I => \N__28487\
        );

    \I__4957\ : Odrv4
    port map (
            O => \N__28490\,
            I => \current_shift_inst.elapsed_time_ns_phase_4\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__28487\,
            I => \current_shift_inst.elapsed_time_ns_phase_4\
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__28482\,
            I => \N__28479\
        );

    \I__4954\ : InMux
    port map (
            O => \N__28479\,
            I => \N__28476\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__28476\,
            I => \N__28473\
        );

    \I__4952\ : Span4Mux_h
    port map (
            O => \N__28473\,
            I => \N__28470\
        );

    \I__4951\ : Odrv4
    port map (
            O => \N__28470\,
            I => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0\
        );

    \I__4950\ : CascadeMux
    port map (
            O => \N__28467\,
            I => \N__28464\
        );

    \I__4949\ : InMux
    port map (
            O => \N__28464\,
            I => \N__28461\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__28461\,
            I => \G_406\
        );

    \I__4947\ : CascadeMux
    port map (
            O => \N__28458\,
            I => \N__28454\
        );

    \I__4946\ : InMux
    port map (
            O => \N__28457\,
            I => \N__28447\
        );

    \I__4945\ : InMux
    port map (
            O => \N__28454\,
            I => \N__28444\
        );

    \I__4944\ : InMux
    port map (
            O => \N__28453\,
            I => \N__28435\
        );

    \I__4943\ : InMux
    port map (
            O => \N__28452\,
            I => \N__28435\
        );

    \I__4942\ : InMux
    port map (
            O => \N__28451\,
            I => \N__28435\
        );

    \I__4941\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28435\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__28447\,
            I => \N__28430\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__28444\,
            I => \N__28430\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__28435\,
            I => \current_shift_inst.elapsed_time_ns_phase_1\
        );

    \I__4937\ : Odrv4
    port map (
            O => \N__28430\,
            I => \current_shift_inst.elapsed_time_ns_phase_1\
        );

    \I__4936\ : CascadeMux
    port map (
            O => \N__28425\,
            I => \N__28422\
        );

    \I__4935\ : InMux
    port map (
            O => \N__28422\,
            I => \N__28419\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__28419\,
            I => \G_405\
        );

    \I__4933\ : InMux
    port map (
            O => \N__28416\,
            I => \N__28409\
        );

    \I__4932\ : InMux
    port map (
            O => \N__28415\,
            I => \N__28409\
        );

    \I__4931\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28406\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__28409\,
            I => \N__28403\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__28406\,
            I => \N__28400\
        );

    \I__4928\ : Span4Mux_h
    port map (
            O => \N__28403\,
            I => \N__28394\
        );

    \I__4927\ : Span4Mux_h
    port map (
            O => \N__28400\,
            I => \N__28394\
        );

    \I__4926\ : InMux
    port map (
            O => \N__28399\,
            I => \N__28391\
        );

    \I__4925\ : Odrv4
    port map (
            O => \N__28394\,
            I => \current_shift_inst.elapsed_time_ns_phase_14\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__28391\,
            I => \current_shift_inst.elapsed_time_ns_phase_14\
        );

    \I__4923\ : CascadeMux
    port map (
            O => \N__28386\,
            I => \N__28383\
        );

    \I__4922\ : InMux
    port map (
            O => \N__28383\,
            I => \N__28380\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__28380\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14\
        );

    \I__4920\ : InMux
    port map (
            O => \N__28377\,
            I => \N__28368\
        );

    \I__4919\ : InMux
    port map (
            O => \N__28376\,
            I => \N__28368\
        );

    \I__4918\ : InMux
    port map (
            O => \N__28375\,
            I => \N__28368\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__28368\,
            I => \N__28365\
        );

    \I__4916\ : Span4Mux_h
    port map (
            O => \N__28365\,
            I => \N__28361\
        );

    \I__4915\ : InMux
    port map (
            O => \N__28364\,
            I => \N__28358\
        );

    \I__4914\ : Odrv4
    port map (
            O => \N__28361\,
            I => \current_shift_inst.elapsed_time_ns_phase_16\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__28358\,
            I => \current_shift_inst.elapsed_time_ns_phase_16\
        );

    \I__4912\ : InMux
    port map (
            O => \N__28353\,
            I => \N__28350\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__28350\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIBU361_16\
        );

    \I__4910\ : InMux
    port map (
            O => \N__28347\,
            I => \N__28342\
        );

    \I__4909\ : InMux
    port map (
            O => \N__28346\,
            I => \N__28339\
        );

    \I__4908\ : InMux
    port map (
            O => \N__28345\,
            I => \N__28336\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__28342\,
            I => \N__28331\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__28339\,
            I => \N__28331\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__28336\,
            I => \N__28325\
        );

    \I__4904\ : Span4Mux_h
    port map (
            O => \N__28331\,
            I => \N__28325\
        );

    \I__4903\ : InMux
    port map (
            O => \N__28330\,
            I => \N__28322\
        );

    \I__4902\ : Span4Mux_v
    port map (
            O => \N__28325\,
            I => \N__28319\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__28322\,
            I => \N__28316\
        );

    \I__4900\ : Odrv4
    port map (
            O => \N__28319\,
            I => \current_shift_inst.elapsed_time_ns_phase_17\
        );

    \I__4899\ : Odrv4
    port map (
            O => \N__28316\,
            I => \current_shift_inst.elapsed_time_ns_phase_17\
        );

    \I__4898\ : CascadeMux
    port map (
            O => \N__28311\,
            I => \N__28308\
        );

    \I__4897\ : InMux
    port map (
            O => \N__28308\,
            I => \N__28305\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__28305\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17\
        );

    \I__4895\ : InMux
    port map (
            O => \N__28302\,
            I => \N__28297\
        );

    \I__4894\ : InMux
    port map (
            O => \N__28301\,
            I => \N__28294\
        );

    \I__4893\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28291\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__28297\,
            I => \N__28284\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__28294\,
            I => \N__28284\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__28291\,
            I => \N__28284\
        );

    \I__4889\ : Span4Mux_v
    port map (
            O => \N__28284\,
            I => \N__28281\
        );

    \I__4888\ : Span4Mux_v
    port map (
            O => \N__28281\,
            I => \N__28277\
        );

    \I__4887\ : InMux
    port map (
            O => \N__28280\,
            I => \N__28274\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__28277\,
            I => \current_shift_inst.elapsed_time_ns_phase_12\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__28274\,
            I => \current_shift_inst.elapsed_time_ns_phase_12\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__28269\,
            I => \N__28266\
        );

    \I__4883\ : InMux
    port map (
            O => \N__28266\,
            I => \N__28263\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__28263\,
            I => \N__28258\
        );

    \I__4881\ : InMux
    port map (
            O => \N__28262\,
            I => \N__28253\
        );

    \I__4880\ : InMux
    port map (
            O => \N__28261\,
            I => \N__28253\
        );

    \I__4879\ : Span4Mux_h
    port map (
            O => \N__28258\,
            I => \N__28248\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__28253\,
            I => \N__28248\
        );

    \I__4877\ : Span4Mux_h
    port map (
            O => \N__28248\,
            I => \N__28244\
        );

    \I__4876\ : InMux
    port map (
            O => \N__28247\,
            I => \N__28241\
        );

    \I__4875\ : Odrv4
    port map (
            O => \N__28244\,
            I => \current_shift_inst.elapsed_time_ns_phase_11\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__28241\,
            I => \current_shift_inst.elapsed_time_ns_phase_11\
        );

    \I__4873\ : InMux
    port map (
            O => \N__28236\,
            I => \N__28233\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__28233\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11\
        );

    \I__4871\ : CascadeMux
    port map (
            O => \N__28230\,
            I => \N__28227\
        );

    \I__4870\ : InMux
    port map (
            O => \N__28227\,
            I => \N__28224\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__28224\,
            I => \N__28221\
        );

    \I__4868\ : Span4Mux_v
    port map (
            O => \N__28221\,
            I => \N__28218\
        );

    \I__4867\ : Odrv4
    port map (
            O => \N__28218\,
            I => \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0\
        );

    \I__4866\ : CascadeMux
    port map (
            O => \N__28215\,
            I => \N__28212\
        );

    \I__4865\ : InMux
    port map (
            O => \N__28212\,
            I => \N__28209\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__28209\,
            I => \N__28206\
        );

    \I__4863\ : Odrv4
    port map (
            O => \N__28206\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIER9V_5\
        );

    \I__4862\ : InMux
    port map (
            O => \N__28203\,
            I => \N__28200\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__28200\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12\
        );

    \I__4860\ : InMux
    port map (
            O => \N__28197\,
            I => \N__28188\
        );

    \I__4859\ : InMux
    port map (
            O => \N__28196\,
            I => \N__28188\
        );

    \I__4858\ : InMux
    port map (
            O => \N__28195\,
            I => \N__28188\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__28188\,
            I => \N__28184\
        );

    \I__4856\ : CascadeMux
    port map (
            O => \N__28187\,
            I => \N__28181\
        );

    \I__4855\ : Span4Mux_h
    port map (
            O => \N__28184\,
            I => \N__28178\
        );

    \I__4854\ : InMux
    port map (
            O => \N__28181\,
            I => \N__28175\
        );

    \I__4853\ : Odrv4
    port map (
            O => \N__28178\,
            I => \current_shift_inst.elapsed_time_ns_phase_7\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__28175\,
            I => \current_shift_inst.elapsed_time_ns_phase_7\
        );

    \I__4851\ : InMux
    port map (
            O => \N__28170\,
            I => \N__28167\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__28167\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7\
        );

    \I__4849\ : CascadeMux
    port map (
            O => \N__28164\,
            I => \N__28161\
        );

    \I__4848\ : InMux
    port map (
            O => \N__28161\,
            I => \N__28154\
        );

    \I__4847\ : InMux
    port map (
            O => \N__28160\,
            I => \N__28154\
        );

    \I__4846\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28151\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__28154\,
            I => \N__28148\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__28151\,
            I => \N__28142\
        );

    \I__4843\ : Span4Mux_h
    port map (
            O => \N__28148\,
            I => \N__28142\
        );

    \I__4842\ : InMux
    port map (
            O => \N__28147\,
            I => \N__28139\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__28142\,
            I => \current_shift_inst.elapsed_time_ns_phase_8\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__28139\,
            I => \current_shift_inst.elapsed_time_ns_phase_8\
        );

    \I__4839\ : CascadeMux
    port map (
            O => \N__28134\,
            I => \N__28131\
        );

    \I__4838\ : InMux
    port map (
            O => \N__28131\,
            I => \N__28128\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__28128\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8\
        );

    \I__4836\ : InMux
    port map (
            O => \N__28125\,
            I => \N__28122\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__28122\,
            I => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0\
        );

    \I__4834\ : InMux
    port map (
            O => \N__28119\,
            I => \N__28116\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__28116\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5M161_15\
        );

    \I__4832\ : CascadeMux
    port map (
            O => \N__28113\,
            I => \N__28110\
        );

    \I__4831\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28107\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__28107\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI190J_15\
        );

    \I__4829\ : CascadeMux
    port map (
            O => \N__28104\,
            I => \N__28101\
        );

    \I__4828\ : InMux
    port map (
            O => \N__28101\,
            I => \N__28098\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__28098\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16\
        );

    \I__4826\ : InMux
    port map (
            O => \N__28095\,
            I => \N__28086\
        );

    \I__4825\ : InMux
    port map (
            O => \N__28094\,
            I => \N__28086\
        );

    \I__4824\ : InMux
    port map (
            O => \N__28093\,
            I => \N__28086\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__28086\,
            I => \N__28083\
        );

    \I__4822\ : Span4Mux_h
    port map (
            O => \N__28083\,
            I => \N__28079\
        );

    \I__4821\ : InMux
    port map (
            O => \N__28082\,
            I => \N__28076\
        );

    \I__4820\ : Odrv4
    port map (
            O => \N__28079\,
            I => \current_shift_inst.elapsed_time_ns_phase_15\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__28076\,
            I => \current_shift_inst.elapsed_time_ns_phase_15\
        );

    \I__4818\ : InMux
    port map (
            O => \N__28071\,
            I => \N__28068\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__28068\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14\
        );

    \I__4816\ : CascadeMux
    port map (
            O => \N__28065\,
            I => \N__28062\
        );

    \I__4815\ : InMux
    port map (
            O => \N__28062\,
            I => \N__28059\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__28059\,
            I => \N__28056\
        );

    \I__4813\ : Odrv4
    port map (
            O => \N__28056\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12\
        );

    \I__4812\ : CascadeMux
    port map (
            O => \N__28053\,
            I => \N__28050\
        );

    \I__4811\ : InMux
    port map (
            O => \N__28050\,
            I => \N__28043\
        );

    \I__4810\ : InMux
    port map (
            O => \N__28049\,
            I => \N__28043\
        );

    \I__4809\ : InMux
    port map (
            O => \N__28048\,
            I => \N__28040\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__28043\,
            I => \N__28037\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__28040\,
            I => \N__28032\
        );

    \I__4806\ : Span4Mux_h
    port map (
            O => \N__28037\,
            I => \N__28032\
        );

    \I__4805\ : Sp12to4
    port map (
            O => \N__28032\,
            I => \N__28028\
        );

    \I__4804\ : InMux
    port map (
            O => \N__28031\,
            I => \N__28025\
        );

    \I__4803\ : Odrv12
    port map (
            O => \N__28028\,
            I => \current_shift_inst.elapsed_time_ns_phase_13\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__28025\,
            I => \current_shift_inst.elapsed_time_ns_phase_13\
        );

    \I__4801\ : InMux
    port map (
            O => \N__28020\,
            I => \N__28017\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__28017\,
            I => \N__28014\
        );

    \I__4799\ : Odrv4
    port map (
            O => \N__28014\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13\
        );

    \I__4798\ : InMux
    port map (
            O => \N__28011\,
            I => \N__28008\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__28008\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6\
        );

    \I__4796\ : CascadeMux
    port map (
            O => \N__28005\,
            I => \N__28002\
        );

    \I__4795\ : InMux
    port map (
            O => \N__28002\,
            I => \N__27999\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__27999\,
            I => \N__27996\
        );

    \I__4793\ : Odrv4
    port map (
            O => \N__27996\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6\
        );

    \I__4792\ : CascadeMux
    port map (
            O => \N__27993\,
            I => \N__27990\
        );

    \I__4791\ : InMux
    port map (
            O => \N__27990\,
            I => \N__27987\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__27987\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7\
        );

    \I__4789\ : CascadeMux
    port map (
            O => \N__27984\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_5_cascade_\
        );

    \I__4788\ : CascadeMux
    port map (
            O => \N__27981\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13_cascade_\
        );

    \I__4787\ : InMux
    port map (
            O => \N__27978\,
            I => \N__27975\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__27975\,
            I => \N__27972\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__27972\,
            I => \il_min_comp1_D1\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__27969\,
            I => \N__27966\
        );

    \I__4783\ : InMux
    port map (
            O => \N__27966\,
            I => \N__27961\
        );

    \I__4782\ : InMux
    port map (
            O => \N__27965\,
            I => \N__27956\
        );

    \I__4781\ : InMux
    port map (
            O => \N__27964\,
            I => \N__27956\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__27961\,
            I => measured_delay_hc_22
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__27956\,
            I => measured_delay_hc_22
        );

    \I__4778\ : CascadeMux
    port map (
            O => \N__27951\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_2_cascade_\
        );

    \I__4777\ : InMux
    port map (
            O => \N__27948\,
            I => \current_shift_inst.z_5_cry_25\
        );

    \I__4776\ : CascadeMux
    port map (
            O => \N__27945\,
            I => \N__27941\
        );

    \I__4775\ : InMux
    port map (
            O => \N__27944\,
            I => \N__27933\
        );

    \I__4774\ : InMux
    port map (
            O => \N__27941\,
            I => \N__27933\
        );

    \I__4773\ : InMux
    port map (
            O => \N__27940\,
            I => \N__27933\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__27933\,
            I => \N__27930\
        );

    \I__4771\ : Span4Mux_h
    port map (
            O => \N__27930\,
            I => \N__27926\
        );

    \I__4770\ : InMux
    port map (
            O => \N__27929\,
            I => \N__27923\
        );

    \I__4769\ : Odrv4
    port map (
            O => \N__27926\,
            I => \current_shift_inst.elapsed_time_ns_phase_27\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__27923\,
            I => \current_shift_inst.elapsed_time_ns_phase_27\
        );

    \I__4767\ : InMux
    port map (
            O => \N__27918\,
            I => \current_shift_inst.z_5_cry_26\
        );

    \I__4766\ : InMux
    port map (
            O => \N__27915\,
            I => \N__27906\
        );

    \I__4765\ : InMux
    port map (
            O => \N__27914\,
            I => \N__27906\
        );

    \I__4764\ : InMux
    port map (
            O => \N__27913\,
            I => \N__27906\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__27906\,
            I => \N__27903\
        );

    \I__4762\ : Span4Mux_h
    port map (
            O => \N__27903\,
            I => \N__27899\
        );

    \I__4761\ : InMux
    port map (
            O => \N__27902\,
            I => \N__27896\
        );

    \I__4760\ : Odrv4
    port map (
            O => \N__27899\,
            I => \current_shift_inst.elapsed_time_ns_phase_28\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__27896\,
            I => \current_shift_inst.elapsed_time_ns_phase_28\
        );

    \I__4758\ : InMux
    port map (
            O => \N__27891\,
            I => \current_shift_inst.z_5_cry_27\
        );

    \I__4757\ : CascadeMux
    port map (
            O => \N__27888\,
            I => \N__27884\
        );

    \I__4756\ : InMux
    port map (
            O => \N__27887\,
            I => \N__27879\
        );

    \I__4755\ : InMux
    port map (
            O => \N__27884\,
            I => \N__27879\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__27879\,
            I => \N__27876\
        );

    \I__4753\ : Span4Mux_h
    port map (
            O => \N__27876\,
            I => \N__27872\
        );

    \I__4752\ : InMux
    port map (
            O => \N__27875\,
            I => \N__27869\
        );

    \I__4751\ : Odrv4
    port map (
            O => \N__27872\,
            I => \current_shift_inst.elapsed_time_ns_phase_29\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__27869\,
            I => \current_shift_inst.elapsed_time_ns_phase_29\
        );

    \I__4749\ : InMux
    port map (
            O => \N__27864\,
            I => \current_shift_inst.z_5_cry_28\
        );

    \I__4748\ : CascadeMux
    port map (
            O => \N__27861\,
            I => \N__27854\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__27860\,
            I => \N__27851\
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__27859\,
            I => \N__27848\
        );

    \I__4745\ : CascadeMux
    port map (
            O => \N__27858\,
            I => \N__27845\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__27857\,
            I => \N__27842\
        );

    \I__4743\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27823\
        );

    \I__4742\ : InMux
    port map (
            O => \N__27851\,
            I => \N__27814\
        );

    \I__4741\ : InMux
    port map (
            O => \N__27848\,
            I => \N__27814\
        );

    \I__4740\ : InMux
    port map (
            O => \N__27845\,
            I => \N__27814\
        );

    \I__4739\ : InMux
    port map (
            O => \N__27842\,
            I => \N__27814\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__27841\,
            I => \N__27811\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__27840\,
            I => \N__27808\
        );

    \I__4736\ : CascadeMux
    port map (
            O => \N__27839\,
            I => \N__27805\
        );

    \I__4735\ : CascadeMux
    port map (
            O => \N__27838\,
            I => \N__27802\
        );

    \I__4734\ : InMux
    port map (
            O => \N__27837\,
            I => \N__27791\
        );

    \I__4733\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27791\
        );

    \I__4732\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27791\
        );

    \I__4731\ : InMux
    port map (
            O => \N__27834\,
            I => \N__27788\
        );

    \I__4730\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27779\
        );

    \I__4729\ : InMux
    port map (
            O => \N__27832\,
            I => \N__27779\
        );

    \I__4728\ : InMux
    port map (
            O => \N__27831\,
            I => \N__27779\
        );

    \I__4727\ : InMux
    port map (
            O => \N__27830\,
            I => \N__27779\
        );

    \I__4726\ : CascadeMux
    port map (
            O => \N__27829\,
            I => \N__27769\
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__27828\,
            I => \N__27766\
        );

    \I__4724\ : CascadeMux
    port map (
            O => \N__27827\,
            I => \N__27763\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__27826\,
            I => \N__27760\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__27823\,
            I => \N__27755\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__27814\,
            I => \N__27755\
        );

    \I__4720\ : InMux
    port map (
            O => \N__27811\,
            I => \N__27746\
        );

    \I__4719\ : InMux
    port map (
            O => \N__27808\,
            I => \N__27746\
        );

    \I__4718\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27746\
        );

    \I__4717\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27746\
        );

    \I__4716\ : CascadeMux
    port map (
            O => \N__27801\,
            I => \N__27743\
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__27800\,
            I => \N__27740\
        );

    \I__4714\ : CascadeMux
    port map (
            O => \N__27799\,
            I => \N__27737\
        );

    \I__4713\ : CascadeMux
    port map (
            O => \N__27798\,
            I => \N__27734\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__27791\,
            I => \N__27731\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__27788\,
            I => \N__27726\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__27779\,
            I => \N__27726\
        );

    \I__4709\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27723\
        );

    \I__4708\ : CascadeMux
    port map (
            O => \N__27777\,
            I => \N__27720\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__27776\,
            I => \N__27717\
        );

    \I__4706\ : CascadeMux
    port map (
            O => \N__27775\,
            I => \N__27706\
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__27774\,
            I => \N__27702\
        );

    \I__4704\ : CascadeMux
    port map (
            O => \N__27773\,
            I => \N__27699\
        );

    \I__4703\ : CascadeMux
    port map (
            O => \N__27772\,
            I => \N__27695\
        );

    \I__4702\ : InMux
    port map (
            O => \N__27769\,
            I => \N__27686\
        );

    \I__4701\ : InMux
    port map (
            O => \N__27766\,
            I => \N__27686\
        );

    \I__4700\ : InMux
    port map (
            O => \N__27763\,
            I => \N__27686\
        );

    \I__4699\ : InMux
    port map (
            O => \N__27760\,
            I => \N__27686\
        );

    \I__4698\ : Span4Mux_v
    port map (
            O => \N__27755\,
            I => \N__27681\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__27746\,
            I => \N__27681\
        );

    \I__4696\ : InMux
    port map (
            O => \N__27743\,
            I => \N__27672\
        );

    \I__4695\ : InMux
    port map (
            O => \N__27740\,
            I => \N__27672\
        );

    \I__4694\ : InMux
    port map (
            O => \N__27737\,
            I => \N__27672\
        );

    \I__4693\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27672\
        );

    \I__4692\ : Span4Mux_v
    port map (
            O => \N__27731\,
            I => \N__27659\
        );

    \I__4691\ : Span4Mux_v
    port map (
            O => \N__27726\,
            I => \N__27659\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__27723\,
            I => \N__27659\
        );

    \I__4689\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27656\
        );

    \I__4688\ : InMux
    port map (
            O => \N__27717\,
            I => \N__27651\
        );

    \I__4687\ : InMux
    port map (
            O => \N__27716\,
            I => \N__27651\
        );

    \I__4686\ : InMux
    port map (
            O => \N__27715\,
            I => \N__27644\
        );

    \I__4685\ : InMux
    port map (
            O => \N__27714\,
            I => \N__27644\
        );

    \I__4684\ : InMux
    port map (
            O => \N__27713\,
            I => \N__27644\
        );

    \I__4683\ : InMux
    port map (
            O => \N__27712\,
            I => \N__27635\
        );

    \I__4682\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27635\
        );

    \I__4681\ : InMux
    port map (
            O => \N__27710\,
            I => \N__27635\
        );

    \I__4680\ : InMux
    port map (
            O => \N__27709\,
            I => \N__27635\
        );

    \I__4679\ : InMux
    port map (
            O => \N__27706\,
            I => \N__27622\
        );

    \I__4678\ : InMux
    port map (
            O => \N__27705\,
            I => \N__27622\
        );

    \I__4677\ : InMux
    port map (
            O => \N__27702\,
            I => \N__27622\
        );

    \I__4676\ : InMux
    port map (
            O => \N__27699\,
            I => \N__27622\
        );

    \I__4675\ : InMux
    port map (
            O => \N__27698\,
            I => \N__27622\
        );

    \I__4674\ : InMux
    port map (
            O => \N__27695\,
            I => \N__27622\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__27686\,
            I => \N__27619\
        );

    \I__4672\ : Span4Mux_h
    port map (
            O => \N__27681\,
            I => \N__27614\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__27672\,
            I => \N__27614\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__27671\,
            I => \N__27611\
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__27670\,
            I => \N__27608\
        );

    \I__4668\ : CascadeMux
    port map (
            O => \N__27669\,
            I => \N__27605\
        );

    \I__4667\ : CascadeMux
    port map (
            O => \N__27668\,
            I => \N__27602\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__27667\,
            I => \N__27599\
        );

    \I__4665\ : CascadeMux
    port map (
            O => \N__27666\,
            I => \N__27596\
        );

    \I__4664\ : Span4Mux_v
    port map (
            O => \N__27659\,
            I => \N__27592\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__27656\,
            I => \N__27587\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__27651\,
            I => \N__27587\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__27644\,
            I => \N__27582\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__27635\,
            I => \N__27582\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__27622\,
            I => \N__27579\
        );

    \I__4658\ : Span4Mux_v
    port map (
            O => \N__27619\,
            I => \N__27574\
        );

    \I__4657\ : Span4Mux_v
    port map (
            O => \N__27614\,
            I => \N__27574\
        );

    \I__4656\ : InMux
    port map (
            O => \N__27611\,
            I => \N__27567\
        );

    \I__4655\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27567\
        );

    \I__4654\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27567\
        );

    \I__4653\ : InMux
    port map (
            O => \N__27602\,
            I => \N__27560\
        );

    \I__4652\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27560\
        );

    \I__4651\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27560\
        );

    \I__4650\ : InMux
    port map (
            O => \N__27595\,
            I => \N__27557\
        );

    \I__4649\ : Sp12to4
    port map (
            O => \N__27592\,
            I => \N__27553\
        );

    \I__4648\ : Span4Mux_v
    port map (
            O => \N__27587\,
            I => \N__27548\
        );

    \I__4647\ : Span4Mux_s2_h
    port map (
            O => \N__27582\,
            I => \N__27548\
        );

    \I__4646\ : Span4Mux_v
    port map (
            O => \N__27579\,
            I => \N__27539\
        );

    \I__4645\ : Span4Mux_v
    port map (
            O => \N__27574\,
            I => \N__27539\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__27567\,
            I => \N__27539\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__27560\,
            I => \N__27539\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__27557\,
            I => \N__27536\
        );

    \I__4641\ : InMux
    port map (
            O => \N__27556\,
            I => \N__27532\
        );

    \I__4640\ : Span12Mux_h
    port map (
            O => \N__27553\,
            I => \N__27526\
        );

    \I__4639\ : Sp12to4
    port map (
            O => \N__27548\,
            I => \N__27526\
        );

    \I__4638\ : Sp12to4
    port map (
            O => \N__27539\,
            I => \N__27523\
        );

    \I__4637\ : Span12Mux_s3_h
    port map (
            O => \N__27536\,
            I => \N__27520\
        );

    \I__4636\ : InMux
    port map (
            O => \N__27535\,
            I => \N__27517\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__27532\,
            I => \N__27514\
        );

    \I__4634\ : InMux
    port map (
            O => \N__27531\,
            I => \N__27511\
        );

    \I__4633\ : Span12Mux_v
    port map (
            O => \N__27526\,
            I => \N__27508\
        );

    \I__4632\ : Span12Mux_v
    port map (
            O => \N__27523\,
            I => \N__27501\
        );

    \I__4631\ : Span12Mux_h
    port map (
            O => \N__27520\,
            I => \N__27501\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__27517\,
            I => \N__27501\
        );

    \I__4629\ : Span4Mux_s1_v
    port map (
            O => \N__27514\,
            I => \N__27496\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__27511\,
            I => \N__27496\
        );

    \I__4627\ : Odrv12
    port map (
            O => \N__27508\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4626\ : Odrv12
    port map (
            O => \N__27501\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4625\ : Odrv4
    port map (
            O => \N__27496\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4624\ : InMux
    port map (
            O => \N__27489\,
            I => \current_shift_inst.z_5_cry_29\
        );

    \I__4623\ : InMux
    port map (
            O => \N__27486\,
            I => \current_shift_inst.z_5_cry_30\
        );

    \I__4622\ : InMux
    port map (
            O => \N__27483\,
            I => \N__27480\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__27480\,
            I => \N__27477\
        );

    \I__4620\ : Span4Mux_h
    port map (
            O => \N__27477\,
            I => \N__27474\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__27474\,
            I => \il_min_comp2_D1\
        );

    \I__4618\ : InMux
    port map (
            O => \N__27471\,
            I => \N__27468\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__27468\,
            I => \N__27462\
        );

    \I__4616\ : InMux
    port map (
            O => \N__27467\,
            I => \N__27457\
        );

    \I__4615\ : InMux
    port map (
            O => \N__27466\,
            I => \N__27457\
        );

    \I__4614\ : InMux
    port map (
            O => \N__27465\,
            I => \N__27454\
        );

    \I__4613\ : Span4Mux_h
    port map (
            O => \N__27462\,
            I => \N__27449\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__27457\,
            I => \N__27449\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__27454\,
            I => \N__27446\
        );

    \I__4610\ : Odrv4
    port map (
            O => \N__27449\,
            I => \current_shift_inst.elapsed_time_ns_phase_18\
        );

    \I__4609\ : Odrv4
    port map (
            O => \N__27446\,
            I => \current_shift_inst.elapsed_time_ns_phase_18\
        );

    \I__4608\ : InMux
    port map (
            O => \N__27441\,
            I => \current_shift_inst.z_5_cry_17\
        );

    \I__4607\ : CascadeMux
    port map (
            O => \N__27438\,
            I => \N__27434\
        );

    \I__4606\ : InMux
    port map (
            O => \N__27437\,
            I => \N__27426\
        );

    \I__4605\ : InMux
    port map (
            O => \N__27434\,
            I => \N__27426\
        );

    \I__4604\ : InMux
    port map (
            O => \N__27433\,
            I => \N__27426\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__27426\,
            I => \N__27423\
        );

    \I__4602\ : Span4Mux_h
    port map (
            O => \N__27423\,
            I => \N__27419\
        );

    \I__4601\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27416\
        );

    \I__4600\ : Odrv4
    port map (
            O => \N__27419\,
            I => \current_shift_inst.elapsed_time_ns_phase_19\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__27416\,
            I => \current_shift_inst.elapsed_time_ns_phase_19\
        );

    \I__4598\ : InMux
    port map (
            O => \N__27411\,
            I => \current_shift_inst.z_5_cry_18\
        );

    \I__4597\ : InMux
    port map (
            O => \N__27408\,
            I => \N__27399\
        );

    \I__4596\ : InMux
    port map (
            O => \N__27407\,
            I => \N__27399\
        );

    \I__4595\ : InMux
    port map (
            O => \N__27406\,
            I => \N__27399\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__27399\,
            I => \N__27396\
        );

    \I__4593\ : Span4Mux_h
    port map (
            O => \N__27396\,
            I => \N__27392\
        );

    \I__4592\ : InMux
    port map (
            O => \N__27395\,
            I => \N__27389\
        );

    \I__4591\ : Odrv4
    port map (
            O => \N__27392\,
            I => \current_shift_inst.elapsed_time_ns_phase_20\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__27389\,
            I => \current_shift_inst.elapsed_time_ns_phase_20\
        );

    \I__4589\ : InMux
    port map (
            O => \N__27384\,
            I => \current_shift_inst.z_5_cry_19\
        );

    \I__4588\ : CascadeMux
    port map (
            O => \N__27381\,
            I => \N__27376\
        );

    \I__4587\ : InMux
    port map (
            O => \N__27380\,
            I => \N__27373\
        );

    \I__4586\ : InMux
    port map (
            O => \N__27379\,
            I => \N__27368\
        );

    \I__4585\ : InMux
    port map (
            O => \N__27376\,
            I => \N__27368\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__27373\,
            I => \N__27363\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__27368\,
            I => \N__27363\
        );

    \I__4582\ : Span4Mux_h
    port map (
            O => \N__27363\,
            I => \N__27359\
        );

    \I__4581\ : InMux
    port map (
            O => \N__27362\,
            I => \N__27356\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__27359\,
            I => \current_shift_inst.elapsed_time_ns_phase_21\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__27356\,
            I => \current_shift_inst.elapsed_time_ns_phase_21\
        );

    \I__4578\ : InMux
    port map (
            O => \N__27351\,
            I => \current_shift_inst.z_5_cry_20\
        );

    \I__4577\ : InMux
    port map (
            O => \N__27348\,
            I => \current_shift_inst.z_5_cry_21\
        );

    \I__4576\ : InMux
    port map (
            O => \N__27345\,
            I => \current_shift_inst.z_5_cry_22\
        );

    \I__4575\ : InMux
    port map (
            O => \N__27342\,
            I => \current_shift_inst.z_5_cry_23\
        );

    \I__4574\ : InMux
    port map (
            O => \N__27339\,
            I => \bfn_9_21_0_\
        );

    \I__4573\ : InMux
    port map (
            O => \N__27336\,
            I => \N__27327\
        );

    \I__4572\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27327\
        );

    \I__4571\ : InMux
    port map (
            O => \N__27334\,
            I => \N__27327\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__27327\,
            I => \N__27323\
        );

    \I__4569\ : InMux
    port map (
            O => \N__27326\,
            I => \N__27320\
        );

    \I__4568\ : Span4Mux_h
    port map (
            O => \N__27323\,
            I => \N__27317\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__27320\,
            I => \N__27314\
        );

    \I__4566\ : Odrv4
    port map (
            O => \N__27317\,
            I => \current_shift_inst.elapsed_time_ns_phase_9\
        );

    \I__4565\ : Odrv4
    port map (
            O => \N__27314\,
            I => \current_shift_inst.elapsed_time_ns_phase_9\
        );

    \I__4564\ : InMux
    port map (
            O => \N__27309\,
            I => \bfn_9_19_0_\
        );

    \I__4563\ : InMux
    port map (
            O => \N__27306\,
            I => \N__27297\
        );

    \I__4562\ : InMux
    port map (
            O => \N__27305\,
            I => \N__27297\
        );

    \I__4561\ : InMux
    port map (
            O => \N__27304\,
            I => \N__27297\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__27297\,
            I => \N__27293\
        );

    \I__4559\ : InMux
    port map (
            O => \N__27296\,
            I => \N__27290\
        );

    \I__4558\ : Span4Mux_h
    port map (
            O => \N__27293\,
            I => \N__27287\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__27290\,
            I => \N__27284\
        );

    \I__4556\ : Odrv4
    port map (
            O => \N__27287\,
            I => \current_shift_inst.elapsed_time_ns_phase_10\
        );

    \I__4555\ : Odrv4
    port map (
            O => \N__27284\,
            I => \current_shift_inst.elapsed_time_ns_phase_10\
        );

    \I__4554\ : InMux
    port map (
            O => \N__27279\,
            I => \current_shift_inst.z_5_cry_9\
        );

    \I__4553\ : InMux
    port map (
            O => \N__27276\,
            I => \current_shift_inst.z_5_cry_10\
        );

    \I__4552\ : InMux
    port map (
            O => \N__27273\,
            I => \current_shift_inst.z_5_cry_11\
        );

    \I__4551\ : InMux
    port map (
            O => \N__27270\,
            I => \current_shift_inst.z_5_cry_12\
        );

    \I__4550\ : InMux
    port map (
            O => \N__27267\,
            I => \current_shift_inst.z_5_cry_13\
        );

    \I__4549\ : InMux
    port map (
            O => \N__27264\,
            I => \current_shift_inst.z_5_cry_14\
        );

    \I__4548\ : InMux
    port map (
            O => \N__27261\,
            I => \current_shift_inst.z_5_cry_15\
        );

    \I__4547\ : InMux
    port map (
            O => \N__27258\,
            I => \bfn_9_20_0_\
        );

    \I__4546\ : CascadeMux
    port map (
            O => \N__27255\,
            I => \N__27252\
        );

    \I__4545\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27249\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__27249\,
            I => \current_shift_inst.control_input_1_cry_24_THRU_CO\
        );

    \I__4543\ : InMux
    port map (
            O => \N__27246\,
            I => \bfn_9_17_0_\
        );

    \I__4542\ : CascadeMux
    port map (
            O => \N__27243\,
            I => \N__27240\
        );

    \I__4541\ : InMux
    port map (
            O => \N__27240\,
            I => \N__27234\
        );

    \I__4540\ : CascadeMux
    port map (
            O => \N__27239\,
            I => \N__27229\
        );

    \I__4539\ : CascadeMux
    port map (
            O => \N__27238\,
            I => \N__27226\
        );

    \I__4538\ : CascadeMux
    port map (
            O => \N__27237\,
            I => \N__27222\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__27234\,
            I => \N__27218\
        );

    \I__4536\ : InMux
    port map (
            O => \N__27233\,
            I => \N__27215\
        );

    \I__4535\ : InMux
    port map (
            O => \N__27232\,
            I => \N__27202\
        );

    \I__4534\ : InMux
    port map (
            O => \N__27229\,
            I => \N__27202\
        );

    \I__4533\ : InMux
    port map (
            O => \N__27226\,
            I => \N__27202\
        );

    \I__4532\ : InMux
    port map (
            O => \N__27225\,
            I => \N__27202\
        );

    \I__4531\ : InMux
    port map (
            O => \N__27222\,
            I => \N__27202\
        );

    \I__4530\ : InMux
    port map (
            O => \N__27221\,
            I => \N__27202\
        );

    \I__4529\ : Span4Mux_h
    port map (
            O => \N__27218\,
            I => \N__27199\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__27215\,
            I => \N__27194\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__27202\,
            I => \N__27194\
        );

    \I__4526\ : Span4Mux_h
    port map (
            O => \N__27199\,
            I => \N__27189\
        );

    \I__4525\ : Span4Mux_h
    port map (
            O => \N__27194\,
            I => \N__27189\
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__27189\,
            I => \current_shift_inst.control_inputZ0Z_25\
        );

    \I__4523\ : CEMux
    port map (
            O => \N__27186\,
            I => \N__27181\
        );

    \I__4522\ : CEMux
    port map (
            O => \N__27185\,
            I => \N__27178\
        );

    \I__4521\ : CEMux
    port map (
            O => \N__27184\,
            I => \N__27175\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__27181\,
            I => \N__27171\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__27178\,
            I => \N__27166\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__27175\,
            I => \N__27166\
        );

    \I__4517\ : CEMux
    port map (
            O => \N__27174\,
            I => \N__27163\
        );

    \I__4516\ : Span4Mux_v
    port map (
            O => \N__27171\,
            I => \N__27155\
        );

    \I__4515\ : Span4Mux_v
    port map (
            O => \N__27166\,
            I => \N__27155\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__27163\,
            I => \N__27155\
        );

    \I__4513\ : CEMux
    port map (
            O => \N__27162\,
            I => \N__27152\
        );

    \I__4512\ : Span4Mux_v
    port map (
            O => \N__27155\,
            I => \N__27149\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__27152\,
            I => \N__27146\
        );

    \I__4510\ : Span4Mux_v
    port map (
            O => \N__27149\,
            I => \N__27143\
        );

    \I__4509\ : Span4Mux_v
    port map (
            O => \N__27146\,
            I => \N__27140\
        );

    \I__4508\ : Odrv4
    port map (
            O => \N__27143\,
            I => \current_shift_inst.phase_valid_RNISLORZ0Z2\
        );

    \I__4507\ : Odrv4
    port map (
            O => \N__27140\,
            I => \current_shift_inst.phase_valid_RNISLORZ0Z2\
        );

    \I__4506\ : InMux
    port map (
            O => \N__27135\,
            I => \current_shift_inst.z_5_cry_1\
        );

    \I__4505\ : InMux
    port map (
            O => \N__27132\,
            I => \current_shift_inst.z_5_cry_2\
        );

    \I__4504\ : InMux
    port map (
            O => \N__27129\,
            I => \current_shift_inst.z_5_cry_3\
        );

    \I__4503\ : InMux
    port map (
            O => \N__27126\,
            I => \current_shift_inst.z_5_cry_4\
        );

    \I__4502\ : InMux
    port map (
            O => \N__27123\,
            I => \current_shift_inst.z_5_cry_5\
        );

    \I__4501\ : InMux
    port map (
            O => \N__27120\,
            I => \current_shift_inst.z_5_cry_6\
        );

    \I__4500\ : InMux
    port map (
            O => \N__27117\,
            I => \current_shift_inst.z_5_cry_7\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__27114\,
            I => \N__27111\
        );

    \I__4498\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27108\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__27108\,
            I => \N__27105\
        );

    \I__4496\ : Span4Mux_h
    port map (
            O => \N__27105\,
            I => \N__27102\
        );

    \I__4495\ : Odrv4
    port map (
            O => \N__27102\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIR32K_22\
        );

    \I__4494\ : InMux
    port map (
            O => \N__27099\,
            I => \N__27096\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__27096\,
            I => \current_shift_inst.control_input_1_axb_17\
        );

    \I__4492\ : InMux
    port map (
            O => \N__27093\,
            I => \bfn_9_16_0_\
        );

    \I__4491\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27087\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__27087\,
            I => \current_shift_inst.control_input_1_axb_18\
        );

    \I__4489\ : InMux
    port map (
            O => \N__27084\,
            I => \current_shift_inst.un38_control_input_0_cry_23\
        );

    \I__4488\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27078\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__27078\,
            I => \current_shift_inst.control_input_1_axb_19\
        );

    \I__4486\ : InMux
    port map (
            O => \N__27075\,
            I => \current_shift_inst.un38_control_input_0_cry_24\
        );

    \I__4485\ : InMux
    port map (
            O => \N__27072\,
            I => \N__27069\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__27069\,
            I => \current_shift_inst.control_input_1_axb_20\
        );

    \I__4483\ : InMux
    port map (
            O => \N__27066\,
            I => \current_shift_inst.un38_control_input_0_cry_25\
        );

    \I__4482\ : InMux
    port map (
            O => \N__27063\,
            I => \N__27060\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__27060\,
            I => \N__27057\
        );

    \I__4480\ : Odrv4
    port map (
            O => \N__27057\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26\
        );

    \I__4479\ : InMux
    port map (
            O => \N__27054\,
            I => \N__27051\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__27051\,
            I => \current_shift_inst.control_input_1_axb_21\
        );

    \I__4477\ : InMux
    port map (
            O => \N__27048\,
            I => \current_shift_inst.un38_control_input_0_cry_26\
        );

    \I__4476\ : InMux
    port map (
            O => \N__27045\,
            I => \N__27042\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__27042\,
            I => \N__27039\
        );

    \I__4474\ : Odrv4
    port map (
            O => \N__27039\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINKG81_27\
        );

    \I__4473\ : CascadeMux
    port map (
            O => \N__27036\,
            I => \N__27033\
        );

    \I__4472\ : InMux
    port map (
            O => \N__27033\,
            I => \N__27030\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__27030\,
            I => \N__27027\
        );

    \I__4470\ : Odrv4
    port map (
            O => \N__27027\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27\
        );

    \I__4469\ : InMux
    port map (
            O => \N__27024\,
            I => \N__27021\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__27021\,
            I => \current_shift_inst.control_input_1_axb_22\
        );

    \I__4467\ : InMux
    port map (
            O => \N__27018\,
            I => \current_shift_inst.un38_control_input_0_cry_27\
        );

    \I__4466\ : InMux
    port map (
            O => \N__27015\,
            I => \N__27012\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__27012\,
            I => \N__27009\
        );

    \I__4464\ : Odrv12
    port map (
            O => \N__27009\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29\
        );

    \I__4463\ : CascadeMux
    port map (
            O => \N__27006\,
            I => \N__27003\
        );

    \I__4462\ : InMux
    port map (
            O => \N__27003\,
            I => \N__27000\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__27000\,
            I => \N__26997\
        );

    \I__4460\ : Odrv12
    port map (
            O => \N__26997\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28\
        );

    \I__4459\ : InMux
    port map (
            O => \N__26994\,
            I => \N__26991\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__26991\,
            I => \current_shift_inst.control_input_1_axb_23\
        );

    \I__4457\ : InMux
    port map (
            O => \N__26988\,
            I => \current_shift_inst.un38_control_input_0_cry_28\
        );

    \I__4456\ : InMux
    port map (
            O => \N__26985\,
            I => \N__26982\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__26982\,
            I => \N__26979\
        );

    \I__4454\ : Span4Mux_h
    port map (
            O => \N__26979\,
            I => \N__26976\
        );

    \I__4453\ : Odrv4
    port map (
            O => \N__26976\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30\
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__26973\,
            I => \N__26970\
        );

    \I__4451\ : InMux
    port map (
            O => \N__26970\,
            I => \N__26966\
        );

    \I__4450\ : InMux
    port map (
            O => \N__26969\,
            I => \N__26963\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__26966\,
            I => \N__26960\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__26963\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\
        );

    \I__4447\ : Odrv12
    port map (
            O => \N__26960\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\
        );

    \I__4446\ : InMux
    port map (
            O => \N__26955\,
            I => \N__26952\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__26952\,
            I => \current_shift_inst.control_input_1_axb_24\
        );

    \I__4444\ : InMux
    port map (
            O => \N__26949\,
            I => \current_shift_inst.un38_control_input_0_cry_29\
        );

    \I__4443\ : InMux
    port map (
            O => \N__26946\,
            I => \N__26943\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__26943\,
            I => \current_shift_inst.control_input_1_axb_9\
        );

    \I__4441\ : InMux
    port map (
            O => \N__26940\,
            I => \bfn_9_15_0_\
        );

    \I__4440\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26934\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__26934\,
            I => \current_shift_inst.control_input_1_axb_10\
        );

    \I__4438\ : InMux
    port map (
            O => \N__26931\,
            I => \current_shift_inst.un38_control_input_0_cry_15\
        );

    \I__4437\ : InMux
    port map (
            O => \N__26928\,
            I => \N__26925\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__26925\,
            I => \current_shift_inst.control_input_1_axb_11\
        );

    \I__4435\ : InMux
    port map (
            O => \N__26922\,
            I => \current_shift_inst.un38_control_input_0_cry_16\
        );

    \I__4434\ : InMux
    port map (
            O => \N__26919\,
            I => \N__26916\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__26916\,
            I => \N__26913\
        );

    \I__4432\ : Span4Mux_v
    port map (
            O => \N__26913\,
            I => \N__26910\
        );

    \I__4431\ : Odrv4
    port map (
            O => \N__26910\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIH6661_17\
        );

    \I__4430\ : InMux
    port map (
            O => \N__26907\,
            I => \N__26904\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__26904\,
            I => \current_shift_inst.control_input_1_axb_12\
        );

    \I__4428\ : InMux
    port map (
            O => \N__26901\,
            I => \current_shift_inst.un38_control_input_0_cry_17\
        );

    \I__4427\ : InMux
    port map (
            O => \N__26898\,
            I => \N__26895\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__26895\,
            I => \N__26892\
        );

    \I__4425\ : Odrv4
    port map (
            O => \N__26892\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIE6961_18\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__26889\,
            I => \N__26886\
        );

    \I__4423\ : InMux
    port map (
            O => \N__26886\,
            I => \N__26883\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__26883\,
            I => \N__26880\
        );

    \I__4421\ : Span4Mux_v
    port map (
            O => \N__26880\,
            I => \N__26877\
        );

    \I__4420\ : Odrv4
    port map (
            O => \N__26877\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18\
        );

    \I__4419\ : InMux
    port map (
            O => \N__26874\,
            I => \N__26871\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__26871\,
            I => \current_shift_inst.control_input_1_axb_13\
        );

    \I__4417\ : InMux
    port map (
            O => \N__26868\,
            I => \current_shift_inst.un38_control_input_0_cry_18\
        );

    \I__4416\ : InMux
    port map (
            O => \N__26865\,
            I => \N__26862\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__26862\,
            I => \N__26859\
        );

    \I__4414\ : Odrv4
    port map (
            O => \N__26859\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPC571_19\
        );

    \I__4413\ : CascadeMux
    port map (
            O => \N__26856\,
            I => \N__26853\
        );

    \I__4412\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26850\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__26850\,
            I => \N__26847\
        );

    \I__4410\ : Odrv12
    port map (
            O => \N__26847\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19\
        );

    \I__4409\ : InMux
    port map (
            O => \N__26844\,
            I => \N__26841\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__26841\,
            I => \current_shift_inst.control_input_1_axb_14\
        );

    \I__4407\ : InMux
    port map (
            O => \N__26838\,
            I => \current_shift_inst.un38_control_input_0_cry_19\
        );

    \I__4406\ : InMux
    port map (
            O => \N__26835\,
            I => \N__26832\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__26832\,
            I => \N__26829\
        );

    \I__4404\ : Odrv4
    port map (
            O => \N__26829\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIDR081_20\
        );

    \I__4403\ : CascadeMux
    port map (
            O => \N__26826\,
            I => \N__26823\
        );

    \I__4402\ : InMux
    port map (
            O => \N__26823\,
            I => \N__26820\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__26820\,
            I => \N__26817\
        );

    \I__4400\ : Odrv12
    port map (
            O => \N__26817\,
            I => \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20\
        );

    \I__4399\ : InMux
    port map (
            O => \N__26814\,
            I => \N__26811\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__26811\,
            I => \current_shift_inst.control_input_1_axb_15\
        );

    \I__4397\ : InMux
    port map (
            O => \N__26808\,
            I => \current_shift_inst.un38_control_input_0_cry_20\
        );

    \I__4396\ : InMux
    port map (
            O => \N__26805\,
            I => \N__26802\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__26802\,
            I => \N__26799\
        );

    \I__4394\ : Odrv4
    port map (
            O => \N__26799\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21\
        );

    \I__4393\ : CascadeMux
    port map (
            O => \N__26796\,
            I => \N__26793\
        );

    \I__4392\ : InMux
    port map (
            O => \N__26793\,
            I => \N__26790\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__26790\,
            I => \N__26787\
        );

    \I__4390\ : Odrv4
    port map (
            O => \N__26787\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21\
        );

    \I__4389\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26781\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__26781\,
            I => \current_shift_inst.control_input_1_axb_16\
        );

    \I__4387\ : InMux
    port map (
            O => \N__26778\,
            I => \current_shift_inst.un38_control_input_0_cry_21\
        );

    \I__4386\ : InMux
    port map (
            O => \N__26775\,
            I => \bfn_9_14_0_\
        );

    \I__4385\ : InMux
    port map (
            O => \N__26772\,
            I => \N__26769\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__26769\,
            I => \current_shift_inst.control_input_1_axb_2\
        );

    \I__4383\ : InMux
    port map (
            O => \N__26766\,
            I => \current_shift_inst.un38_control_input_0_cry_7\
        );

    \I__4382\ : InMux
    port map (
            O => \N__26763\,
            I => \N__26760\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__26760\,
            I => \N__26757\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__26757\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8\
        );

    \I__4379\ : InMux
    port map (
            O => \N__26754\,
            I => \N__26751\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__26751\,
            I => \current_shift_inst.control_input_1_axb_3\
        );

    \I__4377\ : InMux
    port map (
            O => \N__26748\,
            I => \current_shift_inst.un38_control_input_0_cry_8\
        );

    \I__4376\ : InMux
    port map (
            O => \N__26745\,
            I => \N__26742\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__26742\,
            I => \N__26739\
        );

    \I__4374\ : Odrv4
    port map (
            O => \N__26739\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10\
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__26736\,
            I => \N__26733\
        );

    \I__4372\ : InMux
    port map (
            O => \N__26733\,
            I => \N__26730\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__26730\,
            I => \N__26727\
        );

    \I__4370\ : Span4Mux_h
    port map (
            O => \N__26727\,
            I => \N__26724\
        );

    \I__4369\ : Odrv4
    port map (
            O => \N__26724\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9\
        );

    \I__4368\ : InMux
    port map (
            O => \N__26721\,
            I => \N__26718\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__26718\,
            I => \current_shift_inst.control_input_1_axb_4\
        );

    \I__4366\ : InMux
    port map (
            O => \N__26715\,
            I => \current_shift_inst.un38_control_input_0_cry_9\
        );

    \I__4365\ : InMux
    port map (
            O => \N__26712\,
            I => \N__26709\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__26709\,
            I => \N__26706\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__26706\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10\
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__26703\,
            I => \N__26700\
        );

    \I__4361\ : InMux
    port map (
            O => \N__26700\,
            I => \N__26697\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__26697\,
            I => \N__26694\
        );

    \I__4359\ : Span4Mux_h
    port map (
            O => \N__26694\,
            I => \N__26691\
        );

    \I__4358\ : Odrv4
    port map (
            O => \N__26691\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10\
        );

    \I__4357\ : InMux
    port map (
            O => \N__26688\,
            I => \N__26685\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__26685\,
            I => \current_shift_inst.control_input_1_axb_5\
        );

    \I__4355\ : InMux
    port map (
            O => \N__26682\,
            I => \current_shift_inst.un38_control_input_0_cry_10\
        );

    \I__4354\ : CascadeMux
    port map (
            O => \N__26679\,
            I => \N__26676\
        );

    \I__4353\ : InMux
    port map (
            O => \N__26676\,
            I => \N__26673\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__26673\,
            I => \N__26670\
        );

    \I__4351\ : Odrv4
    port map (
            O => \N__26670\,
            I => \current_shift_inst.elapsed_time_ns_1_RNILORI_11\
        );

    \I__4350\ : InMux
    port map (
            O => \N__26667\,
            I => \N__26664\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__26664\,
            I => \current_shift_inst.control_input_1_axb_6\
        );

    \I__4348\ : InMux
    port map (
            O => \N__26661\,
            I => \current_shift_inst.un38_control_input_0_cry_11\
        );

    \I__4347\ : InMux
    port map (
            O => \N__26658\,
            I => \N__26655\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__26655\,
            I => \current_shift_inst.control_input_1_axb_7\
        );

    \I__4345\ : InMux
    port map (
            O => \N__26652\,
            I => \current_shift_inst.un38_control_input_0_cry_12\
        );

    \I__4344\ : CascadeMux
    port map (
            O => \N__26649\,
            I => \N__26646\
        );

    \I__4343\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26643\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__26643\,
            I => \N__26640\
        );

    \I__4341\ : Odrv4
    port map (
            O => \N__26640\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13\
        );

    \I__4340\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26634\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__26634\,
            I => \current_shift_inst.control_input_1_axb_8\
        );

    \I__4338\ : InMux
    port map (
            O => \N__26631\,
            I => \current_shift_inst.un38_control_input_0_cry_13\
        );

    \I__4337\ : InMux
    port map (
            O => \N__26628\,
            I => \N__26625\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__26625\,
            I => \current_shift_inst.z_i_0_31\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__26622\,
            I => \N__26619\
        );

    \I__4334\ : InMux
    port map (
            O => \N__26619\,
            I => \N__26616\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__26616\,
            I => \current_shift_inst.un38_control_input_0_cry_3_c_invZ0\
        );

    \I__4332\ : InMux
    port map (
            O => \N__26613\,
            I => \N__26610\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__26610\,
            I => \current_shift_inst.control_input_1_axb_0\
        );

    \I__4330\ : InMux
    port map (
            O => \N__26607\,
            I => \current_shift_inst.un38_control_input_0_cry_5\
        );

    \I__4329\ : InMux
    port map (
            O => \N__26604\,
            I => \N__26601\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__26601\,
            I => \current_shift_inst.control_input_1_axb_1\
        );

    \I__4327\ : InMux
    port map (
            O => \N__26598\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29\
        );

    \I__4326\ : InMux
    port map (
            O => \N__26595\,
            I => \N__26571\
        );

    \I__4325\ : InMux
    port map (
            O => \N__26594\,
            I => \N__26571\
        );

    \I__4324\ : InMux
    port map (
            O => \N__26593\,
            I => \N__26571\
        );

    \I__4323\ : InMux
    port map (
            O => \N__26592\,
            I => \N__26571\
        );

    \I__4322\ : InMux
    port map (
            O => \N__26591\,
            I => \N__26562\
        );

    \I__4321\ : InMux
    port map (
            O => \N__26590\,
            I => \N__26562\
        );

    \I__4320\ : InMux
    port map (
            O => \N__26589\,
            I => \N__26562\
        );

    \I__4319\ : InMux
    port map (
            O => \N__26588\,
            I => \N__26562\
        );

    \I__4318\ : InMux
    port map (
            O => \N__26587\,
            I => \N__26553\
        );

    \I__4317\ : InMux
    port map (
            O => \N__26586\,
            I => \N__26553\
        );

    \I__4316\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26553\
        );

    \I__4315\ : InMux
    port map (
            O => \N__26584\,
            I => \N__26553\
        );

    \I__4314\ : InMux
    port map (
            O => \N__26583\,
            I => \N__26544\
        );

    \I__4313\ : InMux
    port map (
            O => \N__26582\,
            I => \N__26544\
        );

    \I__4312\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26544\
        );

    \I__4311\ : InMux
    port map (
            O => \N__26580\,
            I => \N__26544\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__26571\,
            I => \N__26525\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__26562\,
            I => \N__26525\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__26553\,
            I => \N__26520\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__26544\,
            I => \N__26520\
        );

    \I__4306\ : InMux
    port map (
            O => \N__26543\,
            I => \N__26511\
        );

    \I__4305\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26511\
        );

    \I__4304\ : InMux
    port map (
            O => \N__26541\,
            I => \N__26511\
        );

    \I__4303\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26511\
        );

    \I__4302\ : InMux
    port map (
            O => \N__26539\,
            I => \N__26502\
        );

    \I__4301\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26502\
        );

    \I__4300\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26502\
        );

    \I__4299\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26502\
        );

    \I__4298\ : InMux
    port map (
            O => \N__26535\,
            I => \N__26497\
        );

    \I__4297\ : InMux
    port map (
            O => \N__26534\,
            I => \N__26497\
        );

    \I__4296\ : InMux
    port map (
            O => \N__26533\,
            I => \N__26488\
        );

    \I__4295\ : InMux
    port map (
            O => \N__26532\,
            I => \N__26488\
        );

    \I__4294\ : InMux
    port map (
            O => \N__26531\,
            I => \N__26488\
        );

    \I__4293\ : InMux
    port map (
            O => \N__26530\,
            I => \N__26488\
        );

    \I__4292\ : Span4Mux_h
    port map (
            O => \N__26525\,
            I => \N__26485\
        );

    \I__4291\ : Span4Mux_v
    port map (
            O => \N__26520\,
            I => \N__26482\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__26511\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__26502\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__26497\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__26488\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__4286\ : Odrv4
    port map (
            O => \N__26485\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__4285\ : Odrv4
    port map (
            O => \N__26482\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__4284\ : InMux
    port map (
            O => \N__26469\,
            I => \N__26466\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__26466\,
            I => \N__26463\
        );

    \I__4282\ : Odrv12
    port map (
            O => \N__26463\,
            I => il_min_comp1_c
        );

    \I__4281\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26457\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__26457\,
            I => \current_shift_inst.S1_syncZ0Z0\
        );

    \I__4279\ : InMux
    port map (
            O => \N__26454\,
            I => \N__26448\
        );

    \I__4278\ : InMux
    port map (
            O => \N__26453\,
            I => \N__26448\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__26448\,
            I => \current_shift_inst.S1_syncZ0Z1\
        );

    \I__4276\ : InMux
    port map (
            O => \N__26445\,
            I => \N__26442\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__26442\,
            I => \current_shift_inst.S1_sync_prevZ0\
        );

    \I__4274\ : CascadeMux
    port map (
            O => \N__26439\,
            I => \N__26436\
        );

    \I__4273\ : InMux
    port map (
            O => \N__26436\,
            I => \N__26432\
        );

    \I__4272\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26429\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__26432\,
            I => \N__26423\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__26429\,
            I => \N__26423\
        );

    \I__4269\ : InMux
    port map (
            O => \N__26428\,
            I => \N__26420\
        );

    \I__4268\ : Span4Mux_h
    port map (
            O => \N__26423\,
            I => \N__26417\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__26420\,
            I => \current_shift_inst.timer_phase.counterZ0Z_20\
        );

    \I__4266\ : Odrv4
    port map (
            O => \N__26417\,
            I => \current_shift_inst.timer_phase.counterZ0Z_20\
        );

    \I__4265\ : InMux
    port map (
            O => \N__26412\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\
        );

    \I__4264\ : CascadeMux
    port map (
            O => \N__26409\,
            I => \N__26406\
        );

    \I__4263\ : InMux
    port map (
            O => \N__26406\,
            I => \N__26402\
        );

    \I__4262\ : InMux
    port map (
            O => \N__26405\,
            I => \N__26399\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__26402\,
            I => \N__26393\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__26399\,
            I => \N__26393\
        );

    \I__4259\ : InMux
    port map (
            O => \N__26398\,
            I => \N__26390\
        );

    \I__4258\ : Span4Mux_h
    port map (
            O => \N__26393\,
            I => \N__26387\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__26390\,
            I => \current_shift_inst.timer_phase.counterZ0Z_21\
        );

    \I__4256\ : Odrv4
    port map (
            O => \N__26387\,
            I => \current_shift_inst.timer_phase.counterZ0Z_21\
        );

    \I__4255\ : InMux
    port map (
            O => \N__26382\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\
        );

    \I__4254\ : InMux
    port map (
            O => \N__26379\,
            I => \N__26372\
        );

    \I__4253\ : InMux
    port map (
            O => \N__26378\,
            I => \N__26372\
        );

    \I__4252\ : InMux
    port map (
            O => \N__26377\,
            I => \N__26369\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__26372\,
            I => \N__26366\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__26369\,
            I => \current_shift_inst.timer_phase.counterZ0Z_22\
        );

    \I__4249\ : Odrv4
    port map (
            O => \N__26366\,
            I => \current_shift_inst.timer_phase.counterZ0Z_22\
        );

    \I__4248\ : InMux
    port map (
            O => \N__26361\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\
        );

    \I__4247\ : InMux
    port map (
            O => \N__26358\,
            I => \N__26351\
        );

    \I__4246\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26351\
        );

    \I__4245\ : InMux
    port map (
            O => \N__26356\,
            I => \N__26348\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__26351\,
            I => \N__26345\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__26348\,
            I => \current_shift_inst.timer_phase.counterZ0Z_23\
        );

    \I__4242\ : Odrv4
    port map (
            O => \N__26345\,
            I => \current_shift_inst.timer_phase.counterZ0Z_23\
        );

    \I__4241\ : InMux
    port map (
            O => \N__26340\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\
        );

    \I__4240\ : CascadeMux
    port map (
            O => \N__26337\,
            I => \N__26333\
        );

    \I__4239\ : InMux
    port map (
            O => \N__26336\,
            I => \N__26329\
        );

    \I__4238\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26326\
        );

    \I__4237\ : InMux
    port map (
            O => \N__26332\,
            I => \N__26323\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__26329\,
            I => \N__26318\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__26326\,
            I => \N__26318\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__26323\,
            I => \current_shift_inst.timer_phase.counterZ0Z_24\
        );

    \I__4233\ : Odrv4
    port map (
            O => \N__26318\,
            I => \current_shift_inst.timer_phase.counterZ0Z_24\
        );

    \I__4232\ : InMux
    port map (
            O => \N__26313\,
            I => \bfn_8_20_0_\
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__26310\,
            I => \N__26306\
        );

    \I__4230\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26302\
        );

    \I__4229\ : InMux
    port map (
            O => \N__26306\,
            I => \N__26299\
        );

    \I__4228\ : InMux
    port map (
            O => \N__26305\,
            I => \N__26296\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__26302\,
            I => \N__26291\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__26299\,
            I => \N__26291\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__26296\,
            I => \current_shift_inst.timer_phase.counterZ0Z_25\
        );

    \I__4224\ : Odrv4
    port map (
            O => \N__26291\,
            I => \current_shift_inst.timer_phase.counterZ0Z_25\
        );

    \I__4223\ : InMux
    port map (
            O => \N__26286\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\
        );

    \I__4222\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26280\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__26280\,
            I => \N__26276\
        );

    \I__4220\ : InMux
    port map (
            O => \N__26279\,
            I => \N__26273\
        );

    \I__4219\ : Span4Mux_h
    port map (
            O => \N__26276\,
            I => \N__26270\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__26273\,
            I => \current_shift_inst.timer_phase.counterZ0Z_28\
        );

    \I__4217\ : Odrv4
    port map (
            O => \N__26270\,
            I => \current_shift_inst.timer_phase.counterZ0Z_28\
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__26265\,
            I => \N__26261\
        );

    \I__4215\ : CascadeMux
    port map (
            O => \N__26264\,
            I => \N__26258\
        );

    \I__4214\ : InMux
    port map (
            O => \N__26261\,
            I => \N__26252\
        );

    \I__4213\ : InMux
    port map (
            O => \N__26258\,
            I => \N__26252\
        );

    \I__4212\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26249\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__26252\,
            I => \N__26246\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__26249\,
            I => \current_shift_inst.timer_phase.counterZ0Z_26\
        );

    \I__4209\ : Odrv4
    port map (
            O => \N__26246\,
            I => \current_shift_inst.timer_phase.counterZ0Z_26\
        );

    \I__4208\ : InMux
    port map (
            O => \N__26241\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\
        );

    \I__4207\ : InMux
    port map (
            O => \N__26238\,
            I => \N__26235\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__26235\,
            I => \N__26231\
        );

    \I__4205\ : InMux
    port map (
            O => \N__26234\,
            I => \N__26228\
        );

    \I__4204\ : Span4Mux_h
    port map (
            O => \N__26231\,
            I => \N__26225\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__26228\,
            I => \current_shift_inst.timer_phase.counterZ0Z_29\
        );

    \I__4202\ : Odrv4
    port map (
            O => \N__26225\,
            I => \current_shift_inst.timer_phase.counterZ0Z_29\
        );

    \I__4201\ : CascadeMux
    port map (
            O => \N__26220\,
            I => \N__26216\
        );

    \I__4200\ : CascadeMux
    port map (
            O => \N__26219\,
            I => \N__26213\
        );

    \I__4199\ : InMux
    port map (
            O => \N__26216\,
            I => \N__26207\
        );

    \I__4198\ : InMux
    port map (
            O => \N__26213\,
            I => \N__26207\
        );

    \I__4197\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26204\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__26207\,
            I => \N__26201\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__26204\,
            I => \current_shift_inst.timer_phase.counterZ0Z_27\
        );

    \I__4194\ : Odrv4
    port map (
            O => \N__26201\,
            I => \current_shift_inst.timer_phase.counterZ0Z_27\
        );

    \I__4193\ : InMux
    port map (
            O => \N__26196\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\
        );

    \I__4192\ : CascadeMux
    port map (
            O => \N__26193\,
            I => \N__26190\
        );

    \I__4191\ : InMux
    port map (
            O => \N__26190\,
            I => \N__26186\
        );

    \I__4190\ : InMux
    port map (
            O => \N__26189\,
            I => \N__26183\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__26186\,
            I => \N__26177\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__26183\,
            I => \N__26177\
        );

    \I__4187\ : InMux
    port map (
            O => \N__26182\,
            I => \N__26174\
        );

    \I__4186\ : Span4Mux_h
    port map (
            O => \N__26177\,
            I => \N__26171\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__26174\,
            I => \current_shift_inst.timer_phase.counterZ0Z_12\
        );

    \I__4184\ : Odrv4
    port map (
            O => \N__26171\,
            I => \current_shift_inst.timer_phase.counterZ0Z_12\
        );

    \I__4183\ : InMux
    port map (
            O => \N__26166\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__26163\,
            I => \N__26160\
        );

    \I__4181\ : InMux
    port map (
            O => \N__26160\,
            I => \N__26156\
        );

    \I__4180\ : InMux
    port map (
            O => \N__26159\,
            I => \N__26153\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__26156\,
            I => \N__26147\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__26153\,
            I => \N__26147\
        );

    \I__4177\ : InMux
    port map (
            O => \N__26152\,
            I => \N__26144\
        );

    \I__4176\ : Span4Mux_h
    port map (
            O => \N__26147\,
            I => \N__26141\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__26144\,
            I => \current_shift_inst.timer_phase.counterZ0Z_13\
        );

    \I__4174\ : Odrv4
    port map (
            O => \N__26141\,
            I => \current_shift_inst.timer_phase.counterZ0Z_13\
        );

    \I__4173\ : InMux
    port map (
            O => \N__26136\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\
        );

    \I__4172\ : InMux
    port map (
            O => \N__26133\,
            I => \N__26126\
        );

    \I__4171\ : InMux
    port map (
            O => \N__26132\,
            I => \N__26126\
        );

    \I__4170\ : InMux
    port map (
            O => \N__26131\,
            I => \N__26123\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__26126\,
            I => \N__26120\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__26123\,
            I => \current_shift_inst.timer_phase.counterZ0Z_14\
        );

    \I__4167\ : Odrv4
    port map (
            O => \N__26120\,
            I => \current_shift_inst.timer_phase.counterZ0Z_14\
        );

    \I__4166\ : InMux
    port map (
            O => \N__26115\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\
        );

    \I__4165\ : InMux
    port map (
            O => \N__26112\,
            I => \N__26105\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26111\,
            I => \N__26105\
        );

    \I__4163\ : InMux
    port map (
            O => \N__26110\,
            I => \N__26102\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__26105\,
            I => \N__26099\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__26102\,
            I => \current_shift_inst.timer_phase.counterZ0Z_15\
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__26099\,
            I => \current_shift_inst.timer_phase.counterZ0Z_15\
        );

    \I__4159\ : InMux
    port map (
            O => \N__26094\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__26091\,
            I => \N__26087\
        );

    \I__4157\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26083\
        );

    \I__4156\ : InMux
    port map (
            O => \N__26087\,
            I => \N__26080\
        );

    \I__4155\ : InMux
    port map (
            O => \N__26086\,
            I => \N__26077\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__26083\,
            I => \N__26072\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__26080\,
            I => \N__26072\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__26077\,
            I => \current_shift_inst.timer_phase.counterZ0Z_16\
        );

    \I__4151\ : Odrv4
    port map (
            O => \N__26072\,
            I => \current_shift_inst.timer_phase.counterZ0Z_16\
        );

    \I__4150\ : InMux
    port map (
            O => \N__26067\,
            I => \bfn_8_19_0_\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__26064\,
            I => \N__26060\
        );

    \I__4148\ : InMux
    port map (
            O => \N__26063\,
            I => \N__26056\
        );

    \I__4147\ : InMux
    port map (
            O => \N__26060\,
            I => \N__26053\
        );

    \I__4146\ : InMux
    port map (
            O => \N__26059\,
            I => \N__26050\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__26056\,
            I => \N__26045\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__26053\,
            I => \N__26045\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__26050\,
            I => \current_shift_inst.timer_phase.counterZ0Z_17\
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__26045\,
            I => \current_shift_inst.timer_phase.counterZ0Z_17\
        );

    \I__4141\ : InMux
    port map (
            O => \N__26040\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\
        );

    \I__4140\ : CascadeMux
    port map (
            O => \N__26037\,
            I => \N__26033\
        );

    \I__4139\ : CascadeMux
    port map (
            O => \N__26036\,
            I => \N__26030\
        );

    \I__4138\ : InMux
    port map (
            O => \N__26033\,
            I => \N__26024\
        );

    \I__4137\ : InMux
    port map (
            O => \N__26030\,
            I => \N__26024\
        );

    \I__4136\ : InMux
    port map (
            O => \N__26029\,
            I => \N__26021\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__26024\,
            I => \N__26018\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__26021\,
            I => \current_shift_inst.timer_phase.counterZ0Z_18\
        );

    \I__4133\ : Odrv4
    port map (
            O => \N__26018\,
            I => \current_shift_inst.timer_phase.counterZ0Z_18\
        );

    \I__4132\ : InMux
    port map (
            O => \N__26013\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\
        );

    \I__4131\ : CascadeMux
    port map (
            O => \N__26010\,
            I => \N__26006\
        );

    \I__4130\ : CascadeMux
    port map (
            O => \N__26009\,
            I => \N__26003\
        );

    \I__4129\ : InMux
    port map (
            O => \N__26006\,
            I => \N__25997\
        );

    \I__4128\ : InMux
    port map (
            O => \N__26003\,
            I => \N__25997\
        );

    \I__4127\ : InMux
    port map (
            O => \N__26002\,
            I => \N__25994\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__25997\,
            I => \N__25991\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__25994\,
            I => \current_shift_inst.timer_phase.counterZ0Z_19\
        );

    \I__4124\ : Odrv4
    port map (
            O => \N__25991\,
            I => \current_shift_inst.timer_phase.counterZ0Z_19\
        );

    \I__4123\ : InMux
    port map (
            O => \N__25986\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\
        );

    \I__4122\ : CascadeMux
    port map (
            O => \N__25983\,
            I => \N__25979\
        );

    \I__4121\ : CascadeMux
    port map (
            O => \N__25982\,
            I => \N__25976\
        );

    \I__4120\ : InMux
    port map (
            O => \N__25979\,
            I => \N__25970\
        );

    \I__4119\ : InMux
    port map (
            O => \N__25976\,
            I => \N__25970\
        );

    \I__4118\ : InMux
    port map (
            O => \N__25975\,
            I => \N__25967\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__25970\,
            I => \N__25964\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__25967\,
            I => \current_shift_inst.timer_phase.counterZ0Z_3\
        );

    \I__4115\ : Odrv4
    port map (
            O => \N__25964\,
            I => \current_shift_inst.timer_phase.counterZ0Z_3\
        );

    \I__4114\ : InMux
    port map (
            O => \N__25959\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\
        );

    \I__4113\ : InMux
    port map (
            O => \N__25956\,
            I => \N__25950\
        );

    \I__4112\ : InMux
    port map (
            O => \N__25955\,
            I => \N__25950\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__25950\,
            I => \N__25946\
        );

    \I__4110\ : InMux
    port map (
            O => \N__25949\,
            I => \N__25943\
        );

    \I__4109\ : Span4Mux_h
    port map (
            O => \N__25946\,
            I => \N__25940\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__25943\,
            I => \current_shift_inst.timer_phase.counterZ0Z_4\
        );

    \I__4107\ : Odrv4
    port map (
            O => \N__25940\,
            I => \current_shift_inst.timer_phase.counterZ0Z_4\
        );

    \I__4106\ : InMux
    port map (
            O => \N__25935\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\
        );

    \I__4105\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25925\
        );

    \I__4104\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25925\
        );

    \I__4103\ : InMux
    port map (
            O => \N__25930\,
            I => \N__25922\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__25925\,
            I => \N__25919\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__25922\,
            I => \current_shift_inst.timer_phase.counterZ0Z_5\
        );

    \I__4100\ : Odrv4
    port map (
            O => \N__25919\,
            I => \current_shift_inst.timer_phase.counterZ0Z_5\
        );

    \I__4099\ : InMux
    port map (
            O => \N__25914\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\
        );

    \I__4098\ : CascadeMux
    port map (
            O => \N__25911\,
            I => \N__25907\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__25910\,
            I => \N__25904\
        );

    \I__4096\ : InMux
    port map (
            O => \N__25907\,
            I => \N__25899\
        );

    \I__4095\ : InMux
    port map (
            O => \N__25904\,
            I => \N__25899\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__25899\,
            I => \N__25895\
        );

    \I__4093\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25892\
        );

    \I__4092\ : Span4Mux_h
    port map (
            O => \N__25895\,
            I => \N__25889\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__25892\,
            I => \current_shift_inst.timer_phase.counterZ0Z_6\
        );

    \I__4090\ : Odrv4
    port map (
            O => \N__25889\,
            I => \current_shift_inst.timer_phase.counterZ0Z_6\
        );

    \I__4089\ : InMux
    port map (
            O => \N__25884\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__25881\,
            I => \N__25877\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__25880\,
            I => \N__25874\
        );

    \I__4086\ : InMux
    port map (
            O => \N__25877\,
            I => \N__25869\
        );

    \I__4085\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25869\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__25869\,
            I => \N__25865\
        );

    \I__4083\ : InMux
    port map (
            O => \N__25868\,
            I => \N__25862\
        );

    \I__4082\ : Span4Mux_h
    port map (
            O => \N__25865\,
            I => \N__25859\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__25862\,
            I => \current_shift_inst.timer_phase.counterZ0Z_7\
        );

    \I__4080\ : Odrv4
    port map (
            O => \N__25859\,
            I => \current_shift_inst.timer_phase.counterZ0Z_7\
        );

    \I__4079\ : InMux
    port map (
            O => \N__25854\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\
        );

    \I__4078\ : InMux
    port map (
            O => \N__25851\,
            I => \N__25847\
        );

    \I__4077\ : InMux
    port map (
            O => \N__25850\,
            I => \N__25844\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__25847\,
            I => \N__25840\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__25844\,
            I => \N__25837\
        );

    \I__4074\ : InMux
    port map (
            O => \N__25843\,
            I => \N__25834\
        );

    \I__4073\ : Span4Mux_h
    port map (
            O => \N__25840\,
            I => \N__25831\
        );

    \I__4072\ : Odrv4
    port map (
            O => \N__25837\,
            I => \current_shift_inst.timer_phase.counterZ0Z_8\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__25834\,
            I => \current_shift_inst.timer_phase.counterZ0Z_8\
        );

    \I__4070\ : Odrv4
    port map (
            O => \N__25831\,
            I => \current_shift_inst.timer_phase.counterZ0Z_8\
        );

    \I__4069\ : InMux
    port map (
            O => \N__25824\,
            I => \bfn_8_18_0_\
        );

    \I__4068\ : InMux
    port map (
            O => \N__25821\,
            I => \N__25817\
        );

    \I__4067\ : InMux
    port map (
            O => \N__25820\,
            I => \N__25814\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__25817\,
            I => \N__25810\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__25814\,
            I => \N__25807\
        );

    \I__4064\ : InMux
    port map (
            O => \N__25813\,
            I => \N__25804\
        );

    \I__4063\ : Span4Mux_h
    port map (
            O => \N__25810\,
            I => \N__25801\
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__25807\,
            I => \current_shift_inst.timer_phase.counterZ0Z_9\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__25804\,
            I => \current_shift_inst.timer_phase.counterZ0Z_9\
        );

    \I__4060\ : Odrv4
    port map (
            O => \N__25801\,
            I => \current_shift_inst.timer_phase.counterZ0Z_9\
        );

    \I__4059\ : InMux
    port map (
            O => \N__25794\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\
        );

    \I__4058\ : CascadeMux
    port map (
            O => \N__25791\,
            I => \N__25787\
        );

    \I__4057\ : CascadeMux
    port map (
            O => \N__25790\,
            I => \N__25784\
        );

    \I__4056\ : InMux
    port map (
            O => \N__25787\,
            I => \N__25778\
        );

    \I__4055\ : InMux
    port map (
            O => \N__25784\,
            I => \N__25778\
        );

    \I__4054\ : InMux
    port map (
            O => \N__25783\,
            I => \N__25775\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__25778\,
            I => \N__25772\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__25775\,
            I => \current_shift_inst.timer_phase.counterZ0Z_10\
        );

    \I__4051\ : Odrv4
    port map (
            O => \N__25772\,
            I => \current_shift_inst.timer_phase.counterZ0Z_10\
        );

    \I__4050\ : InMux
    port map (
            O => \N__25767\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__25764\,
            I => \N__25760\
        );

    \I__4048\ : CascadeMux
    port map (
            O => \N__25763\,
            I => \N__25757\
        );

    \I__4047\ : InMux
    port map (
            O => \N__25760\,
            I => \N__25751\
        );

    \I__4046\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25751\
        );

    \I__4045\ : InMux
    port map (
            O => \N__25756\,
            I => \N__25748\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__25751\,
            I => \N__25745\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__25748\,
            I => \current_shift_inst.timer_phase.counterZ0Z_11\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__25745\,
            I => \current_shift_inst.timer_phase.counterZ0Z_11\
        );

    \I__4041\ : InMux
    port map (
            O => \N__25740\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\
        );

    \I__4040\ : CascadeMux
    port map (
            O => \N__25737\,
            I => \N__25734\
        );

    \I__4039\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25730\
        );

    \I__4038\ : InMux
    port map (
            O => \N__25733\,
            I => \N__25727\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__25730\,
            I => \N__25724\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__25727\,
            I => \N__25721\
        );

    \I__4035\ : Span4Mux_v
    port map (
            O => \N__25724\,
            I => \N__25718\
        );

    \I__4034\ : Odrv4
    port map (
            O => \N__25721\,
            I => \current_shift_inst.control_inputZ0Z_21\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__25718\,
            I => \current_shift_inst.control_inputZ0Z_21\
        );

    \I__4032\ : InMux
    port map (
            O => \N__25713\,
            I => \current_shift_inst.control_input_1_cry_20\
        );

    \I__4031\ : CascadeMux
    port map (
            O => \N__25710\,
            I => \N__25706\
        );

    \I__4030\ : InMux
    port map (
            O => \N__25709\,
            I => \N__25703\
        );

    \I__4029\ : InMux
    port map (
            O => \N__25706\,
            I => \N__25700\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__25703\,
            I => \N__25697\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__25700\,
            I => \N__25694\
        );

    \I__4026\ : Span4Mux_h
    port map (
            O => \N__25697\,
            I => \N__25689\
        );

    \I__4025\ : Span4Mux_h
    port map (
            O => \N__25694\,
            I => \N__25689\
        );

    \I__4024\ : Odrv4
    port map (
            O => \N__25689\,
            I => \current_shift_inst.control_inputZ0Z_22\
        );

    \I__4023\ : InMux
    port map (
            O => \N__25686\,
            I => \current_shift_inst.control_input_1_cry_21\
        );

    \I__4022\ : CascadeMux
    port map (
            O => \N__25683\,
            I => \N__25679\
        );

    \I__4021\ : InMux
    port map (
            O => \N__25682\,
            I => \N__25676\
        );

    \I__4020\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25673\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__25676\,
            I => \N__25670\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__25673\,
            I => \N__25667\
        );

    \I__4017\ : Span4Mux_h
    port map (
            O => \N__25670\,
            I => \N__25662\
        );

    \I__4016\ : Span4Mux_h
    port map (
            O => \N__25667\,
            I => \N__25662\
        );

    \I__4015\ : Odrv4
    port map (
            O => \N__25662\,
            I => \current_shift_inst.control_inputZ0Z_23\
        );

    \I__4014\ : InMux
    port map (
            O => \N__25659\,
            I => \current_shift_inst.control_input_1_cry_22\
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__25656\,
            I => \N__25653\
        );

    \I__4012\ : InMux
    port map (
            O => \N__25653\,
            I => \N__25649\
        );

    \I__4011\ : InMux
    port map (
            O => \N__25652\,
            I => \N__25646\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__25649\,
            I => \N__25643\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__25646\,
            I => \N__25640\
        );

    \I__4008\ : Span4Mux_h
    port map (
            O => \N__25643\,
            I => \N__25637\
        );

    \I__4007\ : Odrv12
    port map (
            O => \N__25640\,
            I => \current_shift_inst.control_inputZ0Z_24\
        );

    \I__4006\ : Odrv4
    port map (
            O => \N__25637\,
            I => \current_shift_inst.control_inputZ0Z_24\
        );

    \I__4005\ : InMux
    port map (
            O => \N__25632\,
            I => \bfn_8_16_0_\
        );

    \I__4004\ : InMux
    port map (
            O => \N__25629\,
            I => \current_shift_inst.control_input_1_cry_24\
        );

    \I__4003\ : InMux
    port map (
            O => \N__25626\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__25623\,
            I => \N__25619\
        );

    \I__4001\ : CascadeMux
    port map (
            O => \N__25622\,
            I => \N__25616\
        );

    \I__4000\ : InMux
    port map (
            O => \N__25619\,
            I => \N__25610\
        );

    \I__3999\ : InMux
    port map (
            O => \N__25616\,
            I => \N__25610\
        );

    \I__3998\ : InMux
    port map (
            O => \N__25615\,
            I => \N__25607\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__25610\,
            I => \N__25604\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__25607\,
            I => \current_shift_inst.timer_phase.counterZ0Z_2\
        );

    \I__3995\ : Odrv4
    port map (
            O => \N__25604\,
            I => \current_shift_inst.timer_phase.counterZ0Z_2\
        );

    \I__3994\ : InMux
    port map (
            O => \N__25599\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\
        );

    \I__3993\ : InMux
    port map (
            O => \N__25596\,
            I => \N__25592\
        );

    \I__3992\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25589\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__25592\,
            I => \N__25584\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__25589\,
            I => \N__25584\
        );

    \I__3989\ : Span4Mux_v
    port map (
            O => \N__25584\,
            I => \N__25581\
        );

    \I__3988\ : Odrv4
    port map (
            O => \N__25581\,
            I => \current_shift_inst.control_inputZ0Z_12\
        );

    \I__3987\ : InMux
    port map (
            O => \N__25578\,
            I => \current_shift_inst.control_input_1_cry_11\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__25575\,
            I => \N__25571\
        );

    \I__3985\ : InMux
    port map (
            O => \N__25574\,
            I => \N__25568\
        );

    \I__3984\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25565\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__25568\,
            I => \N__25560\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__25565\,
            I => \N__25560\
        );

    \I__3981\ : Span4Mux_v
    port map (
            O => \N__25560\,
            I => \N__25557\
        );

    \I__3980\ : Odrv4
    port map (
            O => \N__25557\,
            I => \current_shift_inst.control_inputZ0Z_13\
        );

    \I__3979\ : InMux
    port map (
            O => \N__25554\,
            I => \current_shift_inst.control_input_1_cry_12\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__25551\,
            I => \N__25547\
        );

    \I__3977\ : InMux
    port map (
            O => \N__25550\,
            I => \N__25544\
        );

    \I__3976\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25541\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__25544\,
            I => \N__25536\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__25541\,
            I => \N__25536\
        );

    \I__3973\ : Span4Mux_v
    port map (
            O => \N__25536\,
            I => \N__25533\
        );

    \I__3972\ : Odrv4
    port map (
            O => \N__25533\,
            I => \current_shift_inst.control_inputZ0Z_14\
        );

    \I__3971\ : InMux
    port map (
            O => \N__25530\,
            I => \current_shift_inst.control_input_1_cry_13\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__25527\,
            I => \N__25523\
        );

    \I__3969\ : InMux
    port map (
            O => \N__25526\,
            I => \N__25520\
        );

    \I__3968\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25517\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__25520\,
            I => \N__25512\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__25517\,
            I => \N__25512\
        );

    \I__3965\ : Span4Mux_v
    port map (
            O => \N__25512\,
            I => \N__25509\
        );

    \I__3964\ : Odrv4
    port map (
            O => \N__25509\,
            I => \current_shift_inst.control_inputZ0Z_15\
        );

    \I__3963\ : InMux
    port map (
            O => \N__25506\,
            I => \current_shift_inst.control_input_1_cry_14\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__25503\,
            I => \N__25500\
        );

    \I__3961\ : InMux
    port map (
            O => \N__25500\,
            I => \N__25496\
        );

    \I__3960\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25493\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__25496\,
            I => \N__25490\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__25493\,
            I => \N__25487\
        );

    \I__3957\ : Span4Mux_h
    port map (
            O => \N__25490\,
            I => \N__25484\
        );

    \I__3956\ : Odrv12
    port map (
            O => \N__25487\,
            I => \current_shift_inst.control_inputZ0Z_16\
        );

    \I__3955\ : Odrv4
    port map (
            O => \N__25484\,
            I => \current_shift_inst.control_inputZ0Z_16\
        );

    \I__3954\ : InMux
    port map (
            O => \N__25479\,
            I => \bfn_8_15_0_\
        );

    \I__3953\ : CascadeMux
    port map (
            O => \N__25476\,
            I => \N__25473\
        );

    \I__3952\ : InMux
    port map (
            O => \N__25473\,
            I => \N__25469\
        );

    \I__3951\ : InMux
    port map (
            O => \N__25472\,
            I => \N__25466\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__25469\,
            I => \N__25463\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__25466\,
            I => \N__25460\
        );

    \I__3948\ : Span12Mux_s8_h
    port map (
            O => \N__25463\,
            I => \N__25457\
        );

    \I__3947\ : Odrv12
    port map (
            O => \N__25460\,
            I => \current_shift_inst.control_inputZ0Z_17\
        );

    \I__3946\ : Odrv12
    port map (
            O => \N__25457\,
            I => \current_shift_inst.control_inputZ0Z_17\
        );

    \I__3945\ : InMux
    port map (
            O => \N__25452\,
            I => \current_shift_inst.control_input_1_cry_16\
        );

    \I__3944\ : CascadeMux
    port map (
            O => \N__25449\,
            I => \N__25446\
        );

    \I__3943\ : InMux
    port map (
            O => \N__25446\,
            I => \N__25443\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__25443\,
            I => \N__25439\
        );

    \I__3941\ : InMux
    port map (
            O => \N__25442\,
            I => \N__25436\
        );

    \I__3940\ : Span4Mux_v
    port map (
            O => \N__25439\,
            I => \N__25433\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__25436\,
            I => \N__25430\
        );

    \I__3938\ : Span4Mux_h
    port map (
            O => \N__25433\,
            I => \N__25427\
        );

    \I__3937\ : Odrv12
    port map (
            O => \N__25430\,
            I => \current_shift_inst.control_inputZ0Z_18\
        );

    \I__3936\ : Odrv4
    port map (
            O => \N__25427\,
            I => \current_shift_inst.control_inputZ0Z_18\
        );

    \I__3935\ : InMux
    port map (
            O => \N__25422\,
            I => \current_shift_inst.control_input_1_cry_17\
        );

    \I__3934\ : CascadeMux
    port map (
            O => \N__25419\,
            I => \N__25416\
        );

    \I__3933\ : InMux
    port map (
            O => \N__25416\,
            I => \N__25412\
        );

    \I__3932\ : InMux
    port map (
            O => \N__25415\,
            I => \N__25409\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__25412\,
            I => \N__25406\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__25409\,
            I => \N__25403\
        );

    \I__3929\ : Span4Mux_h
    port map (
            O => \N__25406\,
            I => \N__25400\
        );

    \I__3928\ : Odrv4
    port map (
            O => \N__25403\,
            I => \current_shift_inst.control_inputZ0Z_19\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__25400\,
            I => \current_shift_inst.control_inputZ0Z_19\
        );

    \I__3926\ : InMux
    port map (
            O => \N__25395\,
            I => \current_shift_inst.control_input_1_cry_18\
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__25392\,
            I => \N__25389\
        );

    \I__3924\ : InMux
    port map (
            O => \N__25389\,
            I => \N__25385\
        );

    \I__3923\ : InMux
    port map (
            O => \N__25388\,
            I => \N__25382\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__25385\,
            I => \N__25379\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__25382\,
            I => \N__25374\
        );

    \I__3920\ : Span4Mux_v
    port map (
            O => \N__25379\,
            I => \N__25374\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__25374\,
            I => \current_shift_inst.control_inputZ0Z_20\
        );

    \I__3918\ : InMux
    port map (
            O => \N__25371\,
            I => \current_shift_inst.control_input_1_cry_19\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__25368\,
            I => \N__25365\
        );

    \I__3916\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25362\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__25362\,
            I => \N__25358\
        );

    \I__3914\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25355\
        );

    \I__3913\ : Span4Mux_v
    port map (
            O => \N__25358\,
            I => \N__25352\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__25355\,
            I => \current_shift_inst.control_inputZ0Z_4\
        );

    \I__3911\ : Odrv4
    port map (
            O => \N__25352\,
            I => \current_shift_inst.control_inputZ0Z_4\
        );

    \I__3910\ : InMux
    port map (
            O => \N__25347\,
            I => \current_shift_inst.control_input_1_cry_3\
        );

    \I__3909\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25340\
        );

    \I__3908\ : CascadeMux
    port map (
            O => \N__25343\,
            I => \N__25337\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__25340\,
            I => \N__25334\
        );

    \I__3906\ : InMux
    port map (
            O => \N__25337\,
            I => \N__25331\
        );

    \I__3905\ : Span4Mux_h
    port map (
            O => \N__25334\,
            I => \N__25328\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__25331\,
            I => \N__25325\
        );

    \I__3903\ : Span4Mux_v
    port map (
            O => \N__25328\,
            I => \N__25322\
        );

    \I__3902\ : Span4Mux_v
    port map (
            O => \N__25325\,
            I => \N__25319\
        );

    \I__3901\ : Odrv4
    port map (
            O => \N__25322\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__25319\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__3899\ : InMux
    port map (
            O => \N__25314\,
            I => \current_shift_inst.control_input_1_cry_4\
        );

    \I__3898\ : CascadeMux
    port map (
            O => \N__25311\,
            I => \N__25307\
        );

    \I__3897\ : InMux
    port map (
            O => \N__25310\,
            I => \N__25304\
        );

    \I__3896\ : InMux
    port map (
            O => \N__25307\,
            I => \N__25301\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__25304\,
            I => \N__25298\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__25301\,
            I => \N__25295\
        );

    \I__3893\ : Span4Mux_h
    port map (
            O => \N__25298\,
            I => \N__25290\
        );

    \I__3892\ : Span4Mux_h
    port map (
            O => \N__25295\,
            I => \N__25290\
        );

    \I__3891\ : Odrv4
    port map (
            O => \N__25290\,
            I => \current_shift_inst.control_inputZ0Z_6\
        );

    \I__3890\ : InMux
    port map (
            O => \N__25287\,
            I => \current_shift_inst.control_input_1_cry_5\
        );

    \I__3889\ : InMux
    port map (
            O => \N__25284\,
            I => \N__25280\
        );

    \I__3888\ : CascadeMux
    port map (
            O => \N__25283\,
            I => \N__25277\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__25280\,
            I => \N__25274\
        );

    \I__3886\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25271\
        );

    \I__3885\ : Span4Mux_v
    port map (
            O => \N__25274\,
            I => \N__25266\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__25271\,
            I => \N__25266\
        );

    \I__3883\ : Span4Mux_h
    port map (
            O => \N__25266\,
            I => \N__25263\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__25263\,
            I => \N__25260\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__25260\,
            I => \current_shift_inst.control_inputZ0Z_7\
        );

    \I__3880\ : InMux
    port map (
            O => \N__25257\,
            I => \current_shift_inst.control_input_1_cry_6\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__25254\,
            I => \N__25250\
        );

    \I__3878\ : InMux
    port map (
            O => \N__25253\,
            I => \N__25247\
        );

    \I__3877\ : InMux
    port map (
            O => \N__25250\,
            I => \N__25244\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__25247\,
            I => \N__25241\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__25244\,
            I => \N__25238\
        );

    \I__3874\ : Span4Mux_h
    port map (
            O => \N__25241\,
            I => \N__25235\
        );

    \I__3873\ : Span4Mux_h
    port map (
            O => \N__25238\,
            I => \N__25232\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__25235\,
            I => \current_shift_inst.control_inputZ0Z_8\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__25232\,
            I => \current_shift_inst.control_inputZ0Z_8\
        );

    \I__3870\ : InMux
    port map (
            O => \N__25227\,
            I => \bfn_8_14_0_\
        );

    \I__3869\ : InMux
    port map (
            O => \N__25224\,
            I => \N__25220\
        );

    \I__3868\ : CascadeMux
    port map (
            O => \N__25223\,
            I => \N__25217\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__25220\,
            I => \N__25214\
        );

    \I__3866\ : InMux
    port map (
            O => \N__25217\,
            I => \N__25211\
        );

    \I__3865\ : Span4Mux_h
    port map (
            O => \N__25214\,
            I => \N__25208\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__25211\,
            I => \N__25205\
        );

    \I__3863\ : Span4Mux_v
    port map (
            O => \N__25208\,
            I => \N__25202\
        );

    \I__3862\ : Span4Mux_h
    port map (
            O => \N__25205\,
            I => \N__25199\
        );

    \I__3861\ : Odrv4
    port map (
            O => \N__25202\,
            I => \current_shift_inst.control_inputZ0Z_9\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__25199\,
            I => \current_shift_inst.control_inputZ0Z_9\
        );

    \I__3859\ : InMux
    port map (
            O => \N__25194\,
            I => \current_shift_inst.control_input_1_cry_8\
        );

    \I__3858\ : InMux
    port map (
            O => \N__25191\,
            I => \N__25187\
        );

    \I__3857\ : InMux
    port map (
            O => \N__25190\,
            I => \N__25184\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__25187\,
            I => \N__25181\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__25184\,
            I => \N__25178\
        );

    \I__3854\ : Span4Mux_h
    port map (
            O => \N__25181\,
            I => \N__25175\
        );

    \I__3853\ : Odrv12
    port map (
            O => \N__25178\,
            I => \current_shift_inst.control_inputZ0Z_10\
        );

    \I__3852\ : Odrv4
    port map (
            O => \N__25175\,
            I => \current_shift_inst.control_inputZ0Z_10\
        );

    \I__3851\ : InMux
    port map (
            O => \N__25170\,
            I => \current_shift_inst.control_input_1_cry_9\
        );

    \I__3850\ : InMux
    port map (
            O => \N__25167\,
            I => \N__25163\
        );

    \I__3849\ : InMux
    port map (
            O => \N__25166\,
            I => \N__25160\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__25163\,
            I => \N__25157\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__25160\,
            I => \N__25154\
        );

    \I__3846\ : Span4Mux_v
    port map (
            O => \N__25157\,
            I => \N__25149\
        );

    \I__3845\ : Span4Mux_v
    port map (
            O => \N__25154\,
            I => \N__25149\
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__25149\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__3843\ : InMux
    port map (
            O => \N__25146\,
            I => \current_shift_inst.control_input_1_cry_10\
        );

    \I__3842\ : InMux
    port map (
            O => \N__25143\,
            I => \N__25140\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__25140\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31\
        );

    \I__3840\ : InMux
    port map (
            O => \N__25137\,
            I => \N__25134\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__25134\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31\
        );

    \I__3838\ : CascadeMux
    port map (
            O => \N__25131\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31_cascade_\
        );

    \I__3837\ : InMux
    port map (
            O => \N__25128\,
            I => \N__25125\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__25125\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31\
        );

    \I__3835\ : InMux
    port map (
            O => \N__25122\,
            I => \N__25118\
        );

    \I__3834\ : InMux
    port map (
            O => \N__25121\,
            I => \N__25115\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__25118\,
            I => \current_shift_inst.PI_CTRL.N_47_21\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__25115\,
            I => \current_shift_inst.PI_CTRL.N_47_21\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__25110\,
            I => \N__25107\
        );

    \I__3830\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25104\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__25104\,
            I => \N__25101\
        );

    \I__3828\ : Span4Mux_v
    port map (
            O => \N__25101\,
            I => \N__25098\
        );

    \I__3827\ : Span4Mux_h
    port map (
            O => \N__25098\,
            I => \N__25095\
        );

    \I__3826\ : Odrv4
    port map (
            O => \N__25095\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__25092\,
            I => \N__25089\
        );

    \I__3824\ : InMux
    port map (
            O => \N__25089\,
            I => \N__25086\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__25086\,
            I => \N__25083\
        );

    \I__3822\ : Span4Mux_h
    port map (
            O => \N__25083\,
            I => \N__25080\
        );

    \I__3821\ : Odrv4
    port map (
            O => \N__25080\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__25077\,
            I => \N__25073\
        );

    \I__3819\ : CascadeMux
    port map (
            O => \N__25076\,
            I => \N__25070\
        );

    \I__3818\ : InMux
    port map (
            O => \N__25073\,
            I => \N__25067\
        );

    \I__3817\ : InMux
    port map (
            O => \N__25070\,
            I => \N__25064\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__25067\,
            I => \N__25061\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__25064\,
            I => \N__25058\
        );

    \I__3814\ : Span4Mux_v
    port map (
            O => \N__25061\,
            I => \N__25053\
        );

    \I__3813\ : Span4Mux_h
    port map (
            O => \N__25058\,
            I => \N__25050\
        );

    \I__3812\ : InMux
    port map (
            O => \N__25057\,
            I => \N__25045\
        );

    \I__3811\ : InMux
    port map (
            O => \N__25056\,
            I => \N__25045\
        );

    \I__3810\ : Span4Mux_h
    port map (
            O => \N__25053\,
            I => \N__25040\
        );

    \I__3809\ : Span4Mux_h
    port map (
            O => \N__25050\,
            I => \N__25040\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__25045\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__25040\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3806\ : InMux
    port map (
            O => \N__25035\,
            I => \N__25031\
        );

    \I__3805\ : InMux
    port map (
            O => \N__25034\,
            I => \N__25028\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__25031\,
            I => \N__25018\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__25028\,
            I => \N__25018\
        );

    \I__3802\ : InMux
    port map (
            O => \N__25027\,
            I => \N__25009\
        );

    \I__3801\ : InMux
    port map (
            O => \N__25026\,
            I => \N__25009\
        );

    \I__3800\ : InMux
    port map (
            O => \N__25025\,
            I => \N__25009\
        );

    \I__3799\ : InMux
    port map (
            O => \N__25024\,
            I => \N__25009\
        );

    \I__3798\ : InMux
    port map (
            O => \N__25023\,
            I => \N__25006\
        );

    \I__3797\ : Span4Mux_v
    port map (
            O => \N__25018\,
            I => \N__24994\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__25009\,
            I => \N__24994\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__25006\,
            I => \N__24994\
        );

    \I__3794\ : InMux
    port map (
            O => \N__25005\,
            I => \N__24983\
        );

    \I__3793\ : InMux
    port map (
            O => \N__25004\,
            I => \N__24983\
        );

    \I__3792\ : InMux
    port map (
            O => \N__25003\,
            I => \N__24983\
        );

    \I__3791\ : InMux
    port map (
            O => \N__25002\,
            I => \N__24983\
        );

    \I__3790\ : InMux
    port map (
            O => \N__25001\,
            I => \N__24983\
        );

    \I__3789\ : Span4Mux_v
    port map (
            O => \N__24994\,
            I => \N__24964\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__24983\,
            I => \N__24964\
        );

    \I__3787\ : InMux
    port map (
            O => \N__24982\,
            I => \N__24951\
        );

    \I__3786\ : InMux
    port map (
            O => \N__24981\,
            I => \N__24951\
        );

    \I__3785\ : InMux
    port map (
            O => \N__24980\,
            I => \N__24951\
        );

    \I__3784\ : InMux
    port map (
            O => \N__24979\,
            I => \N__24951\
        );

    \I__3783\ : InMux
    port map (
            O => \N__24978\,
            I => \N__24951\
        );

    \I__3782\ : InMux
    port map (
            O => \N__24977\,
            I => \N__24951\
        );

    \I__3781\ : InMux
    port map (
            O => \N__24976\,
            I => \N__24936\
        );

    \I__3780\ : InMux
    port map (
            O => \N__24975\,
            I => \N__24936\
        );

    \I__3779\ : InMux
    port map (
            O => \N__24974\,
            I => \N__24936\
        );

    \I__3778\ : InMux
    port map (
            O => \N__24973\,
            I => \N__24936\
        );

    \I__3777\ : InMux
    port map (
            O => \N__24972\,
            I => \N__24936\
        );

    \I__3776\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24936\
        );

    \I__3775\ : InMux
    port map (
            O => \N__24970\,
            I => \N__24931\
        );

    \I__3774\ : InMux
    port map (
            O => \N__24969\,
            I => \N__24931\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__24964\,
            I => \N__24928\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__24951\,
            I => \N__24925\
        );

    \I__3771\ : InMux
    port map (
            O => \N__24950\,
            I => \N__24920\
        );

    \I__3770\ : InMux
    port map (
            O => \N__24949\,
            I => \N__24920\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__24936\,
            I => \N__24915\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__24931\,
            I => \N__24915\
        );

    \I__3767\ : Odrv4
    port map (
            O => \N__24928\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3766\ : Odrv12
    port map (
            O => \N__24925\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__24920\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3764\ : Odrv4
    port map (
            O => \N__24915\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3763\ : InMux
    port map (
            O => \N__24906\,
            I => \N__24903\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__24903\,
            I => \N__24900\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__24900\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__3760\ : CascadeMux
    port map (
            O => \N__24897\,
            I => \N__24882\
        );

    \I__3759\ : CascadeMux
    port map (
            O => \N__24896\,
            I => \N__24879\
        );

    \I__3758\ : CascadeMux
    port map (
            O => \N__24895\,
            I => \N__24876\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__24894\,
            I => \N__24873\
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__24893\,
            I => \N__24868\
        );

    \I__3755\ : CascadeMux
    port map (
            O => \N__24892\,
            I => \N__24864\
        );

    \I__3754\ : CascadeMux
    port map (
            O => \N__24891\,
            I => \N__24861\
        );

    \I__3753\ : CascadeMux
    port map (
            O => \N__24890\,
            I => \N__24858\
        );

    \I__3752\ : CascadeMux
    port map (
            O => \N__24889\,
            I => \N__24855\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__24888\,
            I => \N__24852\
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__24887\,
            I => \N__24847\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__24886\,
            I => \N__24844\
        );

    \I__3748\ : CascadeMux
    port map (
            O => \N__24885\,
            I => \N__24841\
        );

    \I__3747\ : InMux
    port map (
            O => \N__24882\,
            I => \N__24829\
        );

    \I__3746\ : InMux
    port map (
            O => \N__24879\,
            I => \N__24829\
        );

    \I__3745\ : InMux
    port map (
            O => \N__24876\,
            I => \N__24829\
        );

    \I__3744\ : InMux
    port map (
            O => \N__24873\,
            I => \N__24829\
        );

    \I__3743\ : InMux
    port map (
            O => \N__24872\,
            I => \N__24829\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__24871\,
            I => \N__24825\
        );

    \I__3741\ : InMux
    port map (
            O => \N__24868\,
            I => \N__24815\
        );

    \I__3740\ : InMux
    port map (
            O => \N__24867\,
            I => \N__24812\
        );

    \I__3739\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24809\
        );

    \I__3738\ : InMux
    port map (
            O => \N__24861\,
            I => \N__24804\
        );

    \I__3737\ : InMux
    port map (
            O => \N__24858\,
            I => \N__24804\
        );

    \I__3736\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24795\
        );

    \I__3735\ : InMux
    port map (
            O => \N__24852\,
            I => \N__24795\
        );

    \I__3734\ : InMux
    port map (
            O => \N__24851\,
            I => \N__24795\
        );

    \I__3733\ : InMux
    port map (
            O => \N__24850\,
            I => \N__24795\
        );

    \I__3732\ : InMux
    port map (
            O => \N__24847\,
            I => \N__24786\
        );

    \I__3731\ : InMux
    port map (
            O => \N__24844\,
            I => \N__24786\
        );

    \I__3730\ : InMux
    port map (
            O => \N__24841\,
            I => \N__24786\
        );

    \I__3729\ : InMux
    port map (
            O => \N__24840\,
            I => \N__24786\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__24829\,
            I => \N__24783\
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__24828\,
            I => \N__24779\
        );

    \I__3726\ : InMux
    port map (
            O => \N__24825\,
            I => \N__24775\
        );

    \I__3725\ : InMux
    port map (
            O => \N__24824\,
            I => \N__24770\
        );

    \I__3724\ : InMux
    port map (
            O => \N__24823\,
            I => \N__24770\
        );

    \I__3723\ : CascadeMux
    port map (
            O => \N__24822\,
            I => \N__24767\
        );

    \I__3722\ : CascadeMux
    port map (
            O => \N__24821\,
            I => \N__24763\
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__24820\,
            I => \N__24760\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__24819\,
            I => \N__24757\
        );

    \I__3719\ : CascadeMux
    port map (
            O => \N__24818\,
            I => \N__24754\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__24815\,
            I => \N__24749\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__24812\,
            I => \N__24746\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24739\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__24804\,
            I => \N__24739\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__24795\,
            I => \N__24739\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__24786\,
            I => \N__24734\
        );

    \I__3712\ : Span4Mux_h
    port map (
            O => \N__24783\,
            I => \N__24734\
        );

    \I__3711\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24731\
        );

    \I__3710\ : InMux
    port map (
            O => \N__24779\,
            I => \N__24726\
        );

    \I__3709\ : InMux
    port map (
            O => \N__24778\,
            I => \N__24726\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__24775\,
            I => \N__24723\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__24770\,
            I => \N__24720\
        );

    \I__3706\ : InMux
    port map (
            O => \N__24767\,
            I => \N__24715\
        );

    \I__3705\ : InMux
    port map (
            O => \N__24766\,
            I => \N__24715\
        );

    \I__3704\ : InMux
    port map (
            O => \N__24763\,
            I => \N__24702\
        );

    \I__3703\ : InMux
    port map (
            O => \N__24760\,
            I => \N__24702\
        );

    \I__3702\ : InMux
    port map (
            O => \N__24757\,
            I => \N__24702\
        );

    \I__3701\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24702\
        );

    \I__3700\ : InMux
    port map (
            O => \N__24753\,
            I => \N__24702\
        );

    \I__3699\ : InMux
    port map (
            O => \N__24752\,
            I => \N__24702\
        );

    \I__3698\ : Span4Mux_h
    port map (
            O => \N__24749\,
            I => \N__24699\
        );

    \I__3697\ : Span4Mux_v
    port map (
            O => \N__24746\,
            I => \N__24690\
        );

    \I__3696\ : Span4Mux_v
    port map (
            O => \N__24739\,
            I => \N__24690\
        );

    \I__3695\ : Span4Mux_v
    port map (
            O => \N__24734\,
            I => \N__24690\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__24731\,
            I => \N__24690\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__24726\,
            I => \N__24683\
        );

    \I__3692\ : Span4Mux_h
    port map (
            O => \N__24723\,
            I => \N__24683\
        );

    \I__3691\ : Span4Mux_h
    port map (
            O => \N__24720\,
            I => \N__24683\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__24715\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__24702\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3688\ : Odrv4
    port map (
            O => \N__24699\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3687\ : Odrv4
    port map (
            O => \N__24690\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__24683\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3685\ : InMux
    port map (
            O => \N__24672\,
            I => \N__24667\
        );

    \I__3684\ : InMux
    port map (
            O => \N__24671\,
            I => \N__24664\
        );

    \I__3683\ : CascadeMux
    port map (
            O => \N__24670\,
            I => \N__24642\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__24667\,
            I => \N__24636\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__24664\,
            I => \N__24636\
        );

    \I__3680\ : InMux
    port map (
            O => \N__24663\,
            I => \N__24627\
        );

    \I__3679\ : InMux
    port map (
            O => \N__24662\,
            I => \N__24627\
        );

    \I__3678\ : InMux
    port map (
            O => \N__24661\,
            I => \N__24627\
        );

    \I__3677\ : InMux
    port map (
            O => \N__24660\,
            I => \N__24627\
        );

    \I__3676\ : InMux
    port map (
            O => \N__24659\,
            I => \N__24624\
        );

    \I__3675\ : InMux
    port map (
            O => \N__24658\,
            I => \N__24611\
        );

    \I__3674\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24611\
        );

    \I__3673\ : InMux
    port map (
            O => \N__24656\,
            I => \N__24611\
        );

    \I__3672\ : InMux
    port map (
            O => \N__24655\,
            I => \N__24611\
        );

    \I__3671\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24611\
        );

    \I__3670\ : InMux
    port map (
            O => \N__24653\,
            I => \N__24611\
        );

    \I__3669\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24606\
        );

    \I__3668\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24606\
        );

    \I__3667\ : InMux
    port map (
            O => \N__24650\,
            I => \N__24588\
        );

    \I__3666\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24588\
        );

    \I__3665\ : InMux
    port map (
            O => \N__24648\,
            I => \N__24588\
        );

    \I__3664\ : InMux
    port map (
            O => \N__24647\,
            I => \N__24588\
        );

    \I__3663\ : InMux
    port map (
            O => \N__24646\,
            I => \N__24588\
        );

    \I__3662\ : InMux
    port map (
            O => \N__24645\,
            I => \N__24588\
        );

    \I__3661\ : InMux
    port map (
            O => \N__24642\,
            I => \N__24583\
        );

    \I__3660\ : InMux
    port map (
            O => \N__24641\,
            I => \N__24583\
        );

    \I__3659\ : Span4Mux_v
    port map (
            O => \N__24636\,
            I => \N__24574\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__24627\,
            I => \N__24574\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__24624\,
            I => \N__24574\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__24611\,
            I => \N__24574\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__24606\,
            I => \N__24571\
        );

    \I__3654\ : InMux
    port map (
            O => \N__24605\,
            I => \N__24560\
        );

    \I__3653\ : InMux
    port map (
            O => \N__24604\,
            I => \N__24560\
        );

    \I__3652\ : InMux
    port map (
            O => \N__24603\,
            I => \N__24560\
        );

    \I__3651\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24560\
        );

    \I__3650\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24560\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__24588\,
            I => \N__24557\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__24583\,
            I => \N__24554\
        );

    \I__3647\ : Span4Mux_v
    port map (
            O => \N__24574\,
            I => \N__24547\
        );

    \I__3646\ : Span4Mux_v
    port map (
            O => \N__24571\,
            I => \N__24547\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__24560\,
            I => \N__24547\
        );

    \I__3644\ : Odrv12
    port map (
            O => \N__24557\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__3643\ : Odrv4
    port map (
            O => \N__24554\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__3642\ : Odrv4
    port map (
            O => \N__24547\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__3641\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24537\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__24537\,
            I => \N__24531\
        );

    \I__3639\ : InMux
    port map (
            O => \N__24536\,
            I => \N__24528\
        );

    \I__3638\ : InMux
    port map (
            O => \N__24535\,
            I => \N__24523\
        );

    \I__3637\ : InMux
    port map (
            O => \N__24534\,
            I => \N__24523\
        );

    \I__3636\ : Span4Mux_v
    port map (
            O => \N__24531\,
            I => \N__24518\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__24528\,
            I => \N__24518\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__24523\,
            I => \N__24515\
        );

    \I__3633\ : Odrv4
    port map (
            O => \N__24518\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__24515\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3631\ : CEMux
    port map (
            O => \N__24510\,
            I => \N__24503\
        );

    \I__3630\ : CEMux
    port map (
            O => \N__24509\,
            I => \N__24496\
        );

    \I__3629\ : CEMux
    port map (
            O => \N__24508\,
            I => \N__24493\
        );

    \I__3628\ : CEMux
    port map (
            O => \N__24507\,
            I => \N__24489\
        );

    \I__3627\ : CEMux
    port map (
            O => \N__24506\,
            I => \N__24486\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__24503\,
            I => \N__24480\
        );

    \I__3625\ : CEMux
    port map (
            O => \N__24502\,
            I => \N__24477\
        );

    \I__3624\ : CEMux
    port map (
            O => \N__24501\,
            I => \N__24472\
        );

    \I__3623\ : CEMux
    port map (
            O => \N__24500\,
            I => \N__24469\
        );

    \I__3622\ : CEMux
    port map (
            O => \N__24499\,
            I => \N__24462\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__24496\,
            I => \N__24459\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__24493\,
            I => \N__24456\
        );

    \I__3619\ : CEMux
    port map (
            O => \N__24492\,
            I => \N__24453\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__24489\,
            I => \N__24450\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__24486\,
            I => \N__24447\
        );

    \I__3616\ : CEMux
    port map (
            O => \N__24485\,
            I => \N__24444\
        );

    \I__3615\ : CEMux
    port map (
            O => \N__24484\,
            I => \N__24441\
        );

    \I__3614\ : CEMux
    port map (
            O => \N__24483\,
            I => \N__24438\
        );

    \I__3613\ : Span4Mux_s3_h
    port map (
            O => \N__24480\,
            I => \N__24433\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__24477\,
            I => \N__24433\
        );

    \I__3611\ : CEMux
    port map (
            O => \N__24476\,
            I => \N__24430\
        );

    \I__3610\ : CEMux
    port map (
            O => \N__24475\,
            I => \N__24427\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__24472\,
            I => \N__24424\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__24469\,
            I => \N__24421\
        );

    \I__3607\ : CEMux
    port map (
            O => \N__24468\,
            I => \N__24418\
        );

    \I__3606\ : CEMux
    port map (
            O => \N__24467\,
            I => \N__24415\
        );

    \I__3605\ : CEMux
    port map (
            O => \N__24466\,
            I => \N__24412\
        );

    \I__3604\ : CEMux
    port map (
            O => \N__24465\,
            I => \N__24408\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__24462\,
            I => \N__24404\
        );

    \I__3602\ : Span4Mux_v
    port map (
            O => \N__24459\,
            I => \N__24397\
        );

    \I__3601\ : Span4Mux_v
    port map (
            O => \N__24456\,
            I => \N__24397\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__24453\,
            I => \N__24397\
        );

    \I__3599\ : Span4Mux_h
    port map (
            O => \N__24450\,
            I => \N__24394\
        );

    \I__3598\ : Span4Mux_h
    port map (
            O => \N__24447\,
            I => \N__24391\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__24444\,
            I => \N__24388\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__24441\,
            I => \N__24385\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__24438\,
            I => \N__24382\
        );

    \I__3594\ : Span4Mux_h
    port map (
            O => \N__24433\,
            I => \N__24377\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__24430\,
            I => \N__24377\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__24427\,
            I => \N__24374\
        );

    \I__3591\ : Span4Mux_h
    port map (
            O => \N__24424\,
            I => \N__24371\
        );

    \I__3590\ : Span4Mux_s3_h
    port map (
            O => \N__24421\,
            I => \N__24366\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__24418\,
            I => \N__24366\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__24415\,
            I => \N__24363\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__24412\,
            I => \N__24360\
        );

    \I__3586\ : CEMux
    port map (
            O => \N__24411\,
            I => \N__24357\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__24408\,
            I => \N__24354\
        );

    \I__3584\ : CEMux
    port map (
            O => \N__24407\,
            I => \N__24351\
        );

    \I__3583\ : Span4Mux_h
    port map (
            O => \N__24404\,
            I => \N__24348\
        );

    \I__3582\ : Span4Mux_v
    port map (
            O => \N__24397\,
            I => \N__24345\
        );

    \I__3581\ : Span4Mux_v
    port map (
            O => \N__24394\,
            I => \N__24336\
        );

    \I__3580\ : Span4Mux_v
    port map (
            O => \N__24391\,
            I => \N__24336\
        );

    \I__3579\ : Span4Mux_h
    port map (
            O => \N__24388\,
            I => \N__24336\
        );

    \I__3578\ : Span4Mux_h
    port map (
            O => \N__24385\,
            I => \N__24336\
        );

    \I__3577\ : Span4Mux_s3_h
    port map (
            O => \N__24382\,
            I => \N__24333\
        );

    \I__3576\ : Span4Mux_v
    port map (
            O => \N__24377\,
            I => \N__24328\
        );

    \I__3575\ : Span4Mux_h
    port map (
            O => \N__24374\,
            I => \N__24328\
        );

    \I__3574\ : Span4Mux_v
    port map (
            O => \N__24371\,
            I => \N__24317\
        );

    \I__3573\ : Span4Mux_h
    port map (
            O => \N__24366\,
            I => \N__24317\
        );

    \I__3572\ : Span4Mux_h
    port map (
            O => \N__24363\,
            I => \N__24317\
        );

    \I__3571\ : Span4Mux_h
    port map (
            O => \N__24360\,
            I => \N__24317\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__24357\,
            I => \N__24317\
        );

    \I__3569\ : Span4Mux_s3_h
    port map (
            O => \N__24354\,
            I => \N__24312\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__24351\,
            I => \N__24312\
        );

    \I__3567\ : Sp12to4
    port map (
            O => \N__24348\,
            I => \N__24309\
        );

    \I__3566\ : Span4Mux_v
    port map (
            O => \N__24345\,
            I => \N__24306\
        );

    \I__3565\ : Span4Mux_v
    port map (
            O => \N__24336\,
            I => \N__24301\
        );

    \I__3564\ : Span4Mux_h
    port map (
            O => \N__24333\,
            I => \N__24301\
        );

    \I__3563\ : Span4Mux_v
    port map (
            O => \N__24328\,
            I => \N__24298\
        );

    \I__3562\ : Span4Mux_v
    port map (
            O => \N__24317\,
            I => \N__24293\
        );

    \I__3561\ : Span4Mux_h
    port map (
            O => \N__24312\,
            I => \N__24293\
        );

    \I__3560\ : Odrv12
    port map (
            O => \N__24309\,
            I => \N_655_g\
        );

    \I__3559\ : Odrv4
    port map (
            O => \N__24306\,
            I => \N_655_g\
        );

    \I__3558\ : Odrv4
    port map (
            O => \N__24301\,
            I => \N_655_g\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__24298\,
            I => \N_655_g\
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__24293\,
            I => \N_655_g\
        );

    \I__3555\ : InMux
    port map (
            O => \N__24282\,
            I => \N__24278\
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__24281\,
            I => \N__24275\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__24278\,
            I => \N__24272\
        );

    \I__3552\ : InMux
    port map (
            O => \N__24275\,
            I => \N__24269\
        );

    \I__3551\ : Span4Mux_v
    port map (
            O => \N__24272\,
            I => \N__24264\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__24269\,
            I => \N__24264\
        );

    \I__3549\ : Span4Mux_h
    port map (
            O => \N__24264\,
            I => \N__24261\
        );

    \I__3548\ : Odrv4
    port map (
            O => \N__24261\,
            I => \current_shift_inst.control_inputZ0Z_0\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__24258\,
            I => \N__24254\
        );

    \I__3546\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24251\
        );

    \I__3545\ : InMux
    port map (
            O => \N__24254\,
            I => \N__24248\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__24251\,
            I => \N__24243\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__24248\,
            I => \N__24243\
        );

    \I__3542\ : Span4Mux_h
    port map (
            O => \N__24243\,
            I => \N__24240\
        );

    \I__3541\ : Odrv4
    port map (
            O => \N__24240\,
            I => \current_shift_inst.control_inputZ0Z_1\
        );

    \I__3540\ : InMux
    port map (
            O => \N__24237\,
            I => \current_shift_inst.control_input_1_cry_0\
        );

    \I__3539\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24230\
        );

    \I__3538\ : CascadeMux
    port map (
            O => \N__24233\,
            I => \N__24227\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__24230\,
            I => \N__24224\
        );

    \I__3536\ : InMux
    port map (
            O => \N__24227\,
            I => \N__24221\
        );

    \I__3535\ : Span4Mux_v
    port map (
            O => \N__24224\,
            I => \N__24216\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__24221\,
            I => \N__24216\
        );

    \I__3533\ : Span4Mux_h
    port map (
            O => \N__24216\,
            I => \N__24213\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__24213\,
            I => \current_shift_inst.control_inputZ0Z_2\
        );

    \I__3531\ : InMux
    port map (
            O => \N__24210\,
            I => \current_shift_inst.control_input_1_cry_1\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__24207\,
            I => \N__24203\
        );

    \I__3529\ : InMux
    port map (
            O => \N__24206\,
            I => \N__24200\
        );

    \I__3528\ : InMux
    port map (
            O => \N__24203\,
            I => \N__24197\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__24200\,
            I => \N__24194\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__24197\,
            I => \N__24191\
        );

    \I__3525\ : Span4Mux_v
    port map (
            O => \N__24194\,
            I => \N__24186\
        );

    \I__3524\ : Span4Mux_v
    port map (
            O => \N__24191\,
            I => \N__24186\
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__24186\,
            I => \current_shift_inst.control_inputZ0Z_3\
        );

    \I__3522\ : InMux
    port map (
            O => \N__24183\,
            I => \current_shift_inst.control_input_1_cry_2\
        );

    \I__3521\ : InMux
    port map (
            O => \N__24180\,
            I => \N__24175\
        );

    \I__3520\ : InMux
    port map (
            O => \N__24179\,
            I => \N__24172\
        );

    \I__3519\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24169\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__24175\,
            I => \N__24166\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__24172\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__24169\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__3515\ : Odrv4
    port map (
            O => \N__24166\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__3514\ : InMux
    port map (
            O => \N__24159\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__3513\ : InMux
    port map (
            O => \N__24156\,
            I => \N__24151\
        );

    \I__3512\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24148\
        );

    \I__3511\ : InMux
    port map (
            O => \N__24154\,
            I => \N__24145\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__24151\,
            I => \N__24142\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__24148\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__24145\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__3507\ : Odrv4
    port map (
            O => \N__24142\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__3506\ : InMux
    port map (
            O => \N__24135\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__3505\ : InMux
    port map (
            O => \N__24132\,
            I => \N__24127\
        );

    \I__3504\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24124\
        );

    \I__3503\ : InMux
    port map (
            O => \N__24130\,
            I => \N__24121\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__24127\,
            I => \N__24118\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__24124\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__24121\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__3499\ : Odrv4
    port map (
            O => \N__24118\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__3498\ : InMux
    port map (
            O => \N__24111\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__3497\ : InMux
    port map (
            O => \N__24108\,
            I => \N__24103\
        );

    \I__3496\ : InMux
    port map (
            O => \N__24107\,
            I => \N__24100\
        );

    \I__3495\ : InMux
    port map (
            O => \N__24106\,
            I => \N__24097\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__24103\,
            I => \N__24094\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__24100\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__24097\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__3491\ : Odrv4
    port map (
            O => \N__24094\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__3490\ : InMux
    port map (
            O => \N__24087\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__3489\ : InMux
    port map (
            O => \N__24084\,
            I => \N__24080\
        );

    \I__3488\ : InMux
    port map (
            O => \N__24083\,
            I => \N__24076\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__24080\,
            I => \N__24073\
        );

    \I__3486\ : InMux
    port map (
            O => \N__24079\,
            I => \N__24070\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__24076\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__3484\ : Odrv4
    port map (
            O => \N__24073\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__24070\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__3482\ : InMux
    port map (
            O => \N__24063\,
            I => \bfn_8_9_0_\
        );

    \I__3481\ : InMux
    port map (
            O => \N__24060\,
            I => \N__24048\
        );

    \I__3480\ : InMux
    port map (
            O => \N__24059\,
            I => \N__24048\
        );

    \I__3479\ : InMux
    port map (
            O => \N__24058\,
            I => \N__24048\
        );

    \I__3478\ : InMux
    port map (
            O => \N__24057\,
            I => \N__24048\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__24048\,
            I => \N__24039\
        );

    \I__3476\ : InMux
    port map (
            O => \N__24047\,
            I => \N__24034\
        );

    \I__3475\ : InMux
    port map (
            O => \N__24046\,
            I => \N__24034\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24045\,
            I => \N__24025\
        );

    \I__3473\ : InMux
    port map (
            O => \N__24044\,
            I => \N__24025\
        );

    \I__3472\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24025\
        );

    \I__3471\ : InMux
    port map (
            O => \N__24042\,
            I => \N__24025\
        );

    \I__3470\ : Odrv4
    port map (
            O => \N__24039\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__24034\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__24025\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__3467\ : InMux
    port map (
            O => \N__24018\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__3466\ : InMux
    port map (
            O => \N__24015\,
            I => \N__24011\
        );

    \I__3465\ : InMux
    port map (
            O => \N__24014\,
            I => \N__24007\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__24004\
        );

    \I__3463\ : InMux
    port map (
            O => \N__24010\,
            I => \N__24001\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__24007\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__24004\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__24001\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__3459\ : InMux
    port map (
            O => \N__23994\,
            I => \N__23990\
        );

    \I__3458\ : InMux
    port map (
            O => \N__23993\,
            I => \N__23987\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__23990\,
            I => \N__23984\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__23987\,
            I => \N__23981\
        );

    \I__3455\ : Odrv4
    port map (
            O => \N__23984\,
            I => \current_shift_inst.PI_CTRL.N_47_16\
        );

    \I__3454\ : Odrv4
    port map (
            O => \N__23981\,
            I => \current_shift_inst.PI_CTRL.N_47_16\
        );

    \I__3453\ : InMux
    port map (
            O => \N__23976\,
            I => \N__23972\
        );

    \I__3452\ : InMux
    port map (
            O => \N__23975\,
            I => \N__23969\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__23972\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__23969\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__3449\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23958\
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__23963\,
            I => \N__23955\
        );

    \I__3447\ : CascadeMux
    port map (
            O => \N__23962\,
            I => \N__23952\
        );

    \I__3446\ : InMux
    port map (
            O => \N__23961\,
            I => \N__23948\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__23958\,
            I => \N__23945\
        );

    \I__3444\ : InMux
    port map (
            O => \N__23955\,
            I => \N__23941\
        );

    \I__3443\ : InMux
    port map (
            O => \N__23952\,
            I => \N__23936\
        );

    \I__3442\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23936\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__23948\,
            I => \N__23933\
        );

    \I__3440\ : Span4Mux_v
    port map (
            O => \N__23945\,
            I => \N__23930\
        );

    \I__3439\ : InMux
    port map (
            O => \N__23944\,
            I => \N__23927\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__23941\,
            I => \N__23922\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__23936\,
            I => \N__23922\
        );

    \I__3436\ : Span4Mux_h
    port map (
            O => \N__23933\,
            I => \N__23915\
        );

    \I__3435\ : Span4Mux_h
    port map (
            O => \N__23930\,
            I => \N__23915\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__23927\,
            I => \N__23915\
        );

    \I__3433\ : Span4Mux_h
    port map (
            O => \N__23922\,
            I => \N__23912\
        );

    \I__3432\ : Span4Mux_v
    port map (
            O => \N__23915\,
            I => \N__23909\
        );

    \I__3431\ : Odrv4
    port map (
            O => \N__23912\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3430\ : Odrv4
    port map (
            O => \N__23909\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3429\ : CascadeMux
    port map (
            O => \N__23904\,
            I => \N__23899\
        );

    \I__3428\ : InMux
    port map (
            O => \N__23903\,
            I => \N__23895\
        );

    \I__3427\ : InMux
    port map (
            O => \N__23902\,
            I => \N__23892\
        );

    \I__3426\ : InMux
    port map (
            O => \N__23899\,
            I => \N__23889\
        );

    \I__3425\ : CascadeMux
    port map (
            O => \N__23898\,
            I => \N__23886\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__23895\,
            I => \N__23883\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__23892\,
            I => \N__23880\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__23889\,
            I => \N__23877\
        );

    \I__3421\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23874\
        );

    \I__3420\ : Span12Mux_v
    port map (
            O => \N__23883\,
            I => \N__23871\
        );

    \I__3419\ : Span4Mux_v
    port map (
            O => \N__23880\,
            I => \N__23868\
        );

    \I__3418\ : Odrv4
    port map (
            O => \N__23877\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__23874\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__3416\ : Odrv12
    port map (
            O => \N__23871\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__3415\ : Odrv4
    port map (
            O => \N__23868\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__3414\ : InMux
    port map (
            O => \N__23859\,
            I => \N__23856\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__23856\,
            I => \N__23850\
        );

    \I__3412\ : InMux
    port map (
            O => \N__23855\,
            I => \N__23847\
        );

    \I__3411\ : InMux
    port map (
            O => \N__23854\,
            I => \N__23844\
        );

    \I__3410\ : InMux
    port map (
            O => \N__23853\,
            I => \N__23841\
        );

    \I__3409\ : Span4Mux_v
    port map (
            O => \N__23850\,
            I => \N__23836\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__23847\,
            I => \N__23836\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__23844\,
            I => \N__23833\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__23841\,
            I => \N__23830\
        );

    \I__3405\ : Odrv4
    port map (
            O => \N__23836\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3404\ : Odrv4
    port map (
            O => \N__23833\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3403\ : Odrv4
    port map (
            O => \N__23830\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__23823\,
            I => \N__23819\
        );

    \I__3401\ : InMux
    port map (
            O => \N__23822\,
            I => \N__23815\
        );

    \I__3400\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23812\
        );

    \I__3399\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23809\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__23815\,
            I => \N__23805\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__23812\,
            I => \N__23800\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__23809\,
            I => \N__23800\
        );

    \I__3395\ : InMux
    port map (
            O => \N__23808\,
            I => \N__23797\
        );

    \I__3394\ : Span4Mux_v
    port map (
            O => \N__23805\,
            I => \N__23792\
        );

    \I__3393\ : Span4Mux_v
    port map (
            O => \N__23800\,
            I => \N__23792\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__23797\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__23792\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__23787\,
            I => \N__23784\
        );

    \I__3389\ : InMux
    port map (
            O => \N__23784\,
            I => \N__23780\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__23783\,
            I => \N__23776\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__23780\,
            I => \N__23772\
        );

    \I__3386\ : InMux
    port map (
            O => \N__23779\,
            I => \N__23769\
        );

    \I__3385\ : InMux
    port map (
            O => \N__23776\,
            I => \N__23766\
        );

    \I__3384\ : InMux
    port map (
            O => \N__23775\,
            I => \N__23763\
        );

    \I__3383\ : Span4Mux_v
    port map (
            O => \N__23772\,
            I => \N__23758\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__23769\,
            I => \N__23758\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__23766\,
            I => \N__23755\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__23763\,
            I => \N__23752\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__23758\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3378\ : Odrv4
    port map (
            O => \N__23755\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3377\ : Odrv4
    port map (
            O => \N__23752\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3376\ : InMux
    port map (
            O => \N__23745\,
            I => \N__23742\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__23742\,
            I => \N__23739\
        );

    \I__3374\ : Span4Mux_v
    port map (
            O => \N__23739\,
            I => \N__23736\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__23736\,
            I => \pwm_generator_inst.thresholdZ0Z_7\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__23733\,
            I => \N__23730\
        );

    \I__3371\ : InMux
    port map (
            O => \N__23730\,
            I => \N__23727\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__23727\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__23724\,
            I => \N__23721\
        );

    \I__3368\ : InMux
    port map (
            O => \N__23721\,
            I => \N__23718\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__23718\,
            I => \N__23715\
        );

    \I__3366\ : Odrv4
    port map (
            O => \N__23715\,
            I => \pwm_generator_inst.thresholdZ0Z_8\
        );

    \I__3365\ : InMux
    port map (
            O => \N__23712\,
            I => \N__23709\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__23709\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__3363\ : CascadeMux
    port map (
            O => \N__23706\,
            I => \N__23703\
        );

    \I__3362\ : InMux
    port map (
            O => \N__23703\,
            I => \N__23700\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__23700\,
            I => \N__23697\
        );

    \I__3360\ : Span4Mux_v
    port map (
            O => \N__23697\,
            I => \N__23694\
        );

    \I__3359\ : Odrv4
    port map (
            O => \N__23694\,
            I => \pwm_generator_inst.thresholdZ0Z_9\
        );

    \I__3358\ : InMux
    port map (
            O => \N__23691\,
            I => \N__23688\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__23688\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__3356\ : InMux
    port map (
            O => \N__23685\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__3355\ : IoInMux
    port map (
            O => \N__23682\,
            I => \N__23679\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__23679\,
            I => \N__23676\
        );

    \I__3353\ : IoSpan4Mux
    port map (
            O => \N__23676\,
            I => \N__23673\
        );

    \I__3352\ : Span4Mux_s2_v
    port map (
            O => \N__23673\,
            I => \N__23670\
        );

    \I__3351\ : Span4Mux_v
    port map (
            O => \N__23670\,
            I => \N__23667\
        );

    \I__3350\ : Span4Mux_h
    port map (
            O => \N__23667\,
            I => \N__23664\
        );

    \I__3349\ : Span4Mux_h
    port map (
            O => \N__23664\,
            I => \N__23661\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__23661\,
            I => pwm_output_c
        );

    \I__3347\ : InMux
    port map (
            O => \N__23658\,
            I => \N__23654\
        );

    \I__3346\ : InMux
    port map (
            O => \N__23657\,
            I => \N__23650\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__23654\,
            I => \N__23647\
        );

    \I__3344\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23644\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__23650\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3342\ : Odrv4
    port map (
            O => \N__23647\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__23644\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3340\ : InMux
    port map (
            O => \N__23637\,
            I => \bfn_8_8_0_\
        );

    \I__3339\ : InMux
    port map (
            O => \N__23634\,
            I => \N__23629\
        );

    \I__3338\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23626\
        );

    \I__3337\ : InMux
    port map (
            O => \N__23632\,
            I => \N__23623\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__23629\,
            I => \N__23620\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__23626\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__23623\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__3333\ : Odrv4
    port map (
            O => \N__23620\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__3332\ : InMux
    port map (
            O => \N__23613\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__3331\ : InMux
    port map (
            O => \N__23610\,
            I => \N__23606\
        );

    \I__3330\ : InMux
    port map (
            O => \N__23609\,
            I => \N__23602\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__23606\,
            I => \N__23599\
        );

    \I__3328\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23596\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__23602\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__3326\ : Odrv4
    port map (
            O => \N__23599\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__23596\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__3324\ : InMux
    port map (
            O => \N__23589\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__3323\ : InMux
    port map (
            O => \N__23586\,
            I => \N__23581\
        );

    \I__3322\ : InMux
    port map (
            O => \N__23585\,
            I => \N__23578\
        );

    \I__3321\ : InMux
    port map (
            O => \N__23584\,
            I => \N__23575\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__23581\,
            I => \N__23572\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__23578\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__23575\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__3317\ : Odrv4
    port map (
            O => \N__23572\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__3316\ : InMux
    port map (
            O => \N__23565\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__3315\ : InMux
    port map (
            O => \N__23562\,
            I => \N__23559\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__23559\,
            I => \N__23556\
        );

    \I__3313\ : Odrv12
    port map (
            O => \N__23556\,
            I => il_max_comp1_c
        );

    \I__3312\ : CascadeMux
    port map (
            O => \N__23553\,
            I => \N__23550\
        );

    \I__3311\ : InMux
    port map (
            O => \N__23550\,
            I => \N__23547\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__23547\,
            I => \N__23544\
        );

    \I__3309\ : Span4Mux_v
    port map (
            O => \N__23544\,
            I => \N__23541\
        );

    \I__3308\ : Span4Mux_h
    port map (
            O => \N__23541\,
            I => \N__23538\
        );

    \I__3307\ : Odrv4
    port map (
            O => \N__23538\,
            I => \pwm_generator_inst.thresholdZ0Z_0\
        );

    \I__3306\ : InMux
    port map (
            O => \N__23535\,
            I => \N__23532\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__23532\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__23529\,
            I => \N__23526\
        );

    \I__3303\ : InMux
    port map (
            O => \N__23526\,
            I => \N__23523\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__23523\,
            I => \pwm_generator_inst.thresholdZ0Z_1\
        );

    \I__3301\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23517\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__23517\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__3299\ : CascadeMux
    port map (
            O => \N__23514\,
            I => \N__23511\
        );

    \I__3298\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23508\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__23508\,
            I => \N__23505\
        );

    \I__3296\ : Odrv4
    port map (
            O => \N__23505\,
            I => \pwm_generator_inst.thresholdZ0Z_2\
        );

    \I__3295\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23499\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__23499\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__3293\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23493\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__23493\,
            I => \N__23490\
        );

    \I__3291\ : Span4Mux_h
    port map (
            O => \N__23490\,
            I => \N__23487\
        );

    \I__3290\ : Odrv4
    port map (
            O => \N__23487\,
            I => \pwm_generator_inst.thresholdZ0Z_3\
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__23484\,
            I => \N__23481\
        );

    \I__3288\ : InMux
    port map (
            O => \N__23481\,
            I => \N__23478\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__23478\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__3286\ : CascadeMux
    port map (
            O => \N__23475\,
            I => \N__23472\
        );

    \I__3285\ : InMux
    port map (
            O => \N__23472\,
            I => \N__23469\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__23469\,
            I => \N__23466\
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__23466\,
            I => \pwm_generator_inst.thresholdZ0Z_4\
        );

    \I__3282\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23460\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__23460\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__23457\,
            I => \N__23454\
        );

    \I__3279\ : InMux
    port map (
            O => \N__23454\,
            I => \N__23451\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__23451\,
            I => \N__23448\
        );

    \I__3277\ : Span4Mux_v
    port map (
            O => \N__23448\,
            I => \N__23445\
        );

    \I__3276\ : Odrv4
    port map (
            O => \N__23445\,
            I => \pwm_generator_inst.thresholdZ0Z_5\
        );

    \I__3275\ : InMux
    port map (
            O => \N__23442\,
            I => \N__23439\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__23439\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__23436\,
            I => \N__23433\
        );

    \I__3272\ : InMux
    port map (
            O => \N__23433\,
            I => \N__23430\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__23430\,
            I => \N__23427\
        );

    \I__3270\ : Odrv12
    port map (
            O => \N__23427\,
            I => \pwm_generator_inst.thresholdZ0Z_6\
        );

    \I__3269\ : InMux
    port map (
            O => \N__23424\,
            I => \N__23421\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__23421\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__3267\ : InMux
    port map (
            O => \N__23418\,
            I => \current_shift_inst.timer_phase.counter_cry_20\
        );

    \I__3266\ : InMux
    port map (
            O => \N__23415\,
            I => \current_shift_inst.timer_phase.counter_cry_21\
        );

    \I__3265\ : InMux
    port map (
            O => \N__23412\,
            I => \current_shift_inst.timer_phase.counter_cry_22\
        );

    \I__3264\ : InMux
    port map (
            O => \N__23409\,
            I => \bfn_7_22_0_\
        );

    \I__3263\ : InMux
    port map (
            O => \N__23406\,
            I => \current_shift_inst.timer_phase.counter_cry_24\
        );

    \I__3262\ : InMux
    port map (
            O => \N__23403\,
            I => \current_shift_inst.timer_phase.counter_cry_25\
        );

    \I__3261\ : InMux
    port map (
            O => \N__23400\,
            I => \current_shift_inst.timer_phase.counter_cry_26\
        );

    \I__3260\ : InMux
    port map (
            O => \N__23397\,
            I => \current_shift_inst.timer_phase.counter_cry_27\
        );

    \I__3259\ : InMux
    port map (
            O => \N__23394\,
            I => \current_shift_inst.timer_phase.counter_cry_28\
        );

    \I__3258\ : InMux
    port map (
            O => \N__23391\,
            I => \N__23388\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__23388\,
            I => \N__23385\
        );

    \I__3256\ : Span4Mux_h
    port map (
            O => \N__23385\,
            I => \N__23382\
        );

    \I__3255\ : Odrv4
    port map (
            O => \N__23382\,
            I => il_min_comp2_c
        );

    \I__3254\ : InMux
    port map (
            O => \N__23379\,
            I => \current_shift_inst.timer_phase.counter_cry_11\
        );

    \I__3253\ : InMux
    port map (
            O => \N__23376\,
            I => \current_shift_inst.timer_phase.counter_cry_12\
        );

    \I__3252\ : InMux
    port map (
            O => \N__23373\,
            I => \current_shift_inst.timer_phase.counter_cry_13\
        );

    \I__3251\ : InMux
    port map (
            O => \N__23370\,
            I => \current_shift_inst.timer_phase.counter_cry_14\
        );

    \I__3250\ : InMux
    port map (
            O => \N__23367\,
            I => \bfn_7_21_0_\
        );

    \I__3249\ : InMux
    port map (
            O => \N__23364\,
            I => \current_shift_inst.timer_phase.counter_cry_16\
        );

    \I__3248\ : InMux
    port map (
            O => \N__23361\,
            I => \current_shift_inst.timer_phase.counter_cry_17\
        );

    \I__3247\ : InMux
    port map (
            O => \N__23358\,
            I => \current_shift_inst.timer_phase.counter_cry_18\
        );

    \I__3246\ : InMux
    port map (
            O => \N__23355\,
            I => \current_shift_inst.timer_phase.counter_cry_19\
        );

    \I__3245\ : InMux
    port map (
            O => \N__23352\,
            I => \current_shift_inst.timer_phase.counter_cry_2\
        );

    \I__3244\ : InMux
    port map (
            O => \N__23349\,
            I => \current_shift_inst.timer_phase.counter_cry_3\
        );

    \I__3243\ : InMux
    port map (
            O => \N__23346\,
            I => \current_shift_inst.timer_phase.counter_cry_4\
        );

    \I__3242\ : InMux
    port map (
            O => \N__23343\,
            I => \current_shift_inst.timer_phase.counter_cry_5\
        );

    \I__3241\ : InMux
    port map (
            O => \N__23340\,
            I => \current_shift_inst.timer_phase.counter_cry_6\
        );

    \I__3240\ : InMux
    port map (
            O => \N__23337\,
            I => \bfn_7_20_0_\
        );

    \I__3239\ : InMux
    port map (
            O => \N__23334\,
            I => \current_shift_inst.timer_phase.counter_cry_8\
        );

    \I__3238\ : InMux
    port map (
            O => \N__23331\,
            I => \current_shift_inst.timer_phase.counter_cry_9\
        );

    \I__3237\ : InMux
    port map (
            O => \N__23328\,
            I => \current_shift_inst.timer_phase.counter_cry_10\
        );

    \I__3236\ : InMux
    port map (
            O => \N__23325\,
            I => \bfn_7_19_0_\
        );

    \I__3235\ : InMux
    port map (
            O => \N__23322\,
            I => \current_shift_inst.timer_phase.counter_cry_0\
        );

    \I__3234\ : InMux
    port map (
            O => \N__23319\,
            I => \current_shift_inst.timer_phase.counter_cry_1\
        );

    \I__3233\ : CascadeMux
    port map (
            O => \N__23316\,
            I => \N__23313\
        );

    \I__3232\ : InMux
    port map (
            O => \N__23313\,
            I => \N__23310\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__23310\,
            I => \N__23307\
        );

    \I__3230\ : Sp12to4
    port map (
            O => \N__23307\,
            I => \N__23304\
        );

    \I__3229\ : Odrv12
    port map (
            O => \N__23304\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__3228\ : InMux
    port map (
            O => \N__23301\,
            I => \N__23298\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__23298\,
            I => \N__23295\
        );

    \I__3226\ : Odrv12
    port map (
            O => \N__23295\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__3225\ : InMux
    port map (
            O => \N__23292\,
            I => \N__23289\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__23289\,
            I => \N__23284\
        );

    \I__3223\ : InMux
    port map (
            O => \N__23288\,
            I => \N__23281\
        );

    \I__3222\ : CascadeMux
    port map (
            O => \N__23287\,
            I => \N__23277\
        );

    \I__3221\ : Span4Mux_v
    port map (
            O => \N__23284\,
            I => \N__23272\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__23281\,
            I => \N__23272\
        );

    \I__3219\ : InMux
    port map (
            O => \N__23280\,
            I => \N__23267\
        );

    \I__3218\ : InMux
    port map (
            O => \N__23277\,
            I => \N__23267\
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__23272\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__23267\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__3215\ : InMux
    port map (
            O => \N__23262\,
            I => \N__23259\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__23259\,
            I => \N__23254\
        );

    \I__3213\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23251\
        );

    \I__3212\ : InMux
    port map (
            O => \N__23257\,
            I => \N__23247\
        );

    \I__3211\ : Span4Mux_v
    port map (
            O => \N__23254\,
            I => \N__23242\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__23251\,
            I => \N__23242\
        );

    \I__3209\ : InMux
    port map (
            O => \N__23250\,
            I => \N__23239\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__23247\,
            I => \N__23236\
        );

    \I__3207\ : Span4Mux_v
    port map (
            O => \N__23242\,
            I => \N__23233\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__23239\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__3205\ : Odrv12
    port map (
            O => \N__23236\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__23233\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__3203\ : InMux
    port map (
            O => \N__23226\,
            I => \N__23221\
        );

    \I__3202\ : InMux
    port map (
            O => \N__23225\,
            I => \N__23217\
        );

    \I__3201\ : InMux
    port map (
            O => \N__23224\,
            I => \N__23214\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__23221\,
            I => \N__23211\
        );

    \I__3199\ : InMux
    port map (
            O => \N__23220\,
            I => \N__23208\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__23217\,
            I => \N__23205\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__23214\,
            I => \N__23202\
        );

    \I__3196\ : Span4Mux_v
    port map (
            O => \N__23211\,
            I => \N__23195\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__23208\,
            I => \N__23195\
        );

    \I__3194\ : Span4Mux_h
    port map (
            O => \N__23205\,
            I => \N__23195\
        );

    \I__3193\ : Odrv4
    port map (
            O => \N__23202\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__23195\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__23190\,
            I => \N__23185\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__23189\,
            I => \N__23182\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__23188\,
            I => \N__23179\
        );

    \I__3188\ : InMux
    port map (
            O => \N__23185\,
            I => \N__23176\
        );

    \I__3187\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23172\
        );

    \I__3186\ : InMux
    port map (
            O => \N__23179\,
            I => \N__23169\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__23176\,
            I => \N__23166\
        );

    \I__3184\ : InMux
    port map (
            O => \N__23175\,
            I => \N__23163\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__23172\,
            I => \N__23160\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__23169\,
            I => \N__23157\
        );

    \I__3181\ : Span4Mux_v
    port map (
            O => \N__23166\,
            I => \N__23150\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__23163\,
            I => \N__23150\
        );

    \I__3179\ : Span4Mux_h
    port map (
            O => \N__23160\,
            I => \N__23150\
        );

    \I__3178\ : Odrv4
    port map (
            O => \N__23157\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__23150\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3176\ : InMux
    port map (
            O => \N__23145\,
            I => \N__23139\
        );

    \I__3175\ : CascadeMux
    port map (
            O => \N__23144\,
            I => \N__23136\
        );

    \I__3174\ : InMux
    port map (
            O => \N__23143\,
            I => \N__23133\
        );

    \I__3173\ : InMux
    port map (
            O => \N__23142\,
            I => \N__23130\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__23139\,
            I => \N__23127\
        );

    \I__3171\ : InMux
    port map (
            O => \N__23136\,
            I => \N__23124\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__23133\,
            I => \N__23121\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__23130\,
            I => \N__23118\
        );

    \I__3168\ : Span4Mux_v
    port map (
            O => \N__23127\,
            I => \N__23111\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__23124\,
            I => \N__23111\
        );

    \I__3166\ : Span4Mux_h
    port map (
            O => \N__23121\,
            I => \N__23111\
        );

    \I__3165\ : Odrv4
    port map (
            O => \N__23118\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__23111\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__3163\ : InMux
    port map (
            O => \N__23106\,
            I => \N__23101\
        );

    \I__3162\ : InMux
    port map (
            O => \N__23105\,
            I => \N__23095\
        );

    \I__3161\ : InMux
    port map (
            O => \N__23104\,
            I => \N__23095\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__23101\,
            I => \N__23092\
        );

    \I__3159\ : InMux
    port map (
            O => \N__23100\,
            I => \N__23089\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__23095\,
            I => \N__23086\
        );

    \I__3157\ : Odrv12
    port map (
            O => \N__23092\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__23089\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3155\ : Odrv4
    port map (
            O => \N__23086\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3154\ : CascadeMux
    port map (
            O => \N__23079\,
            I => \N__23076\
        );

    \I__3153\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23068\
        );

    \I__3152\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23068\
        );

    \I__3151\ : InMux
    port map (
            O => \N__23074\,
            I => \N__23065\
        );

    \I__3150\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23062\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__23068\,
            I => \N__23059\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__23065\,
            I => \N__23056\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__23062\,
            I => \N__23051\
        );

    \I__3146\ : Span4Mux_h
    port map (
            O => \N__23059\,
            I => \N__23051\
        );

    \I__3145\ : Odrv12
    port map (
            O => \N__23056\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3144\ : Odrv4
    port map (
            O => \N__23051\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3143\ : CascadeMux
    port map (
            O => \N__23046\,
            I => \N__23041\
        );

    \I__3142\ : InMux
    port map (
            O => \N__23045\,
            I => \N__23038\
        );

    \I__3141\ : InMux
    port map (
            O => \N__23044\,
            I => \N__23032\
        );

    \I__3140\ : InMux
    port map (
            O => \N__23041\,
            I => \N__23032\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__23038\,
            I => \N__23029\
        );

    \I__3138\ : InMux
    port map (
            O => \N__23037\,
            I => \N__23026\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__23032\,
            I => \N__23023\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__23029\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__23026\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3134\ : Odrv4
    port map (
            O => \N__23023\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3133\ : InMux
    port map (
            O => \N__23016\,
            I => \N__23012\
        );

    \I__3132\ : InMux
    port map (
            O => \N__23015\,
            I => \N__23009\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__23012\,
            I => \N__23006\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__23009\,
            I => \N__23003\
        );

    \I__3129\ : Odrv12
    port map (
            O => \N__23006\,
            I => \current_shift_inst.PI_CTRL.N_46_16\
        );

    \I__3128\ : Odrv4
    port map (
            O => \N__23003\,
            I => \current_shift_inst.PI_CTRL.N_46_16\
        );

    \I__3127\ : CascadeMux
    port map (
            O => \N__22998\,
            I => \N__22995\
        );

    \I__3126\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22992\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__22992\,
            I => \N__22989\
        );

    \I__3124\ : Span4Mux_h
    port map (
            O => \N__22989\,
            I => \N__22986\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__22986\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__3122\ : InMux
    port map (
            O => \N__22983\,
            I => \N__22979\
        );

    \I__3121\ : CascadeMux
    port map (
            O => \N__22982\,
            I => \N__22975\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__22979\,
            I => \N__22971\
        );

    \I__3119\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22968\
        );

    \I__3118\ : InMux
    port map (
            O => \N__22975\,
            I => \N__22965\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__22974\,
            I => \N__22962\
        );

    \I__3116\ : Span4Mux_v
    port map (
            O => \N__22971\,
            I => \N__22957\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__22968\,
            I => \N__22957\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__22965\,
            I => \N__22954\
        );

    \I__3113\ : InMux
    port map (
            O => \N__22962\,
            I => \N__22951\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__22957\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__3111\ : Odrv4
    port map (
            O => \N__22954\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__22951\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__3109\ : InMux
    port map (
            O => \N__22944\,
            I => \N__22941\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__22941\,
            I => \N__22938\
        );

    \I__3107\ : Odrv12
    port map (
            O => \N__22938\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__3106\ : CascadeMux
    port map (
            O => \N__22935\,
            I => \N__22929\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__22934\,
            I => \N__22926\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__22933\,
            I => \N__22921\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__22932\,
            I => \N__22918\
        );

    \I__3102\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22910\
        );

    \I__3101\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22910\
        );

    \I__3100\ : InMux
    port map (
            O => \N__22925\,
            I => \N__22910\
        );

    \I__3099\ : InMux
    port map (
            O => \N__22924\,
            I => \N__22901\
        );

    \I__3098\ : InMux
    port map (
            O => \N__22921\,
            I => \N__22901\
        );

    \I__3097\ : InMux
    port map (
            O => \N__22918\,
            I => \N__22901\
        );

    \I__3096\ : InMux
    port map (
            O => \N__22917\,
            I => \N__22901\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__22910\,
            I => \N__22896\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__22901\,
            I => \N__22896\
        );

    \I__3093\ : Span4Mux_h
    port map (
            O => \N__22896\,
            I => \N__22893\
        );

    \I__3092\ : Odrv4
    port map (
            O => \N__22893\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__3091\ : InMux
    port map (
            O => \N__22890\,
            I => \N__22887\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__22887\,
            I => \N__22884\
        );

    \I__3089\ : Odrv4
    port map (
            O => \N__22884\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__22881\,
            I => \N__22878\
        );

    \I__3087\ : InMux
    port map (
            O => \N__22878\,
            I => \N__22875\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__22875\,
            I => \N__22872\
        );

    \I__3085\ : Span4Mux_h
    port map (
            O => \N__22872\,
            I => \N__22869\
        );

    \I__3084\ : Odrv4
    port map (
            O => \N__22869\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__3083\ : InMux
    port map (
            O => \N__22866\,
            I => \N__22863\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__22863\,
            I => \N__22860\
        );

    \I__3081\ : Odrv4
    port map (
            O => \N__22860\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__3080\ : CascadeMux
    port map (
            O => \N__22857\,
            I => \N__22853\
        );

    \I__3079\ : InMux
    port map (
            O => \N__22856\,
            I => \N__22850\
        );

    \I__3078\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22847\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__22850\,
            I => \N__22843\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__22847\,
            I => \N__22839\
        );

    \I__3075\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22836\
        );

    \I__3074\ : Span4Mux_h
    port map (
            O => \N__22843\,
            I => \N__22833\
        );

    \I__3073\ : InMux
    port map (
            O => \N__22842\,
            I => \N__22830\
        );

    \I__3072\ : Span4Mux_h
    port map (
            O => \N__22839\,
            I => \N__22825\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__22836\,
            I => \N__22825\
        );

    \I__3070\ : Odrv4
    port map (
            O => \N__22833\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__22830\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__22825\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__3067\ : InMux
    port map (
            O => \N__22818\,
            I => \N__22815\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__22815\,
            I => \current_shift_inst.PI_CTRL.N_46_21\
        );

    \I__3065\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22809\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__22809\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_2\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__22806\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2_cascade_\
        );

    \I__3062\ : InMux
    port map (
            O => \N__22803\,
            I => \N__22797\
        );

    \I__3061\ : InMux
    port map (
            O => \N__22802\,
            I => \N__22790\
        );

    \I__3060\ : InMux
    port map (
            O => \N__22801\,
            I => \N__22790\
        );

    \I__3059\ : InMux
    port map (
            O => \N__22800\,
            I => \N__22790\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__22797\,
            I => \N__22787\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__22790\,
            I => \N__22784\
        );

    \I__3056\ : Odrv12
    port map (
            O => \N__22787\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__3055\ : Odrv4
    port map (
            O => \N__22784\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__3054\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22776\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__22776\,
            I => \N__22773\
        );

    \I__3052\ : Odrv4
    port map (
            O => \N__22773\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__22770\,
            I => \N__22767\
        );

    \I__3050\ : InMux
    port map (
            O => \N__22767\,
            I => \N__22764\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__22764\,
            I => \N__22761\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__22761\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\
        );

    \I__3047\ : InMux
    port map (
            O => \N__22758\,
            I => \N__22755\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__22755\,
            I => \N__22752\
        );

    \I__3045\ : Odrv12
    port map (
            O => \N__22752\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__3044\ : InMux
    port map (
            O => \N__22749\,
            I => \N__22746\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__22746\,
            I => \N__22743\
        );

    \I__3042\ : Span4Mux_h
    port map (
            O => \N__22743\,
            I => \N__22740\
        );

    \I__3041\ : Odrv4
    port map (
            O => \N__22740\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__3040\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22731\
        );

    \I__3039\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22728\
        );

    \I__3038\ : InMux
    port map (
            O => \N__22735\,
            I => \N__22725\
        );

    \I__3037\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22722\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__22731\,
            I => \N__22719\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__22728\,
            I => \N__22716\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__22725\,
            I => \N__22713\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__22722\,
            I => \N__22710\
        );

    \I__3032\ : Span12Mux_v
    port map (
            O => \N__22719\,
            I => \N__22707\
        );

    \I__3031\ : Odrv12
    port map (
            O => \N__22716\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3030\ : Odrv4
    port map (
            O => \N__22713\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3029\ : Odrv4
    port map (
            O => \N__22710\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3028\ : Odrv12
    port map (
            O => \N__22707\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__3027\ : InMux
    port map (
            O => \N__22698\,
            I => \N__22692\
        );

    \I__3026\ : InMux
    port map (
            O => \N__22697\,
            I => \N__22689\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__22696\,
            I => \N__22686\
        );

    \I__3024\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22683\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__22692\,
            I => \N__22680\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__22689\,
            I => \N__22677\
        );

    \I__3021\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22674\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__22683\,
            I => \N__22671\
        );

    \I__3019\ : Span4Mux_h
    port map (
            O => \N__22680\,
            I => \N__22668\
        );

    \I__3018\ : Span4Mux_v
    port map (
            O => \N__22677\,
            I => \N__22661\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__22674\,
            I => \N__22661\
        );

    \I__3016\ : Span4Mux_h
    port map (
            O => \N__22671\,
            I => \N__22661\
        );

    \I__3015\ : Odrv4
    port map (
            O => \N__22668\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__3014\ : Odrv4
    port map (
            O => \N__22661\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__3013\ : InMux
    port map (
            O => \N__22656\,
            I => \N__22653\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__22653\,
            I => \N__22650\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__22650\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__22647\,
            I => \N__22644\
        );

    \I__3009\ : InMux
    port map (
            O => \N__22644\,
            I => \N__22640\
        );

    \I__3008\ : InMux
    port map (
            O => \N__22643\,
            I => \N__22637\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__22640\,
            I => \N__22632\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__22637\,
            I => \N__22632\
        );

    \I__3005\ : Span4Mux_v
    port map (
            O => \N__22632\,
            I => \N__22627\
        );

    \I__3004\ : InMux
    port map (
            O => \N__22631\,
            I => \N__22622\
        );

    \I__3003\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22622\
        );

    \I__3002\ : Odrv4
    port map (
            O => \N__22627\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__22622\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3000\ : InMux
    port map (
            O => \N__22617\,
            I => \N__22614\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__22614\,
            I => \N__22609\
        );

    \I__2998\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22606\
        );

    \I__2997\ : CascadeMux
    port map (
            O => \N__22612\,
            I => \N__22603\
        );

    \I__2996\ : Span4Mux_v
    port map (
            O => \N__22609\,
            I => \N__22597\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__22606\,
            I => \N__22597\
        );

    \I__2994\ : InMux
    port map (
            O => \N__22603\,
            I => \N__22592\
        );

    \I__2993\ : InMux
    port map (
            O => \N__22602\,
            I => \N__22592\
        );

    \I__2992\ : Odrv4
    port map (
            O => \N__22597\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__22592\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2990\ : CascadeMux
    port map (
            O => \N__22587\,
            I => \current_shift_inst.PI_CTRL.N_46_21_cascade_\
        );

    \I__2989\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22581\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__22581\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\
        );

    \I__2987\ : InMux
    port map (
            O => \N__22578\,
            I => \N__22575\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__22575\,
            I => \N__22572\
        );

    \I__2985\ : Span4Mux_v
    port map (
            O => \N__22572\,
            I => \N__22569\
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__22569\,
            I => \current_shift_inst.PI_CTRL.N_34\
        );

    \I__2983\ : InMux
    port map (
            O => \N__22566\,
            I => \N__22561\
        );

    \I__2982\ : InMux
    port map (
            O => \N__22565\,
            I => \N__22557\
        );

    \I__2981\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22554\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__22561\,
            I => \N__22551\
        );

    \I__2979\ : InMux
    port map (
            O => \N__22560\,
            I => \N__22548\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__22557\,
            I => \N__22543\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__22554\,
            I => \N__22543\
        );

    \I__2976\ : Odrv12
    port map (
            O => \N__22551\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__22548\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2974\ : Odrv12
    port map (
            O => \N__22543\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__22536\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__2972\ : InMux
    port map (
            O => \N__22533\,
            I => \N__22530\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__22530\,
            I => \N__22524\
        );

    \I__2970\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22521\
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__22528\,
            I => \N__22518\
        );

    \I__2968\ : InMux
    port map (
            O => \N__22527\,
            I => \N__22515\
        );

    \I__2967\ : Span4Mux_v
    port map (
            O => \N__22524\,
            I => \N__22510\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__22521\,
            I => \N__22510\
        );

    \I__2965\ : InMux
    port map (
            O => \N__22518\,
            I => \N__22507\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__22515\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2963\ : Odrv4
    port map (
            O => \N__22510\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__22507\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2961\ : InMux
    port map (
            O => \N__22500\,
            I => \N__22497\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__22497\,
            I => \current_shift_inst.PI_CTRL.N_44\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__22494\,
            I => \current_shift_inst.PI_CTRL.N_44_cascade_\
        );

    \I__2958\ : InMux
    port map (
            O => \N__22491\,
            I => \N__22486\
        );

    \I__2957\ : InMux
    port map (
            O => \N__22490\,
            I => \N__22480\
        );

    \I__2956\ : InMux
    port map (
            O => \N__22489\,
            I => \N__22480\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__22486\,
            I => \N__22477\
        );

    \I__2954\ : InMux
    port map (
            O => \N__22485\,
            I => \N__22474\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__22480\,
            I => \N__22471\
        );

    \I__2952\ : Odrv12
    port map (
            O => \N__22477\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__22474\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2950\ : Odrv4
    port map (
            O => \N__22471\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2949\ : CascadeMux
    port map (
            O => \N__22464\,
            I => \N__22461\
        );

    \I__2948\ : InMux
    port map (
            O => \N__22461\,
            I => \N__22458\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__22458\,
            I => \N__22452\
        );

    \I__2946\ : InMux
    port map (
            O => \N__22457\,
            I => \N__22447\
        );

    \I__2945\ : InMux
    port map (
            O => \N__22456\,
            I => \N__22447\
        );

    \I__2944\ : InMux
    port map (
            O => \N__22455\,
            I => \N__22444\
        );

    \I__2943\ : Span4Mux_v
    port map (
            O => \N__22452\,
            I => \N__22439\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__22447\,
            I => \N__22439\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__22444\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__2940\ : Odrv4
    port map (
            O => \N__22439\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__22434\,
            I => \N__22429\
        );

    \I__2938\ : InMux
    port map (
            O => \N__22433\,
            I => \N__22426\
        );

    \I__2937\ : InMux
    port map (
            O => \N__22432\,
            I => \N__22420\
        );

    \I__2936\ : InMux
    port map (
            O => \N__22429\,
            I => \N__22420\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__22426\,
            I => \N__22417\
        );

    \I__2934\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22414\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__22420\,
            I => \N__22411\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__22417\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__22414\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2930\ : Odrv4
    port map (
            O => \N__22411\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2929\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22399\
        );

    \I__2928\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22393\
        );

    \I__2927\ : InMux
    port map (
            O => \N__22402\,
            I => \N__22393\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__22399\,
            I => \N__22390\
        );

    \I__2925\ : InMux
    port map (
            O => \N__22398\,
            I => \N__22387\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__22393\,
            I => \N__22384\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__22390\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__22387\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__22384\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__22377\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__22374\,
            I => \N__22371\
        );

    \I__2918\ : InMux
    port map (
            O => \N__22371\,
            I => \N__22368\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__22368\,
            I => \N__22363\
        );

    \I__2916\ : InMux
    port map (
            O => \N__22367\,
            I => \N__22358\
        );

    \I__2915\ : InMux
    port map (
            O => \N__22366\,
            I => \N__22358\
        );

    \I__2914\ : Span4Mux_v
    port map (
            O => \N__22363\,
            I => \N__22352\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__22358\,
            I => \N__22352\
        );

    \I__2912\ : InMux
    port map (
            O => \N__22357\,
            I => \N__22349\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__22352\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__22349\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__2909\ : InMux
    port map (
            O => \N__22344\,
            I => \N__22341\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__22341\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\
        );

    \I__2907\ : CascadeMux
    port map (
            O => \N__22338\,
            I => \clk_10khz_RNIIENAZ0Z2_cascade_\
        );

    \I__2906\ : InMux
    port map (
            O => \N__22335\,
            I => \N__22332\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__22332\,
            I => \clk_10khz_RNIIENAZ0Z2\
        );

    \I__2904\ : InMux
    port map (
            O => \N__22329\,
            I => \N__22325\
        );

    \I__2903\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22322\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__22325\,
            I => \N__22318\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__22322\,
            I => \N__22315\
        );

    \I__2900\ : InMux
    port map (
            O => \N__22321\,
            I => \N__22309\
        );

    \I__2899\ : Span4Mux_v
    port map (
            O => \N__22318\,
            I => \N__22304\
        );

    \I__2898\ : Span4Mux_v
    port map (
            O => \N__22315\,
            I => \N__22304\
        );

    \I__2897\ : InMux
    port map (
            O => \N__22314\,
            I => \N__22301\
        );

    \I__2896\ : InMux
    port map (
            O => \N__22313\,
            I => \N__22296\
        );

    \I__2895\ : InMux
    port map (
            O => \N__22312\,
            I => \N__22296\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__22309\,
            I => \N__22293\
        );

    \I__2893\ : Odrv4
    port map (
            O => \N__22304\,
            I => un2_counter_8
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__22301\,
            I => un2_counter_8
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__22296\,
            I => un2_counter_8
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__22293\,
            I => un2_counter_8
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__22284\,
            I => \N__22280\
        );

    \I__2888\ : InMux
    port map (
            O => \N__22283\,
            I => \N__22277\
        );

    \I__2887\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22274\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__22277\,
            I => \N__22267\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__22274\,
            I => \N__22264\
        );

    \I__2884\ : InMux
    port map (
            O => \N__22273\,
            I => \N__22261\
        );

    \I__2883\ : InMux
    port map (
            O => \N__22272\,
            I => \N__22258\
        );

    \I__2882\ : InMux
    port map (
            O => \N__22271\,
            I => \N__22253\
        );

    \I__2881\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22253\
        );

    \I__2880\ : Span4Mux_v
    port map (
            O => \N__22267\,
            I => \N__22248\
        );

    \I__2879\ : Span4Mux_v
    port map (
            O => \N__22264\,
            I => \N__22248\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__22261\,
            I => \N__22245\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__22258\,
            I => un2_counter_7
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__22253\,
            I => un2_counter_7
        );

    \I__2875\ : Odrv4
    port map (
            O => \N__22248\,
            I => un2_counter_7
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__22245\,
            I => un2_counter_7
        );

    \I__2873\ : InMux
    port map (
            O => \N__22236\,
            I => \N__22232\
        );

    \I__2872\ : InMux
    port map (
            O => \N__22235\,
            I => \N__22229\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__22232\,
            I => \N__22222\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__22229\,
            I => \N__22219\
        );

    \I__2869\ : InMux
    port map (
            O => \N__22228\,
            I => \N__22216\
        );

    \I__2868\ : InMux
    port map (
            O => \N__22227\,
            I => \N__22213\
        );

    \I__2867\ : InMux
    port map (
            O => \N__22226\,
            I => \N__22208\
        );

    \I__2866\ : InMux
    port map (
            O => \N__22225\,
            I => \N__22208\
        );

    \I__2865\ : Span4Mux_v
    port map (
            O => \N__22222\,
            I => \N__22201\
        );

    \I__2864\ : Span4Mux_v
    port map (
            O => \N__22219\,
            I => \N__22201\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__22216\,
            I => \N__22201\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__22213\,
            I => un2_counter_9
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__22208\,
            I => un2_counter_9
        );

    \I__2860\ : Odrv4
    port map (
            O => \N__22201\,
            I => un2_counter_9
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__22194\,
            I => \N__22188\
        );

    \I__2858\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22183\
        );

    \I__2857\ : InMux
    port map (
            O => \N__22192\,
            I => \N__22183\
        );

    \I__2856\ : InMux
    port map (
            O => \N__22191\,
            I => \N__22178\
        );

    \I__2855\ : InMux
    port map (
            O => \N__22188\,
            I => \N__22178\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__22183\,
            I => clk_10khz_i
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__22178\,
            I => clk_10khz_i
        );

    \I__2852\ : InMux
    port map (
            O => \N__22173\,
            I => \N__22170\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__22170\,
            I => \N__22167\
        );

    \I__2850\ : Odrv4
    port map (
            O => \N__22167\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_1\
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__22164\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__2848\ : CascadeMux
    port map (
            O => \N__22161\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__2847\ : InMux
    port map (
            O => \N__22158\,
            I => \N__22155\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__22155\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__22152\,
            I => \N__22149\
        );

    \I__2844\ : InMux
    port map (
            O => \N__22149\,
            I => \N__22146\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__22146\,
            I => \N__22143\
        );

    \I__2842\ : Span4Mux_h
    port map (
            O => \N__22143\,
            I => \N__22140\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__22140\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__22137\,
            I => \N__22134\
        );

    \I__2839\ : InMux
    port map (
            O => \N__22134\,
            I => \N__22131\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__22131\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__22128\,
            I => \N__22125\
        );

    \I__2836\ : InMux
    port map (
            O => \N__22125\,
            I => \N__22122\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__22122\,
            I => \N__22119\
        );

    \I__2834\ : Span4Mux_h
    port map (
            O => \N__22119\,
            I => \N__22116\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__22116\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__22113\,
            I => \N__22110\
        );

    \I__2831\ : InMux
    port map (
            O => \N__22110\,
            I => \N__22107\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__22107\,
            I => \N__22104\
        );

    \I__2829\ : Odrv4
    port map (
            O => \N__22104\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__22101\,
            I => \N__22098\
        );

    \I__2827\ : InMux
    port map (
            O => \N__22098\,
            I => \N__22095\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__22095\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__2825\ : CascadeMux
    port map (
            O => \N__22092\,
            I => \N__22089\
        );

    \I__2824\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22086\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__22086\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__2822\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22080\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__22080\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__22077\,
            I => \N__22074\
        );

    \I__2819\ : InMux
    port map (
            O => \N__22074\,
            I => \N__22068\
        );

    \I__2818\ : InMux
    port map (
            O => \N__22073\,
            I => \N__22065\
        );

    \I__2817\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22062\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__22071\,
            I => \N__22059\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__22068\,
            I => \N__22054\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__22065\,
            I => \N__22054\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__22062\,
            I => \N__22051\
        );

    \I__2812\ : InMux
    port map (
            O => \N__22059\,
            I => \N__22048\
        );

    \I__2811\ : Span4Mux_h
    port map (
            O => \N__22054\,
            I => \N__22045\
        );

    \I__2810\ : Odrv4
    port map (
            O => \N__22051\,
            I => \counterZ0Z_0\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__22048\,
            I => \counterZ0Z_0\
        );

    \I__2808\ : Odrv4
    port map (
            O => \N__22045\,
            I => \counterZ0Z_0\
        );

    \I__2807\ : InMux
    port map (
            O => \N__22038\,
            I => \N__22035\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__22035\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__22032\,
            I => \N__22029\
        );

    \I__2804\ : InMux
    port map (
            O => \N__22029\,
            I => \N__22026\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__22026\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__22023\,
            I => \N__22020\
        );

    \I__2801\ : InMux
    port map (
            O => \N__22020\,
            I => \N__22017\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__22017\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__2799\ : InMux
    port map (
            O => \N__22014\,
            I => \N__22011\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__22011\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__22008\,
            I => \N__22005\
        );

    \I__2796\ : InMux
    port map (
            O => \N__22005\,
            I => \N__22002\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__22002\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__2794\ : InMux
    port map (
            O => \N__21999\,
            I => \N__21996\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__21996\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__21993\,
            I => \N__21990\
        );

    \I__2791\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21987\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__21987\,
            I => \N__21984\
        );

    \I__2789\ : Odrv4
    port map (
            O => \N__21984\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__21981\,
            I => \N__21978\
        );

    \I__2787\ : InMux
    port map (
            O => \N__21978\,
            I => \N__21975\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__21975\,
            I => \N__21972\
        );

    \I__2785\ : Odrv4
    port map (
            O => \N__21972\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__2784\ : InMux
    port map (
            O => \N__21969\,
            I => \N__21966\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__21966\,
            I => \N__21963\
        );

    \I__2782\ : Odrv12
    port map (
            O => \N__21963\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__21960\,
            I => \N__21957\
        );

    \I__2780\ : InMux
    port map (
            O => \N__21957\,
            I => \N__21954\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__21954\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__2778\ : InMux
    port map (
            O => \N__21951\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\
        );

    \I__2777\ : InMux
    port map (
            O => \N__21948\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__2776\ : InMux
    port map (
            O => \N__21945\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__2775\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21939\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__21939\,
            I => \N__21936\
        );

    \I__2773\ : Odrv4
    port map (
            O => \N__21936\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__2772\ : InMux
    port map (
            O => \N__21933\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__2771\ : InMux
    port map (
            O => \N__21930\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__2770\ : InMux
    port map (
            O => \N__21927\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__2769\ : InMux
    port map (
            O => \N__21924\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__21921\,
            I => \N__21918\
        );

    \I__2767\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21915\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__21915\,
            I => \N__21912\
        );

    \I__2765\ : Odrv12
    port map (
            O => \N__21912\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__21909\,
            I => \N__21906\
        );

    \I__2763\ : InMux
    port map (
            O => \N__21906\,
            I => \N__21903\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__21903\,
            I => \N__21900\
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__21900\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__2760\ : InMux
    port map (
            O => \N__21897\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\
        );

    \I__2759\ : InMux
    port map (
            O => \N__21894\,
            I => \N__21891\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__21891\,
            I => \N__21888\
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__21888\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__2756\ : InMux
    port map (
            O => \N__21885\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__2755\ : InMux
    port map (
            O => \N__21882\,
            I => \N__21879\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__21879\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__2753\ : InMux
    port map (
            O => \N__21876\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__21873\,
            I => \N__21870\
        );

    \I__2751\ : InMux
    port map (
            O => \N__21870\,
            I => \N__21867\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__21867\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__2749\ : InMux
    port map (
            O => \N__21864\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__2748\ : InMux
    port map (
            O => \N__21861\,
            I => \N__21858\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__21858\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__2746\ : InMux
    port map (
            O => \N__21855\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__21852\,
            I => \N__21849\
        );

    \I__2744\ : InMux
    port map (
            O => \N__21849\,
            I => \N__21846\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__21846\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__2742\ : InMux
    port map (
            O => \N__21843\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__2741\ : InMux
    port map (
            O => \N__21840\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__2740\ : InMux
    port map (
            O => \N__21837\,
            I => \bfn_5_13_0_\
        );

    \I__2739\ : InMux
    port map (
            O => \N__21834\,
            I => \N__21831\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__21831\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__2737\ : InMux
    port map (
            O => \N__21828\,
            I => \bfn_5_11_0_\
        );

    \I__2736\ : CascadeMux
    port map (
            O => \N__21825\,
            I => \N__21822\
        );

    \I__2735\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21819\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__21819\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__2733\ : InMux
    port map (
            O => \N__21816\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\
        );

    \I__2732\ : InMux
    port map (
            O => \N__21813\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__2731\ : InMux
    port map (
            O => \N__21810\,
            I => \N__21807\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__21807\,
            I => \N__21804\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__21804\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__2728\ : InMux
    port map (
            O => \N__21801\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__2727\ : InMux
    port map (
            O => \N__21798\,
            I => \N__21795\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__21795\,
            I => \N__21792\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__21792\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__2724\ : InMux
    port map (
            O => \N__21789\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__21786\,
            I => \N__21783\
        );

    \I__2722\ : InMux
    port map (
            O => \N__21783\,
            I => \N__21780\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__21780\,
            I => \N__21777\
        );

    \I__2720\ : Odrv4
    port map (
            O => \N__21777\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__2719\ : InMux
    port map (
            O => \N__21774\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__2718\ : InMux
    port map (
            O => \N__21771\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__2717\ : InMux
    port map (
            O => \N__21768\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__2716\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21762\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__21762\,
            I => \N__21759\
        );

    \I__2714\ : Odrv4
    port map (
            O => \N__21759\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__2713\ : InMux
    port map (
            O => \N__21756\,
            I => \bfn_5_12_0_\
        );

    \I__2712\ : InMux
    port map (
            O => \N__21753\,
            I => \N__21750\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__21750\,
            I => \N__21747\
        );

    \I__2710\ : Span4Mux_v
    port map (
            O => \N__21747\,
            I => \N__21742\
        );

    \I__2709\ : InMux
    port map (
            O => \N__21746\,
            I => \N__21739\
        );

    \I__2708\ : InMux
    port map (
            O => \N__21745\,
            I => \N__21736\
        );

    \I__2707\ : Odrv4
    port map (
            O => \N__21742\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__21739\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__21736\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__2704\ : InMux
    port map (
            O => \N__21729\,
            I => \N__21726\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__21726\,
            I => \N__21723\
        );

    \I__2702\ : Span4Mux_v
    port map (
            O => \N__21723\,
            I => \N__21718\
        );

    \I__2701\ : InMux
    port map (
            O => \N__21722\,
            I => \N__21715\
        );

    \I__2700\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21712\
        );

    \I__2699\ : Odrv4
    port map (
            O => \N__21718\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__21715\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__21712\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2696\ : InMux
    port map (
            O => \N__21705\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__21702\,
            I => \N__21699\
        );

    \I__2694\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21694\
        );

    \I__2693\ : InMux
    port map (
            O => \N__21698\,
            I => \N__21691\
        );

    \I__2692\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21688\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__21694\,
            I => \N__21683\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__21691\,
            I => \N__21683\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__21688\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2688\ : Odrv4
    port map (
            O => \N__21683\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2687\ : InMux
    port map (
            O => \N__21678\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__2686\ : InMux
    port map (
            O => \N__21675\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__2685\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21669\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__21669\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__2683\ : InMux
    port map (
            O => \N__21666\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__2682\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21660\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__21660\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__2680\ : InMux
    port map (
            O => \N__21657\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__2679\ : InMux
    port map (
            O => \N__21654\,
            I => \N__21651\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__21651\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__2677\ : InMux
    port map (
            O => \N__21648\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__2676\ : InMux
    port map (
            O => \N__21645\,
            I => \N__21642\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__21642\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__2674\ : InMux
    port map (
            O => \N__21639\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__2673\ : InMux
    port map (
            O => \N__21636\,
            I => \N__21633\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__21633\,
            I => \N__21630\
        );

    \I__2671\ : Odrv4
    port map (
            O => \N__21630\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_8\
        );

    \I__2670\ : InMux
    port map (
            O => \N__21627\,
            I => \N__21624\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__21624\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_3\
        );

    \I__2668\ : InMux
    port map (
            O => \N__21621\,
            I => \N__21618\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__21618\,
            I => \N__21615\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__21615\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_7\
        );

    \I__2665\ : InMux
    port map (
            O => \N__21612\,
            I => \N__21609\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__21609\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_5\
        );

    \I__2663\ : InMux
    port map (
            O => \N__21606\,
            I => \N__21603\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__21603\,
            I => \N__21600\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__21600\,
            I => \N__21597\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__21597\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__2659\ : InMux
    port map (
            O => \N__21594\,
            I => \N__21590\
        );

    \I__2658\ : InMux
    port map (
            O => \N__21593\,
            I => \N__21587\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__21590\,
            I => \counterZ0Z_2\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__21587\,
            I => \counterZ0Z_2\
        );

    \I__2655\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21577\
        );

    \I__2654\ : InMux
    port map (
            O => \N__21581\,
            I => \N__21574\
        );

    \I__2653\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21571\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__21577\,
            I => \counterZ0Z_1\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__21574\,
            I => \counterZ0Z_1\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__21571\,
            I => \counterZ0Z_1\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__21564\,
            I => \un2_counter_5_cascade_\
        );

    \I__2648\ : InMux
    port map (
            O => \N__21561\,
            I => \N__21557\
        );

    \I__2647\ : InMux
    port map (
            O => \N__21560\,
            I => \N__21554\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__21557\,
            I => \counterZ0Z_8\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__21554\,
            I => \counterZ0Z_8\
        );

    \I__2644\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21545\
        );

    \I__2643\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21542\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__21545\,
            I => \counterZ0Z_11\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__21542\,
            I => \counterZ0Z_11\
        );

    \I__2640\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21533\
        );

    \I__2639\ : InMux
    port map (
            O => \N__21536\,
            I => \N__21530\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__21533\,
            I => \counterZ0Z_9\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__21530\,
            I => \counterZ0Z_9\
        );

    \I__2636\ : InMux
    port map (
            O => \N__21525\,
            I => \N__21521\
        );

    \I__2635\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21518\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__21521\,
            I => \counterZ0Z_5\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__21518\,
            I => \counterZ0Z_5\
        );

    \I__2632\ : InMux
    port map (
            O => \N__21513\,
            I => \N__21509\
        );

    \I__2631\ : InMux
    port map (
            O => \N__21512\,
            I => \N__21506\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__21509\,
            I => \counterZ0Z_4\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__21506\,
            I => \counterZ0Z_4\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__21501\,
            I => \N__21497\
        );

    \I__2627\ : InMux
    port map (
            O => \N__21500\,
            I => \N__21494\
        );

    \I__2626\ : InMux
    port map (
            O => \N__21497\,
            I => \N__21491\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__21494\,
            I => \counterZ0Z_6\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__21491\,
            I => \counterZ0Z_6\
        );

    \I__2623\ : InMux
    port map (
            O => \N__21486\,
            I => \N__21482\
        );

    \I__2622\ : InMux
    port map (
            O => \N__21485\,
            I => \N__21479\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__21482\,
            I => \counterZ0Z_3\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__21479\,
            I => \counterZ0Z_3\
        );

    \I__2619\ : InMux
    port map (
            O => \N__21474\,
            I => \N__21471\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__21471\,
            I => \N__21468\
        );

    \I__2617\ : Span4Mux_h
    port map (
            O => \N__21468\,
            I => \N__21465\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__21465\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_4\
        );

    \I__2615\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21459\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__21459\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_2\
        );

    \I__2613\ : InMux
    port map (
            O => \N__21456\,
            I => \N__21453\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__21453\,
            I => \N__21450\
        );

    \I__2611\ : Span4Mux_v
    port map (
            O => \N__21450\,
            I => \N__21447\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__21447\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_6\
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__21444\,
            I => \N__21441\
        );

    \I__2608\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21438\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__21438\,
            I => \counter_RNO_0Z0Z_12\
        );

    \I__2606\ : CascadeMux
    port map (
            O => \N__21435\,
            I => \N__21431\
        );

    \I__2605\ : InMux
    port map (
            O => \N__21434\,
            I => \N__21428\
        );

    \I__2604\ : InMux
    port map (
            O => \N__21431\,
            I => \N__21425\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__21428\,
            I => \counterZ0Z_12\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__21425\,
            I => \counterZ0Z_12\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__21420\,
            I => \N__21417\
        );

    \I__2600\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21414\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__21414\,
            I => \counter_RNO_0Z0Z_10\
        );

    \I__2598\ : InMux
    port map (
            O => \N__21411\,
            I => \N__21407\
        );

    \I__2597\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21404\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__21407\,
            I => \counterZ0Z_10\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__21404\,
            I => \counterZ0Z_10\
        );

    \I__2594\ : InMux
    port map (
            O => \N__21399\,
            I => \N__21393\
        );

    \I__2593\ : InMux
    port map (
            O => \N__21398\,
            I => \N__21393\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__21393\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2591\ : InMux
    port map (
            O => \N__21390\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2590\ : InMux
    port map (
            O => \N__21387\,
            I => \N__21383\
        );

    \I__2589\ : InMux
    port map (
            O => \N__21386\,
            I => \N__21380\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__21383\,
            I => \N__21375\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__21380\,
            I => \N__21375\
        );

    \I__2586\ : Span4Mux_v
    port map (
            O => \N__21375\,
            I => \N__21372\
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__21372\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2584\ : InMux
    port map (
            O => \N__21369\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2583\ : InMux
    port map (
            O => \N__21366\,
            I => \N__21360\
        );

    \I__2582\ : InMux
    port map (
            O => \N__21365\,
            I => \N__21360\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__21360\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2580\ : InMux
    port map (
            O => \N__21357\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2579\ : InMux
    port map (
            O => \N__21354\,
            I => \N__21351\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__21351\,
            I => \N__21347\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__21350\,
            I => \N__21344\
        );

    \I__2576\ : Span4Mux_h
    port map (
            O => \N__21347\,
            I => \N__21341\
        );

    \I__2575\ : InMux
    port map (
            O => \N__21344\,
            I => \N__21338\
        );

    \I__2574\ : Odrv4
    port map (
            O => \N__21341\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__21338\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2572\ : InMux
    port map (
            O => \N__21333\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2571\ : CascadeMux
    port map (
            O => \N__21330\,
            I => \N__21327\
        );

    \I__2570\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21324\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__21324\,
            I => \N__21320\
        );

    \I__2568\ : InMux
    port map (
            O => \N__21323\,
            I => \N__21317\
        );

    \I__2567\ : Span4Mux_h
    port map (
            O => \N__21320\,
            I => \N__21314\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__21317\,
            I => \N__21311\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__21314\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2564\ : Odrv4
    port map (
            O => \N__21311\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2563\ : InMux
    port map (
            O => \N__21306\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2562\ : InMux
    port map (
            O => \N__21303\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2561\ : InMux
    port map (
            O => \N__21300\,
            I => \N__21297\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__21297\,
            I => \N__21288\
        );

    \I__2559\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21285\
        );

    \I__2558\ : InMux
    port map (
            O => \N__21295\,
            I => \N__21281\
        );

    \I__2557\ : InMux
    port map (
            O => \N__21294\,
            I => \N__21272\
        );

    \I__2556\ : InMux
    port map (
            O => \N__21293\,
            I => \N__21272\
        );

    \I__2555\ : InMux
    port map (
            O => \N__21292\,
            I => \N__21272\
        );

    \I__2554\ : InMux
    port map (
            O => \N__21291\,
            I => \N__21272\
        );

    \I__2553\ : Span4Mux_v
    port map (
            O => \N__21288\,
            I => \N__21267\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__21285\,
            I => \N__21267\
        );

    \I__2551\ : CascadeMux
    port map (
            O => \N__21284\,
            I => \N__21262\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__21281\,
            I => \N__21259\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__21272\,
            I => \N__21254\
        );

    \I__2548\ : Span4Mux_h
    port map (
            O => \N__21267\,
            I => \N__21254\
        );

    \I__2547\ : InMux
    port map (
            O => \N__21266\,
            I => \N__21251\
        );

    \I__2546\ : InMux
    port map (
            O => \N__21265\,
            I => \N__21246\
        );

    \I__2545\ : InMux
    port map (
            O => \N__21262\,
            I => \N__21246\
        );

    \I__2544\ : Span4Mux_v
    port map (
            O => \N__21259\,
            I => \N__21239\
        );

    \I__2543\ : Span4Mux_v
    port map (
            O => \N__21254\,
            I => \N__21239\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__21251\,
            I => \N__21239\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__21246\,
            I => \N__21234\
        );

    \I__2540\ : Span4Mux_h
    port map (
            O => \N__21239\,
            I => \N__21234\
        );

    \I__2539\ : Span4Mux_v
    port map (
            O => \N__21234\,
            I => \N__21231\
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__21231\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__21228\,
            I => \N__21225\
        );

    \I__2536\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21222\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__21222\,
            I => \counter_RNO_0Z0Z_7\
        );

    \I__2534\ : InMux
    port map (
            O => \N__21219\,
            I => \N__21215\
        );

    \I__2533\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21212\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__21215\,
            I => \counterZ0Z_7\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__21212\,
            I => \counterZ0Z_7\
        );

    \I__2530\ : InMux
    port map (
            O => \N__21207\,
            I => \N__21201\
        );

    \I__2529\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21201\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__21201\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2527\ : InMux
    port map (
            O => \N__21198\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\
        );

    \I__2526\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21189\
        );

    \I__2525\ : InMux
    port map (
            O => \N__21194\,
            I => \N__21189\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__21189\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2523\ : InMux
    port map (
            O => \N__21186\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2522\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21177\
        );

    \I__2521\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21177\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__21177\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2519\ : InMux
    port map (
            O => \N__21174\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2518\ : InMux
    port map (
            O => \N__21171\,
            I => \N__21165\
        );

    \I__2517\ : InMux
    port map (
            O => \N__21170\,
            I => \N__21165\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__21165\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2515\ : InMux
    port map (
            O => \N__21162\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__21159\,
            I => \N__21156\
        );

    \I__2513\ : InMux
    port map (
            O => \N__21156\,
            I => \N__21150\
        );

    \I__2512\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21150\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__21150\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2510\ : InMux
    port map (
            O => \N__21147\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2509\ : InMux
    port map (
            O => \N__21144\,
            I => \N__21141\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__21141\,
            I => \N__21137\
        );

    \I__2507\ : InMux
    port map (
            O => \N__21140\,
            I => \N__21134\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__21137\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__21134\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2504\ : InMux
    port map (
            O => \N__21129\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2503\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21122\
        );

    \I__2502\ : CascadeMux
    port map (
            O => \N__21125\,
            I => \N__21119\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__21122\,
            I => \N__21116\
        );

    \I__2500\ : InMux
    port map (
            O => \N__21119\,
            I => \N__21113\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__21116\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__21113\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2497\ : InMux
    port map (
            O => \N__21108\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2496\ : CascadeMux
    port map (
            O => \N__21105\,
            I => \N__21102\
        );

    \I__2495\ : InMux
    port map (
            O => \N__21102\,
            I => \N__21098\
        );

    \I__2494\ : InMux
    port map (
            O => \N__21101\,
            I => \N__21095\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__21098\,
            I => \N__21090\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__21095\,
            I => \N__21090\
        );

    \I__2491\ : Span4Mux_v
    port map (
            O => \N__21090\,
            I => \N__21087\
        );

    \I__2490\ : Odrv4
    port map (
            O => \N__21087\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2489\ : InMux
    port map (
            O => \N__21084\,
            I => \bfn_4_16_0_\
        );

    \I__2488\ : InMux
    port map (
            O => \N__21081\,
            I => \N__21077\
        );

    \I__2487\ : InMux
    port map (
            O => \N__21080\,
            I => \N__21074\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__21077\,
            I => \N__21071\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__21074\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__21071\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2483\ : InMux
    port map (
            O => \N__21066\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__21063\,
            I => \N__21060\
        );

    \I__2481\ : InMux
    port map (
            O => \N__21060\,
            I => \N__21056\
        );

    \I__2480\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21052\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__21056\,
            I => \N__21049\
        );

    \I__2478\ : InMux
    port map (
            O => \N__21055\,
            I => \N__21046\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__21052\,
            I => \N__21043\
        );

    \I__2476\ : Span4Mux_v
    port map (
            O => \N__21049\,
            I => \N__21036\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__21046\,
            I => \N__21036\
        );

    \I__2474\ : Span4Mux_v
    port map (
            O => \N__21043\,
            I => \N__21036\
        );

    \I__2473\ : Odrv4
    port map (
            O => \N__21036\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2472\ : InMux
    port map (
            O => \N__21033\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\
        );

    \I__2471\ : InMux
    port map (
            O => \N__21030\,
            I => \N__21027\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__21027\,
            I => \N__21024\
        );

    \I__2469\ : Span4Mux_h
    port map (
            O => \N__21024\,
            I => \N__21020\
        );

    \I__2468\ : InMux
    port map (
            O => \N__21023\,
            I => \N__21017\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__21020\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__21017\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2465\ : InMux
    port map (
            O => \N__21012\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__21009\,
            I => \N__21006\
        );

    \I__2463\ : InMux
    port map (
            O => \N__21006\,
            I => \N__21000\
        );

    \I__2462\ : InMux
    port map (
            O => \N__21005\,
            I => \N__21000\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__21000\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2460\ : InMux
    port map (
            O => \N__20997\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2459\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20988\
        );

    \I__2458\ : InMux
    port map (
            O => \N__20993\,
            I => \N__20988\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__20988\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2456\ : InMux
    port map (
            O => \N__20985\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__20982\,
            I => \N__20978\
        );

    \I__2454\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20975\
        );

    \I__2453\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20972\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__20975\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__20972\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2450\ : InMux
    port map (
            O => \N__20967\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2449\ : InMux
    port map (
            O => \N__20964\,
            I => \N__20961\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__20961\,
            I => \N__20957\
        );

    \I__2447\ : InMux
    port map (
            O => \N__20960\,
            I => \N__20954\
        );

    \I__2446\ : Odrv4
    port map (
            O => \N__20957\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__20954\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2444\ : InMux
    port map (
            O => \N__20949\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2443\ : InMux
    port map (
            O => \N__20946\,
            I => \N__20943\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__20943\,
            I => \N__20940\
        );

    \I__2441\ : Span4Mux_h
    port map (
            O => \N__20940\,
            I => \N__20936\
        );

    \I__2440\ : InMux
    port map (
            O => \N__20939\,
            I => \N__20933\
        );

    \I__2439\ : Odrv4
    port map (
            O => \N__20936\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__20933\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2437\ : InMux
    port map (
            O => \N__20928\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2436\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20921\
        );

    \I__2435\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20918\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__20921\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__20918\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2432\ : InMux
    port map (
            O => \N__20913\,
            I => \bfn_4_15_0_\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__20910\,
            I => \N__20907\
        );

    \I__2430\ : InMux
    port map (
            O => \N__20907\,
            I => \N__20904\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__20904\,
            I => \N__20901\
        );

    \I__2428\ : Odrv12
    port map (
            O => \N__20901\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__20898\,
            I => \N__20895\
        );

    \I__2426\ : InMux
    port map (
            O => \N__20895\,
            I => \N__20892\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__20892\,
            I => \N__20889\
        );

    \I__2424\ : Span4Mux_v
    port map (
            O => \N__20889\,
            I => \N__20886\
        );

    \I__2423\ : Span4Mux_h
    port map (
            O => \N__20886\,
            I => \N__20883\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__20883\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2421\ : InMux
    port map (
            O => \N__20880\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\
        );

    \I__2420\ : InMux
    port map (
            O => \N__20877\,
            I => \N__20874\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__20874\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__20871\,
            I => \N__20868\
        );

    \I__2417\ : InMux
    port map (
            O => \N__20868\,
            I => \N__20865\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__20865\,
            I => \N__20862\
        );

    \I__2415\ : Span4Mux_h
    port map (
            O => \N__20862\,
            I => \N__20859\
        );

    \I__2414\ : Span4Mux_v
    port map (
            O => \N__20859\,
            I => \N__20856\
        );

    \I__2413\ : Odrv4
    port map (
            O => \N__20856\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2412\ : InMux
    port map (
            O => \N__20853\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__20850\,
            I => \N__20847\
        );

    \I__2410\ : InMux
    port map (
            O => \N__20847\,
            I => \N__20843\
        );

    \I__2409\ : CascadeMux
    port map (
            O => \N__20846\,
            I => \N__20840\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__20843\,
            I => \N__20837\
        );

    \I__2407\ : InMux
    port map (
            O => \N__20840\,
            I => \N__20833\
        );

    \I__2406\ : Span4Mux_h
    port map (
            O => \N__20837\,
            I => \N__20830\
        );

    \I__2405\ : InMux
    port map (
            O => \N__20836\,
            I => \N__20827\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__20833\,
            I => \N__20820\
        );

    \I__2403\ : Span4Mux_v
    port map (
            O => \N__20830\,
            I => \N__20820\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__20827\,
            I => \N__20820\
        );

    \I__2401\ : Span4Mux_h
    port map (
            O => \N__20820\,
            I => \N__20817\
        );

    \I__2400\ : Odrv4
    port map (
            O => \N__20817\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2399\ : InMux
    port map (
            O => \N__20814\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__20811\,
            I => \N__20806\
        );

    \I__2397\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20800\
        );

    \I__2396\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20800\
        );

    \I__2395\ : InMux
    port map (
            O => \N__20806\,
            I => \N__20797\
        );

    \I__2394\ : InMux
    port map (
            O => \N__20805\,
            I => \N__20794\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__20800\,
            I => \N__20791\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__20797\,
            I => \N__20788\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__20794\,
            I => \N__20785\
        );

    \I__2390\ : Span4Mux_h
    port map (
            O => \N__20791\,
            I => \N__20782\
        );

    \I__2389\ : Odrv4
    port map (
            O => \N__20788\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__20785\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2387\ : Odrv4
    port map (
            O => \N__20782\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2386\ : InMux
    port map (
            O => \N__20775\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2385\ : InMux
    port map (
            O => \N__20772\,
            I => \N__20769\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__20769\,
            I => \N__20766\
        );

    \I__2383\ : Odrv12
    port map (
            O => \N__20766\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__20763\,
            I => \N__20760\
        );

    \I__2381\ : InMux
    port map (
            O => \N__20760\,
            I => \N__20757\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__20757\,
            I => \N__20753\
        );

    \I__2379\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20750\
        );

    \I__2378\ : Span4Mux_v
    port map (
            O => \N__20753\,
            I => \N__20744\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__20750\,
            I => \N__20744\
        );

    \I__2376\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20741\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__20744\,
            I => \N__20736\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__20741\,
            I => \N__20736\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__20736\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2372\ : InMux
    port map (
            O => \N__20733\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2371\ : CascadeMux
    port map (
            O => \N__20730\,
            I => \N__20727\
        );

    \I__2370\ : InMux
    port map (
            O => \N__20727\,
            I => \N__20724\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__20724\,
            I => \N__20719\
        );

    \I__2368\ : InMux
    port map (
            O => \N__20723\,
            I => \N__20716\
        );

    \I__2367\ : InMux
    port map (
            O => \N__20722\,
            I => \N__20713\
        );

    \I__2366\ : Span4Mux_v
    port map (
            O => \N__20719\,
            I => \N__20708\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__20716\,
            I => \N__20708\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__20713\,
            I => \N__20705\
        );

    \I__2363\ : Span4Mux_h
    port map (
            O => \N__20708\,
            I => \N__20702\
        );

    \I__2362\ : Odrv4
    port map (
            O => \N__20705\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2361\ : Odrv4
    port map (
            O => \N__20702\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2360\ : InMux
    port map (
            O => \N__20697\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__20694\,
            I => \N__20691\
        );

    \I__2358\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20688\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__20688\,
            I => \N__20685\
        );

    \I__2356\ : Span4Mux_v
    port map (
            O => \N__20685\,
            I => \N__20682\
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__20682\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__20679\,
            I => \N__20676\
        );

    \I__2353\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20671\
        );

    \I__2352\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20668\
        );

    \I__2351\ : InMux
    port map (
            O => \N__20674\,
            I => \N__20665\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__20671\,
            I => \N__20662\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__20668\,
            I => \N__20659\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__20665\,
            I => \N__20656\
        );

    \I__2347\ : Span4Mux_v
    port map (
            O => \N__20662\,
            I => \N__20653\
        );

    \I__2346\ : Span4Mux_v
    port map (
            O => \N__20659\,
            I => \N__20648\
        );

    \I__2345\ : Span4Mux_s3_h
    port map (
            O => \N__20656\,
            I => \N__20648\
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__20653\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__20648\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2342\ : InMux
    port map (
            O => \N__20643\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__20640\,
            I => \N__20637\
        );

    \I__2340\ : InMux
    port map (
            O => \N__20637\,
            I => \N__20634\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__20634\,
            I => \N__20630\
        );

    \I__2338\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20627\
        );

    \I__2337\ : Span4Mux_v
    port map (
            O => \N__20630\,
            I => \N__20623\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__20627\,
            I => \N__20620\
        );

    \I__2335\ : InMux
    port map (
            O => \N__20626\,
            I => \N__20617\
        );

    \I__2334\ : Span4Mux_s2_h
    port map (
            O => \N__20623\,
            I => \N__20610\
        );

    \I__2333\ : Span4Mux_v
    port map (
            O => \N__20620\,
            I => \N__20610\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__20617\,
            I => \N__20610\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__20610\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2330\ : InMux
    port map (
            O => \N__20607\,
            I => \bfn_4_14_0_\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__20604\,
            I => \N__20601\
        );

    \I__2328\ : InMux
    port map (
            O => \N__20601\,
            I => \N__20598\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__20598\,
            I => \N__20595\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__20595\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__20592\,
            I => \N__20589\
        );

    \I__2324\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20586\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__20586\,
            I => \N__20583\
        );

    \I__2322\ : Span4Mux_v
    port map (
            O => \N__20583\,
            I => \N__20580\
        );

    \I__2321\ : Span4Mux_h
    port map (
            O => \N__20580\,
            I => \N__20577\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__20577\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__20574\,
            I => \N__20571\
        );

    \I__2318\ : InMux
    port map (
            O => \N__20571\,
            I => \N__20568\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__20568\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\
        );

    \I__2316\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20558\
        );

    \I__2315\ : InMux
    port map (
            O => \N__20564\,
            I => \N__20558\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__20563\,
            I => \N__20555\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__20558\,
            I => \N__20545\
        );

    \I__2312\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20542\
        );

    \I__2311\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20535\
        );

    \I__2310\ : InMux
    port map (
            O => \N__20553\,
            I => \N__20535\
        );

    \I__2309\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20535\
        );

    \I__2308\ : InMux
    port map (
            O => \N__20551\,
            I => \N__20526\
        );

    \I__2307\ : InMux
    port map (
            O => \N__20550\,
            I => \N__20526\
        );

    \I__2306\ : InMux
    port map (
            O => \N__20549\,
            I => \N__20526\
        );

    \I__2305\ : InMux
    port map (
            O => \N__20548\,
            I => \N__20526\
        );

    \I__2304\ : Span4Mux_v
    port map (
            O => \N__20545\,
            I => \N__20517\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__20542\,
            I => \N__20517\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__20535\,
            I => \N__20517\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__20526\,
            I => \N__20517\
        );

    \I__2300\ : Span4Mux_h
    port map (
            O => \N__20517\,
            I => \N__20514\
        );

    \I__2299\ : Span4Mux_v
    port map (
            O => \N__20514\,
            I => \N__20510\
        );

    \I__2298\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20507\
        );

    \I__2297\ : Odrv4
    port map (
            O => \N__20510\,
            I => pwm_duty_input_6
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__20507\,
            I => pwm_duty_input_6
        );

    \I__2295\ : InMux
    port map (
            O => \N__20502\,
            I => \N__20493\
        );

    \I__2294\ : InMux
    port map (
            O => \N__20501\,
            I => \N__20493\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__20500\,
            I => \N__20486\
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__20499\,
            I => \N__20483\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__20498\,
            I => \N__20479\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__20493\,
            I => \N__20476\
        );

    \I__2289\ : InMux
    port map (
            O => \N__20492\,
            I => \N__20467\
        );

    \I__2288\ : InMux
    port map (
            O => \N__20491\,
            I => \N__20467\
        );

    \I__2287\ : InMux
    port map (
            O => \N__20490\,
            I => \N__20467\
        );

    \I__2286\ : InMux
    port map (
            O => \N__20489\,
            I => \N__20467\
        );

    \I__2285\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20458\
        );

    \I__2284\ : InMux
    port map (
            O => \N__20483\,
            I => \N__20458\
        );

    \I__2283\ : InMux
    port map (
            O => \N__20482\,
            I => \N__20458\
        );

    \I__2282\ : InMux
    port map (
            O => \N__20479\,
            I => \N__20458\
        );

    \I__2281\ : Span4Mux_v
    port map (
            O => \N__20476\,
            I => \N__20451\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__20467\,
            I => \N__20451\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__20458\,
            I => \N__20451\
        );

    \I__2278\ : Odrv4
    port map (
            O => \N__20451\,
            I => i8_mux
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__20448\,
            I => \N__20441\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__20447\,
            I => \N__20437\
        );

    \I__2275\ : CascadeMux
    port map (
            O => \N__20446\,
            I => \N__20431\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__20445\,
            I => \N__20428\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__20444\,
            I => \N__20425\
        );

    \I__2272\ : InMux
    port map (
            O => \N__20441\,
            I => \N__20419\
        );

    \I__2271\ : InMux
    port map (
            O => \N__20440\,
            I => \N__20419\
        );

    \I__2270\ : InMux
    port map (
            O => \N__20437\,
            I => \N__20416\
        );

    \I__2269\ : InMux
    port map (
            O => \N__20436\,
            I => \N__20409\
        );

    \I__2268\ : InMux
    port map (
            O => \N__20435\,
            I => \N__20409\
        );

    \I__2267\ : InMux
    port map (
            O => \N__20434\,
            I => \N__20409\
        );

    \I__2266\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20400\
        );

    \I__2265\ : InMux
    port map (
            O => \N__20428\,
            I => \N__20400\
        );

    \I__2264\ : InMux
    port map (
            O => \N__20425\,
            I => \N__20400\
        );

    \I__2263\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20400\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__20419\,
            I => \N__20397\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__20416\,
            I => \N__20390\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__20409\,
            I => \N__20390\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__20400\,
            I => \N__20390\
        );

    \I__2258\ : Span4Mux_h
    port map (
            O => \N__20397\,
            I => \N__20387\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__20390\,
            I => \N_28_mux\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__20387\,
            I => \N_28_mux\
        );

    \I__2255\ : InMux
    port map (
            O => \N__20382\,
            I => \N__20379\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__20379\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\
        );

    \I__2253\ : InMux
    port map (
            O => \N__20376\,
            I => \N__20373\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__20373\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_9\
        );

    \I__2251\ : InMux
    port map (
            O => \N__20370\,
            I => \bfn_4_6_0_\
        );

    \I__2250\ : InMux
    port map (
            O => \N__20367\,
            I => un5_counter_cry_9
        );

    \I__2249\ : InMux
    port map (
            O => \N__20364\,
            I => un5_counter_cry_10
        );

    \I__2248\ : InMux
    port map (
            O => \N__20361\,
            I => un5_counter_cry_11
        );

    \I__2247\ : InMux
    port map (
            O => \N__20358\,
            I => \N__20355\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__20355\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\
        );

    \I__2245\ : InMux
    port map (
            O => \N__20352\,
            I => \N__20349\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__20349\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\
        );

    \I__2243\ : InMux
    port map (
            O => \N__20346\,
            I => \N__20343\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__20343\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\
        );

    \I__2241\ : InMux
    port map (
            O => \N__20340\,
            I => \N__20337\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__20337\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\
        );

    \I__2239\ : InMux
    port map (
            O => \N__20334\,
            I => \N__20331\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__20331\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__2237\ : InMux
    port map (
            O => \N__20328\,
            I => un5_counter_cry_1
        );

    \I__2236\ : InMux
    port map (
            O => \N__20325\,
            I => un5_counter_cry_2
        );

    \I__2235\ : InMux
    port map (
            O => \N__20322\,
            I => un5_counter_cry_3
        );

    \I__2234\ : InMux
    port map (
            O => \N__20319\,
            I => un5_counter_cry_4
        );

    \I__2233\ : InMux
    port map (
            O => \N__20316\,
            I => un5_counter_cry_5
        );

    \I__2232\ : InMux
    port map (
            O => \N__20313\,
            I => un5_counter_cry_6
        );

    \I__2231\ : InMux
    port map (
            O => \N__20310\,
            I => un5_counter_cry_7
        );

    \I__2230\ : CascadeMux
    port map (
            O => \N__20307\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__20304\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_\
        );

    \I__2228\ : InMux
    port map (
            O => \N__20301\,
            I => \N__20287\
        );

    \I__2227\ : InMux
    port map (
            O => \N__20300\,
            I => \N__20287\
        );

    \I__2226\ : InMux
    port map (
            O => \N__20299\,
            I => \N__20287\
        );

    \I__2225\ : InMux
    port map (
            O => \N__20298\,
            I => \N__20287\
        );

    \I__2224\ : InMux
    port map (
            O => \N__20297\,
            I => \N__20282\
        );

    \I__2223\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20282\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__20287\,
            I => \N__20279\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__20282\,
            I => \N__20276\
        );

    \I__2220\ : Span4Mux_s3_h
    port map (
            O => \N__20279\,
            I => \N__20272\
        );

    \I__2219\ : Span4Mux_s3_h
    port map (
            O => \N__20276\,
            I => \N__20269\
        );

    \I__2218\ : InMux
    port map (
            O => \N__20275\,
            I => \N__20266\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__20272\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__20269\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__20266\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2214\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20256\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__20256\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2212\ : InMux
    port map (
            O => \N__20253\,
            I => \N__20250\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__20250\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__2210\ : InMux
    port map (
            O => \N__20247\,
            I => \N__20244\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__20244\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__2208\ : InMux
    port map (
            O => \N__20241\,
            I => \N__20238\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__20238\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__20235\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\
        );

    \I__2205\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20229\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__20229\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2203\ : InMux
    port map (
            O => \N__20226\,
            I => \N__20223\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__20223\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9\
        );

    \I__2201\ : InMux
    port map (
            O => \N__20220\,
            I => \N__20215\
        );

    \I__2200\ : InMux
    port map (
            O => \N__20219\,
            I => \N__20212\
        );

    \I__2199\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20209\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__20215\,
            I => \N__20206\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__20212\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__20209\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__20206\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__20199\,
            I => \N__20196\
        );

    \I__2193\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20193\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__20193\,
            I => \N__20190\
        );

    \I__2191\ : Span4Mux_s3_h
    port map (
            O => \N__20190\,
            I => \N__20187\
        );

    \I__2190\ : Odrv4
    port map (
            O => \N__20187\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\
        );

    \I__2189\ : InMux
    port map (
            O => \N__20184\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13\
        );

    \I__2188\ : InMux
    port map (
            O => \N__20181\,
            I => \N__20178\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__20178\,
            I => \N__20174\
        );

    \I__2186\ : InMux
    port map (
            O => \N__20177\,
            I => \N__20171\
        );

    \I__2185\ : Span4Mux_v
    port map (
            O => \N__20174\,
            I => \N__20168\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__20171\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2183\ : Odrv4
    port map (
            O => \N__20168\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2182\ : InMux
    port map (
            O => \N__20163\,
            I => \N__20160\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__20160\,
            I => \N__20157\
        );

    \I__2180\ : Span4Mux_s3_h
    port map (
            O => \N__20157\,
            I => \N__20154\
        );

    \I__2179\ : Odrv4
    port map (
            O => \N__20154\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\
        );

    \I__2178\ : InMux
    port map (
            O => \N__20151\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14\
        );

    \I__2177\ : InMux
    port map (
            O => \N__20148\,
            I => \N__20141\
        );

    \I__2176\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20141\
        );

    \I__2175\ : InMux
    port map (
            O => \N__20146\,
            I => \N__20138\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__20141\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__20138\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2172\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20130\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__20130\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\
        );

    \I__2170\ : InMux
    port map (
            O => \N__20127\,
            I => \bfn_3_13_0_\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__20124\,
            I => \N__20121\
        );

    \I__2168\ : InMux
    port map (
            O => \N__20121\,
            I => \N__20118\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__20118\,
            I => \N__20113\
        );

    \I__2166\ : InMux
    port map (
            O => \N__20117\,
            I => \N__20110\
        );

    \I__2165\ : InMux
    port map (
            O => \N__20116\,
            I => \N__20107\
        );

    \I__2164\ : Span4Mux_v
    port map (
            O => \N__20113\,
            I => \N__20104\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__20110\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__20107\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__20104\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2160\ : InMux
    port map (
            O => \N__20097\,
            I => \N__20094\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__20094\,
            I => \N__20091\
        );

    \I__2158\ : Span4Mux_h
    port map (
            O => \N__20091\,
            I => \N__20088\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__20088\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\
        );

    \I__2156\ : InMux
    port map (
            O => \N__20085\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16\
        );

    \I__2155\ : InMux
    port map (
            O => \N__20082\,
            I => \N__20078\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__20081\,
            I => \N__20074\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__20078\,
            I => \N__20071\
        );

    \I__2152\ : InMux
    port map (
            O => \N__20077\,
            I => \N__20068\
        );

    \I__2151\ : InMux
    port map (
            O => \N__20074\,
            I => \N__20065\
        );

    \I__2150\ : Span4Mux_v
    port map (
            O => \N__20071\,
            I => \N__20062\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__20068\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__20065\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__20062\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2146\ : InMux
    port map (
            O => \N__20055\,
            I => \N__20052\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__20052\,
            I => \N__20049\
        );

    \I__2144\ : Odrv4
    port map (
            O => \N__20049\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\
        );

    \I__2143\ : InMux
    port map (
            O => \N__20046\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17\
        );

    \I__2142\ : InMux
    port map (
            O => \N__20043\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20037\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__20037\,
            I => \N__20034\
        );

    \I__2139\ : Odrv12
    port map (
            O => \N__20034\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\
        );

    \I__2138\ : InMux
    port map (
            O => \N__20031\,
            I => \N__20028\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__20028\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20025\,
            I => \N__20022\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__20022\,
            I => \N__20019\
        );

    \I__2134\ : Span4Mux_v
    port map (
            O => \N__20019\,
            I => \N__20016\
        );

    \I__2133\ : Odrv4
    port map (
            O => \N__20016\,
            I => \pwm_generator_inst.O_6\
        );

    \I__2132\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20010\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__20010\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_6\
        );

    \I__2130\ : InMux
    port map (
            O => \N__20007\,
            I => \N__20004\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__20004\,
            I => \N__20001\
        );

    \I__2128\ : Span4Mux_h
    port map (
            O => \N__20001\,
            I => \N__19998\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__19998\,
            I => \pwm_generator_inst.O_7\
        );

    \I__2126\ : InMux
    port map (
            O => \N__19995\,
            I => \N__19992\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__19992\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_7\
        );

    \I__2124\ : InMux
    port map (
            O => \N__19989\,
            I => \N__19986\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__19986\,
            I => \N__19983\
        );

    \I__2122\ : Span4Mux_h
    port map (
            O => \N__19983\,
            I => \N__19980\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__19980\,
            I => \pwm_generator_inst.O_8\
        );

    \I__2120\ : InMux
    port map (
            O => \N__19977\,
            I => \N__19974\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__19974\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_8\
        );

    \I__2118\ : InMux
    port map (
            O => \N__19971\,
            I => \N__19968\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__19968\,
            I => \N__19965\
        );

    \I__2116\ : Span4Mux_h
    port map (
            O => \N__19965\,
            I => \N__19962\
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__19962\,
            I => \pwm_generator_inst.O_9\
        );

    \I__2114\ : InMux
    port map (
            O => \N__19959\,
            I => \N__19956\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__19956\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_9\
        );

    \I__2112\ : InMux
    port map (
            O => \N__19953\,
            I => \N__19949\
        );

    \I__2111\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19945\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__19949\,
            I => \N__19942\
        );

    \I__2109\ : InMux
    port map (
            O => \N__19948\,
            I => \N__19939\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__19945\,
            I => \N__19936\
        );

    \I__2107\ : Span4Mux_v
    port map (
            O => \N__19942\,
            I => \N__19933\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__19939\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__19936\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__19933\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__19926\,
            I => \N__19923\
        );

    \I__2102\ : InMux
    port map (
            O => \N__19923\,
            I => \N__19920\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__19920\,
            I => \N__19917\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__19917\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\
        );

    \I__2099\ : InMux
    port map (
            O => \N__19914\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__19911\,
            I => \N__19906\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__19910\,
            I => \N__19901\
        );

    \I__2096\ : InMux
    port map (
            O => \N__19909\,
            I => \N__19897\
        );

    \I__2095\ : InMux
    port map (
            O => \N__19906\,
            I => \N__19894\
        );

    \I__2094\ : InMux
    port map (
            O => \N__19905\,
            I => \N__19887\
        );

    \I__2093\ : InMux
    port map (
            O => \N__19904\,
            I => \N__19880\
        );

    \I__2092\ : InMux
    port map (
            O => \N__19901\,
            I => \N__19880\
        );

    \I__2091\ : InMux
    port map (
            O => \N__19900\,
            I => \N__19880\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__19897\,
            I => \N__19875\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__19894\,
            I => \N__19875\
        );

    \I__2088\ : InMux
    port map (
            O => \N__19893\,
            I => \N__19866\
        );

    \I__2087\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19866\
        );

    \I__2086\ : InMux
    port map (
            O => \N__19891\,
            I => \N__19866\
        );

    \I__2085\ : InMux
    port map (
            O => \N__19890\,
            I => \N__19866\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__19887\,
            I => \N__19860\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__19880\,
            I => \N__19860\
        );

    \I__2082\ : Span4Mux_h
    port map (
            O => \N__19875\,
            I => \N__19855\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__19866\,
            I => \N__19855\
        );

    \I__2080\ : InMux
    port map (
            O => \N__19865\,
            I => \N__19852\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__19860\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__19855\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__19852\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2076\ : InMux
    port map (
            O => \N__19845\,
            I => \N__19842\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__19842\,
            I => \N__19838\
        );

    \I__2074\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19835\
        );

    \I__2073\ : Span4Mux_h
    port map (
            O => \N__19838\,
            I => \N__19830\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__19835\,
            I => \N__19830\
        );

    \I__2071\ : Odrv4
    port map (
            O => \N__19830\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__2070\ : InMux
    port map (
            O => \N__19827\,
            I => \N__19824\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__19824\,
            I => \N__19821\
        );

    \I__2068\ : Odrv12
    port map (
            O => \N__19821\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_1\
        );

    \I__2067\ : InMux
    port map (
            O => \N__19818\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_10\
        );

    \I__2066\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19812\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__19812\,
            I => \N__19807\
        );

    \I__2064\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19804\
        );

    \I__2063\ : InMux
    port map (
            O => \N__19810\,
            I => \N__19801\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__19807\,
            I => \N__19798\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__19804\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__19801\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2059\ : Odrv4
    port map (
            O => \N__19798\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__19791\,
            I => \N__19788\
        );

    \I__2057\ : InMux
    port map (
            O => \N__19788\,
            I => \N__19785\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__19785\,
            I => \N__19782\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__19782\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\
        );

    \I__2054\ : InMux
    port map (
            O => \N__19779\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11\
        );

    \I__2053\ : InMux
    port map (
            O => \N__19776\,
            I => \N__19772\
        );

    \I__2052\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19769\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__19772\,
            I => \N__19766\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__19769\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__19766\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2048\ : InMux
    port map (
            O => \N__19761\,
            I => \N__19758\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__19758\,
            I => \N__19755\
        );

    \I__2046\ : Span4Mux_v
    port map (
            O => \N__19755\,
            I => \N__19752\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__19752\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\
        );

    \I__2044\ : InMux
    port map (
            O => \N__19749\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12\
        );

    \I__2043\ : InMux
    port map (
            O => \N__19746\,
            I => \N__19743\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__19743\,
            I => \N__19740\
        );

    \I__2041\ : Span4Mux_h
    port map (
            O => \N__19740\,
            I => \N__19736\
        );

    \I__2040\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19733\
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__19736\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__19733\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__19728\,
            I => \N__19725\
        );

    \I__2036\ : InMux
    port map (
            O => \N__19725\,
            I => \N__19722\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__19722\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_8\
        );

    \I__2034\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19716\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__19716\,
            I => \N__19713\
        );

    \I__2032\ : Span4Mux_h
    port map (
            O => \N__19713\,
            I => \N__19710\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__19710\,
            I => \pwm_generator_inst.O_0\
        );

    \I__2030\ : InMux
    port map (
            O => \N__19707\,
            I => \N__19704\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__19704\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_0\
        );

    \I__2028\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19698\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__19698\,
            I => \N__19695\
        );

    \I__2026\ : Span4Mux_v
    port map (
            O => \N__19695\,
            I => \N__19692\
        );

    \I__2025\ : Odrv4
    port map (
            O => \N__19692\,
            I => \pwm_generator_inst.O_1\
        );

    \I__2024\ : InMux
    port map (
            O => \N__19689\,
            I => \N__19686\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__19686\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_1\
        );

    \I__2022\ : InMux
    port map (
            O => \N__19683\,
            I => \N__19680\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__19680\,
            I => \N__19677\
        );

    \I__2020\ : Span4Mux_h
    port map (
            O => \N__19677\,
            I => \N__19674\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__19674\,
            I => \pwm_generator_inst.O_2\
        );

    \I__2018\ : InMux
    port map (
            O => \N__19671\,
            I => \N__19668\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__19668\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_2\
        );

    \I__2016\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19662\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__19662\,
            I => \N__19659\
        );

    \I__2014\ : Span4Mux_h
    port map (
            O => \N__19659\,
            I => \N__19656\
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__19656\,
            I => \pwm_generator_inst.O_3\
        );

    \I__2012\ : InMux
    port map (
            O => \N__19653\,
            I => \N__19650\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__19650\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_3\
        );

    \I__2010\ : InMux
    port map (
            O => \N__19647\,
            I => \N__19644\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__19644\,
            I => \N__19641\
        );

    \I__2008\ : Span4Mux_v
    port map (
            O => \N__19641\,
            I => \N__19638\
        );

    \I__2007\ : Span4Mux_h
    port map (
            O => \N__19638\,
            I => \N__19635\
        );

    \I__2006\ : Odrv4
    port map (
            O => \N__19635\,
            I => \pwm_generator_inst.O_4\
        );

    \I__2005\ : InMux
    port map (
            O => \N__19632\,
            I => \N__19629\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__19629\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_4\
        );

    \I__2003\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19623\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__19623\,
            I => \N__19620\
        );

    \I__2001\ : Span12Mux_v
    port map (
            O => \N__19620\,
            I => \N__19617\
        );

    \I__2000\ : Odrv12
    port map (
            O => \N__19617\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1999\ : InMux
    port map (
            O => \N__19614\,
            I => \N__19611\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__19611\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_5\
        );

    \I__1997\ : InMux
    port map (
            O => \N__19608\,
            I => \N__19605\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__19605\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_5\
        );

    \I__1995\ : InMux
    port map (
            O => \N__19602\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_4\
        );

    \I__1994\ : InMux
    port map (
            O => \N__19599\,
            I => \N__19596\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__19596\,
            I => \N__19593\
        );

    \I__1992\ : Span4Mux_h
    port map (
            O => \N__19593\,
            I => \N__19590\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__19590\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_6\
        );

    \I__1990\ : InMux
    port map (
            O => \N__19587\,
            I => \N__19584\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__19584\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\
        );

    \I__1988\ : InMux
    port map (
            O => \N__19581\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_5\
        );

    \I__1987\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19575\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__19575\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\
        );

    \I__1985\ : InMux
    port map (
            O => \N__19572\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_6\
        );

    \I__1984\ : InMux
    port map (
            O => \N__19569\,
            I => \bfn_3_9_0_\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__19566\,
            I => \N__19563\
        );

    \I__1982\ : InMux
    port map (
            O => \N__19563\,
            I => \N__19560\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__19560\,
            I => \N__19557\
        );

    \I__1980\ : Span4Mux_v
    port map (
            O => \N__19557\,
            I => \N__19554\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__19554\,
            I => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\
        );

    \I__1978\ : InMux
    port map (
            O => \N__19551\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_8\
        );

    \I__1977\ : InMux
    port map (
            O => \N__19548\,
            I => \N__19545\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__19545\,
            I => \N__19541\
        );

    \I__1975\ : InMux
    port map (
            O => \N__19544\,
            I => \N__19538\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__19541\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__19538\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__1972\ : InMux
    port map (
            O => \N__19533\,
            I => \N__19530\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__19530\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_2\
        );

    \I__1970\ : InMux
    port map (
            O => \N__19527\,
            I => \N__19523\
        );

    \I__1969\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19520\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__19523\,
            I => \N__19517\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__19520\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__19517\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__1965\ : InMux
    port map (
            O => \N__19512\,
            I => \N__19509\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__19509\,
            I => \N__19505\
        );

    \I__1963\ : InMux
    port map (
            O => \N__19508\,
            I => \N__19502\
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__19505\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__19502\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__1960\ : InMux
    port map (
            O => \N__19497\,
            I => \N__19494\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__19494\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_7\
        );

    \I__1958\ : InMux
    port map (
            O => \N__19491\,
            I => \N__19488\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__19488\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_0\
        );

    \I__1956\ : InMux
    port map (
            O => \N__19485\,
            I => \N__19482\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__19482\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_0\
        );

    \I__1954\ : InMux
    port map (
            O => \N__19479\,
            I => \N__19476\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__19476\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\
        );

    \I__1952\ : InMux
    port map (
            O => \N__19473\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_0\
        );

    \I__1951\ : InMux
    port map (
            O => \N__19470\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_1\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__19467\,
            I => \N__19464\
        );

    \I__1949\ : InMux
    port map (
            O => \N__19464\,
            I => \N__19461\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__19461\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_3\
        );

    \I__1947\ : InMux
    port map (
            O => \N__19458\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_2\
        );

    \I__1946\ : InMux
    port map (
            O => \N__19455\,
            I => \N__19452\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__19452\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_4\
        );

    \I__1944\ : InMux
    port map (
            O => \N__19449\,
            I => \N__19446\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__19446\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\
        );

    \I__1942\ : InMux
    port map (
            O => \N__19443\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_3\
        );

    \I__1941\ : InMux
    port map (
            O => \N__19440\,
            I => \N__19437\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__19437\,
            I => \current_shift_inst.PI_CTRL.N_98\
        );

    \I__1939\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19424\
        );

    \I__1938\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19424\
        );

    \I__1937\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19424\
        );

    \I__1936\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19421\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__19424\,
            I => \N__19415\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__19421\,
            I => \N__19415\
        );

    \I__1933\ : InMux
    port map (
            O => \N__19420\,
            I => \N__19412\
        );

    \I__1932\ : Span4Mux_v
    port map (
            O => \N__19415\,
            I => \N__19409\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__19412\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__1930\ : Odrv4
    port map (
            O => \N__19409\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__19404\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_\
        );

    \I__1928\ : InMux
    port map (
            O => \N__19401\,
            I => \N__19392\
        );

    \I__1927\ : InMux
    port map (
            O => \N__19400\,
            I => \N__19383\
        );

    \I__1926\ : InMux
    port map (
            O => \N__19399\,
            I => \N__19383\
        );

    \I__1925\ : InMux
    port map (
            O => \N__19398\,
            I => \N__19383\
        );

    \I__1924\ : InMux
    port map (
            O => \N__19397\,
            I => \N__19383\
        );

    \I__1923\ : InMux
    port map (
            O => \N__19396\,
            I => \N__19377\
        );

    \I__1922\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19377\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__19392\,
            I => \N__19371\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__19383\,
            I => \N__19371\
        );

    \I__1919\ : InMux
    port map (
            O => \N__19382\,
            I => \N__19368\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__19377\,
            I => \N__19365\
        );

    \I__1917\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19362\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__19371\,
            I => \current_shift_inst.PI_CTRL.N_178\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__19368\,
            I => \current_shift_inst.PI_CTRL.N_178\
        );

    \I__1914\ : Odrv12
    port map (
            O => \N__19365\,
            I => \current_shift_inst.PI_CTRL.N_178\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__19362\,
            I => \current_shift_inst.PI_CTRL.N_178\
        );

    \I__1912\ : CascadeMux
    port map (
            O => \N__19353\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\
        );

    \I__1911\ : InMux
    port map (
            O => \N__19350\,
            I => \N__19346\
        );

    \I__1910\ : InMux
    port map (
            O => \N__19349\,
            I => \N__19343\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__19346\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__19343\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__19338\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\
        );

    \I__1906\ : InMux
    port map (
            O => \N__19335\,
            I => \N__19332\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__19332\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__1904\ : InMux
    port map (
            O => \N__19329\,
            I => \N__19326\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__19326\,
            I => \N__19323\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__19323\,
            I => un7_start_stop_0_a3
        );

    \I__1901\ : InMux
    port map (
            O => \N__19320\,
            I => \N__19317\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__19317\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\
        );

    \I__1899\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19311\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__19311\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\
        );

    \I__1897\ : InMux
    port map (
            O => \N__19308\,
            I => \bfn_2_12_0_\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__19305\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_\
        );

    \I__1895\ : InMux
    port map (
            O => \N__19302\,
            I => \N__19298\
        );

    \I__1894\ : InMux
    port map (
            O => \N__19301\,
            I => \N__19295\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__19298\,
            I => \N__19292\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__19295\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1891\ : Odrv12
    port map (
            O => \N__19292\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1890\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19281\
        );

    \I__1889\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19281\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__19281\,
            I => \N__19278\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__19278\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__19275\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__1885\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19269\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__19269\,
            I => \N__19265\
        );

    \I__1883\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19262\
        );

    \I__1882\ : Odrv12
    port map (
            O => \N__19265\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__19262\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__19257\,
            I => \current_shift_inst.PI_CTRL.N_31_cascade_\
        );

    \I__1879\ : InMux
    port map (
            O => \N__19254\,
            I => \N__19251\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__19251\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__1877\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19245\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__19245\,
            I => \N__19242\
        );

    \I__1875\ : Span4Mux_h
    port map (
            O => \N__19242\,
            I => \N__19239\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__19239\,
            I => \pwm_generator_inst.un2_threshold_acc_1_23\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__19236\,
            I => \N__19233\
        );

    \I__1872\ : InMux
    port map (
            O => \N__19233\,
            I => \N__19230\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__19230\,
            I => \N__19227\
        );

    \I__1870\ : Span4Mux_h
    port map (
            O => \N__19227\,
            I => \N__19224\
        );

    \I__1869\ : Span4Mux_v
    port map (
            O => \N__19224\,
            I => \N__19221\
        );

    \I__1868\ : Odrv4
    port map (
            O => \N__19221\,
            I => \pwm_generator_inst.un2_threshold_acc_2_8\
        );

    \I__1867\ : InMux
    port map (
            O => \N__19218\,
            I => \N__19215\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__19215\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\
        );

    \I__1865\ : InMux
    port map (
            O => \N__19212\,
            I => \bfn_2_11_0_\
        );

    \I__1864\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19206\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__19206\,
            I => \N__19203\
        );

    \I__1862\ : Span4Mux_h
    port map (
            O => \N__19203\,
            I => \N__19200\
        );

    \I__1861\ : Odrv4
    port map (
            O => \N__19200\,
            I => \pwm_generator_inst.un2_threshold_acc_1_24\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__19197\,
            I => \N__19194\
        );

    \I__1859\ : InMux
    port map (
            O => \N__19194\,
            I => \N__19191\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__19191\,
            I => \N__19188\
        );

    \I__1857\ : Span4Mux_h
    port map (
            O => \N__19188\,
            I => \N__19185\
        );

    \I__1856\ : Span4Mux_v
    port map (
            O => \N__19185\,
            I => \N__19182\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__19182\,
            I => \pwm_generator_inst.un2_threshold_acc_2_9\
        );

    \I__1854\ : InMux
    port map (
            O => \N__19179\,
            I => \N__19176\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__19176\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\
        );

    \I__1852\ : InMux
    port map (
            O => \N__19173\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__19170\,
            I => \N__19167\
        );

    \I__1850\ : InMux
    port map (
            O => \N__19167\,
            I => \N__19164\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__19164\,
            I => \N__19161\
        );

    \I__1848\ : Span4Mux_h
    port map (
            O => \N__19161\,
            I => \N__19158\
        );

    \I__1847\ : Span4Mux_v
    port map (
            O => \N__19158\,
            I => \N__19155\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__19155\,
            I => \pwm_generator_inst.un2_threshold_acc_2_10\
        );

    \I__1845\ : InMux
    port map (
            O => \N__19152\,
            I => \N__19149\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__19149\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\
        );

    \I__1843\ : InMux
    port map (
            O => \N__19146\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\
        );

    \I__1842\ : InMux
    port map (
            O => \N__19143\,
            I => \N__19140\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__19140\,
            I => \N__19137\
        );

    \I__1840\ : Span4Mux_h
    port map (
            O => \N__19137\,
            I => \N__19134\
        );

    \I__1839\ : Span4Mux_v
    port map (
            O => \N__19134\,
            I => \N__19131\
        );

    \I__1838\ : Odrv4
    port map (
            O => \N__19131\,
            I => \pwm_generator_inst.un2_threshold_acc_2_11\
        );

    \I__1837\ : InMux
    port map (
            O => \N__19128\,
            I => \N__19125\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__19125\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\
        );

    \I__1835\ : InMux
    port map (
            O => \N__19122\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__19119\,
            I => \N__19116\
        );

    \I__1833\ : InMux
    port map (
            O => \N__19116\,
            I => \N__19113\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__19113\,
            I => \N__19110\
        );

    \I__1831\ : Span4Mux_v
    port map (
            O => \N__19110\,
            I => \N__19107\
        );

    \I__1830\ : Span4Mux_v
    port map (
            O => \N__19107\,
            I => \N__19104\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__19104\,
            I => \pwm_generator_inst.un2_threshold_acc_2_12\
        );

    \I__1828\ : InMux
    port map (
            O => \N__19101\,
            I => \N__19098\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__19098\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\
        );

    \I__1826\ : InMux
    port map (
            O => \N__19095\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\
        );

    \I__1825\ : InMux
    port map (
            O => \N__19092\,
            I => \N__19089\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__19089\,
            I => \N__19086\
        );

    \I__1823\ : Span4Mux_v
    port map (
            O => \N__19086\,
            I => \N__19083\
        );

    \I__1822\ : Span4Mux_v
    port map (
            O => \N__19083\,
            I => \N__19080\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__19080\,
            I => \pwm_generator_inst.un2_threshold_acc_2_13\
        );

    \I__1820\ : InMux
    port map (
            O => \N__19077\,
            I => \N__19074\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__19074\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\
        );

    \I__1818\ : InMux
    port map (
            O => \N__19071\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__19068\,
            I => \N__19065\
        );

    \I__1816\ : InMux
    port map (
            O => \N__19065\,
            I => \N__19062\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__19062\,
            I => \N__19059\
        );

    \I__1814\ : Span4Mux_h
    port map (
            O => \N__19059\,
            I => \N__19056\
        );

    \I__1813\ : Span4Mux_v
    port map (
            O => \N__19056\,
            I => \N__19053\
        );

    \I__1812\ : Odrv4
    port map (
            O => \N__19053\,
            I => \pwm_generator_inst.un2_threshold_acc_2_14\
        );

    \I__1811\ : InMux
    port map (
            O => \N__19050\,
            I => \N__19047\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__19047\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\
        );

    \I__1809\ : InMux
    port map (
            O => \N__19044\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\
        );

    \I__1808\ : InMux
    port map (
            O => \N__19041\,
            I => \N__19038\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__19038\,
            I => \N__19035\
        );

    \I__1806\ : Span4Mux_v
    port map (
            O => \N__19035\,
            I => \N__19032\
        );

    \I__1805\ : Odrv4
    port map (
            O => \N__19032\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__19029\,
            I => \N__19022\
        );

    \I__1803\ : CascadeMux
    port map (
            O => \N__19028\,
            I => \N__19018\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__19027\,
            I => \N__19014\
        );

    \I__1801\ : InMux
    port map (
            O => \N__19026\,
            I => \N__19010\
        );

    \I__1800\ : InMux
    port map (
            O => \N__19025\,
            I => \N__19007\
        );

    \I__1799\ : InMux
    port map (
            O => \N__19022\,
            I => \N__18994\
        );

    \I__1798\ : InMux
    port map (
            O => \N__19021\,
            I => \N__18994\
        );

    \I__1797\ : InMux
    port map (
            O => \N__19018\,
            I => \N__18994\
        );

    \I__1796\ : InMux
    port map (
            O => \N__19017\,
            I => \N__18994\
        );

    \I__1795\ : InMux
    port map (
            O => \N__19014\,
            I => \N__18994\
        );

    \I__1794\ : InMux
    port map (
            O => \N__19013\,
            I => \N__18994\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__19010\,
            I => \N__18991\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__19007\,
            I => \N__18986\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__18994\,
            I => \N__18986\
        );

    \I__1790\ : Span4Mux_v
    port map (
            O => \N__18991\,
            I => \N__18983\
        );

    \I__1789\ : Span4Mux_h
    port map (
            O => \N__18986\,
            I => \N__18980\
        );

    \I__1788\ : Odrv4
    port map (
            O => \N__18983\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__18980\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1786\ : InMux
    port map (
            O => \N__18975\,
            I => \N__18972\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__18972\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\
        );

    \I__1784\ : InMux
    port map (
            O => \N__18969\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\
        );

    \I__1783\ : InMux
    port map (
            O => \N__18966\,
            I => \N__18963\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__18963\,
            I => \N__18960\
        );

    \I__1781\ : Span4Mux_h
    port map (
            O => \N__18960\,
            I => \N__18957\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__18957\,
            I => \pwm_generator_inst.un2_threshold_acc_1_16\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__18954\,
            I => \N__18951\
        );

    \I__1778\ : InMux
    port map (
            O => \N__18951\,
            I => \N__18948\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__18948\,
            I => \N__18945\
        );

    \I__1776\ : Span4Mux_h
    port map (
            O => \N__18945\,
            I => \N__18942\
        );

    \I__1775\ : Span4Mux_v
    port map (
            O => \N__18942\,
            I => \N__18939\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__18939\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__18936\,
            I => \N__18933\
        );

    \I__1772\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18930\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__18930\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\
        );

    \I__1770\ : InMux
    port map (
            O => \N__18927\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\
        );

    \I__1769\ : InMux
    port map (
            O => \N__18924\,
            I => \N__18921\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__18921\,
            I => \N__18918\
        );

    \I__1767\ : Span4Mux_h
    port map (
            O => \N__18918\,
            I => \N__18915\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__18915\,
            I => \pwm_generator_inst.un2_threshold_acc_1_17\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__18912\,
            I => \N__18909\
        );

    \I__1764\ : InMux
    port map (
            O => \N__18909\,
            I => \N__18906\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__18906\,
            I => \N__18903\
        );

    \I__1762\ : Span4Mux_h
    port map (
            O => \N__18903\,
            I => \N__18900\
        );

    \I__1761\ : Span4Mux_v
    port map (
            O => \N__18900\,
            I => \N__18897\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__18897\,
            I => \pwm_generator_inst.un2_threshold_acc_2_2\
        );

    \I__1759\ : InMux
    port map (
            O => \N__18894\,
            I => \N__18891\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__18891\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\
        );

    \I__1757\ : InMux
    port map (
            O => \N__18888\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\
        );

    \I__1756\ : InMux
    port map (
            O => \N__18885\,
            I => \N__18882\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__18882\,
            I => \N__18879\
        );

    \I__1754\ : Span4Mux_v
    port map (
            O => \N__18879\,
            I => \N__18876\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__18876\,
            I => \pwm_generator_inst.un2_threshold_acc_1_18\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__18873\,
            I => \N__18870\
        );

    \I__1751\ : InMux
    port map (
            O => \N__18870\,
            I => \N__18867\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__18867\,
            I => \N__18864\
        );

    \I__1749\ : Span4Mux_h
    port map (
            O => \N__18864\,
            I => \N__18861\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__18861\,
            I => \N__18858\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__18858\,
            I => \pwm_generator_inst.un2_threshold_acc_2_3\
        );

    \I__1746\ : InMux
    port map (
            O => \N__18855\,
            I => \N__18852\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__18852\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\
        );

    \I__1744\ : InMux
    port map (
            O => \N__18849\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\
        );

    \I__1743\ : InMux
    port map (
            O => \N__18846\,
            I => \N__18843\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__18843\,
            I => \N__18840\
        );

    \I__1741\ : Span4Mux_v
    port map (
            O => \N__18840\,
            I => \N__18837\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__18837\,
            I => \pwm_generator_inst.un2_threshold_acc_1_19\
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__18834\,
            I => \N__18831\
        );

    \I__1738\ : InMux
    port map (
            O => \N__18831\,
            I => \N__18828\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__18828\,
            I => \N__18825\
        );

    \I__1736\ : Span4Mux_v
    port map (
            O => \N__18825\,
            I => \N__18822\
        );

    \I__1735\ : Span4Mux_v
    port map (
            O => \N__18822\,
            I => \N__18819\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__18819\,
            I => \pwm_generator_inst.un2_threshold_acc_2_4\
        );

    \I__1733\ : InMux
    port map (
            O => \N__18816\,
            I => \N__18813\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__18813\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\
        );

    \I__1731\ : InMux
    port map (
            O => \N__18810\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\
        );

    \I__1730\ : InMux
    port map (
            O => \N__18807\,
            I => \N__18804\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__18804\,
            I => \N__18801\
        );

    \I__1728\ : Span4Mux_h
    port map (
            O => \N__18801\,
            I => \N__18798\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__18798\,
            I => \pwm_generator_inst.un2_threshold_acc_1_20\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__18795\,
            I => \N__18792\
        );

    \I__1725\ : InMux
    port map (
            O => \N__18792\,
            I => \N__18789\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__18789\,
            I => \N__18786\
        );

    \I__1723\ : Span4Mux_v
    port map (
            O => \N__18786\,
            I => \N__18783\
        );

    \I__1722\ : Span4Mux_v
    port map (
            O => \N__18783\,
            I => \N__18780\
        );

    \I__1721\ : Odrv4
    port map (
            O => \N__18780\,
            I => \pwm_generator_inst.un2_threshold_acc_2_5\
        );

    \I__1720\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18774\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__18774\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\
        );

    \I__1718\ : InMux
    port map (
            O => \N__18771\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\
        );

    \I__1717\ : InMux
    port map (
            O => \N__18768\,
            I => \N__18765\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__18765\,
            I => \N__18762\
        );

    \I__1715\ : Span4Mux_h
    port map (
            O => \N__18762\,
            I => \N__18759\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__18759\,
            I => \pwm_generator_inst.un2_threshold_acc_1_21\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__18756\,
            I => \N__18753\
        );

    \I__1712\ : InMux
    port map (
            O => \N__18753\,
            I => \N__18750\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__18750\,
            I => \N__18747\
        );

    \I__1710\ : Span4Mux_h
    port map (
            O => \N__18747\,
            I => \N__18744\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__18744\,
            I => \N__18741\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__18741\,
            I => \pwm_generator_inst.un2_threshold_acc_2_6\
        );

    \I__1707\ : InMux
    port map (
            O => \N__18738\,
            I => \N__18735\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__18735\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\
        );

    \I__1705\ : InMux
    port map (
            O => \N__18732\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\
        );

    \I__1704\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18726\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__18726\,
            I => \N__18723\
        );

    \I__1702\ : Span4Mux_h
    port map (
            O => \N__18723\,
            I => \N__18720\
        );

    \I__1701\ : Odrv4
    port map (
            O => \N__18720\,
            I => \pwm_generator_inst.un2_threshold_acc_1_22\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__18717\,
            I => \N__18714\
        );

    \I__1699\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18711\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__18711\,
            I => \N__18708\
        );

    \I__1697\ : Span4Mux_h
    port map (
            O => \N__18708\,
            I => \N__18705\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__18705\,
            I => \N__18702\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__18702\,
            I => \pwm_generator_inst.un2_threshold_acc_2_7\
        );

    \I__1694\ : InMux
    port map (
            O => \N__18699\,
            I => \N__18696\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__18696\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\
        );

    \I__1692\ : InMux
    port map (
            O => \N__18693\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\
        );

    \I__1691\ : InMux
    port map (
            O => \N__18690\,
            I => \N__18684\
        );

    \I__1690\ : InMux
    port map (
            O => \N__18689\,
            I => \N__18684\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__18684\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__18681\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\
        );

    \I__1687\ : InMux
    port map (
            O => \N__18678\,
            I => \N__18675\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__18675\,
            I => \N__18672\
        );

    \I__1685\ : Span4Mux_v
    port map (
            O => \N__18672\,
            I => \N__18668\
        );

    \I__1684\ : InMux
    port map (
            O => \N__18671\,
            I => \N__18665\
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__18668\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__18665\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1681\ : InMux
    port map (
            O => \N__18660\,
            I => \N__18654\
        );

    \I__1680\ : InMux
    port map (
            O => \N__18659\,
            I => \N__18654\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__18654\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__18651\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13_cascade_\
        );

    \I__1677\ : InMux
    port map (
            O => \N__18648\,
            I => \N__18645\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__18645\,
            I => \N__18642\
        );

    \I__1675\ : Span4Mux_h
    port map (
            O => \N__18642\,
            I => \N__18639\
        );

    \I__1674\ : Span4Mux_v
    port map (
            O => \N__18639\,
            I => \N__18636\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__18636\,
            I => \pwm_generator_inst.un2_threshold_acc_2_0\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__18633\,
            I => \N__18630\
        );

    \I__1671\ : InMux
    port map (
            O => \N__18630\,
            I => \N__18627\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__18627\,
            I => \N__18624\
        );

    \I__1669\ : Span4Mux_h
    port map (
            O => \N__18624\,
            I => \N__18621\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__18621\,
            I => \pwm_generator_inst.un2_threshold_acc_1_15\
        );

    \I__1667\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18615\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__18615\,
            I => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\
        );

    \I__1665\ : InMux
    port map (
            O => \N__18612\,
            I => \N__18606\
        );

    \I__1664\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18606\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__18606\,
            I => \N__18602\
        );

    \I__1662\ : InMux
    port map (
            O => \N__18605\,
            I => \N__18599\
        );

    \I__1661\ : Odrv12
    port map (
            O => \N__18602\,
            I => pwm_duty_input_9
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__18599\,
            I => pwm_duty_input_9
        );

    \I__1659\ : CascadeMux
    port map (
            O => \N__18594\,
            I => \N__18590\
        );

    \I__1658\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18585\
        );

    \I__1657\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18585\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__18585\,
            I => \N__18581\
        );

    \I__1655\ : InMux
    port map (
            O => \N__18584\,
            I => \N__18578\
        );

    \I__1654\ : Odrv12
    port map (
            O => \N__18581\,
            I => pwm_duty_input_8
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__18578\,
            I => pwm_duty_input_8
        );

    \I__1652\ : InMux
    port map (
            O => \N__18573\,
            I => \N__18570\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__18570\,
            I => \N_22_i_i\
        );

    \I__1650\ : InMux
    port map (
            O => \N__18567\,
            I => \N__18564\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__18564\,
            I => \current_shift_inst.PI_CTRL.m14_2\
        );

    \I__1648\ : InMux
    port map (
            O => \N__18561\,
            I => \N__18550\
        );

    \I__1647\ : InMux
    port map (
            O => \N__18560\,
            I => \N__18550\
        );

    \I__1646\ : InMux
    port map (
            O => \N__18559\,
            I => \N__18547\
        );

    \I__1645\ : InMux
    port map (
            O => \N__18558\,
            I => \N__18540\
        );

    \I__1644\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18540\
        );

    \I__1643\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18540\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__18555\,
            I => \N__18537\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__18550\,
            I => \N__18517\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__18547\,
            I => \N__18512\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__18540\,
            I => \N__18512\
        );

    \I__1638\ : InMux
    port map (
            O => \N__18537\,
            I => \N__18509\
        );

    \I__1637\ : InMux
    port map (
            O => \N__18536\,
            I => \N__18506\
        );

    \I__1636\ : InMux
    port map (
            O => \N__18535\,
            I => \N__18503\
        );

    \I__1635\ : InMux
    port map (
            O => \N__18534\,
            I => \N__18486\
        );

    \I__1634\ : InMux
    port map (
            O => \N__18533\,
            I => \N__18486\
        );

    \I__1633\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18486\
        );

    \I__1632\ : InMux
    port map (
            O => \N__18531\,
            I => \N__18486\
        );

    \I__1631\ : InMux
    port map (
            O => \N__18530\,
            I => \N__18486\
        );

    \I__1630\ : InMux
    port map (
            O => \N__18529\,
            I => \N__18486\
        );

    \I__1629\ : InMux
    port map (
            O => \N__18528\,
            I => \N__18486\
        );

    \I__1628\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18486\
        );

    \I__1627\ : InMux
    port map (
            O => \N__18526\,
            I => \N__18471\
        );

    \I__1626\ : InMux
    port map (
            O => \N__18525\,
            I => \N__18471\
        );

    \I__1625\ : InMux
    port map (
            O => \N__18524\,
            I => \N__18471\
        );

    \I__1624\ : InMux
    port map (
            O => \N__18523\,
            I => \N__18471\
        );

    \I__1623\ : InMux
    port map (
            O => \N__18522\,
            I => \N__18471\
        );

    \I__1622\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18471\
        );

    \I__1621\ : InMux
    port map (
            O => \N__18520\,
            I => \N__18471\
        );

    \I__1620\ : Span4Mux_v
    port map (
            O => \N__18517\,
            I => \N__18466\
        );

    \I__1619\ : Span4Mux_v
    port map (
            O => \N__18512\,
            I => \N__18466\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__18509\,
            I => pwm_duty_input_10
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__18506\,
            I => pwm_duty_input_10
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__18503\,
            I => pwm_duty_input_10
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__18486\,
            I => pwm_duty_input_10
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__18471\,
            I => pwm_duty_input_10
        );

    \I__1613\ : Odrv4
    port map (
            O => \N__18466\,
            I => pwm_duty_input_10
        );

    \I__1612\ : InMux
    port map (
            O => \N__18453\,
            I => \N__18448\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__18452\,
            I => \N__18445\
        );

    \I__1610\ : InMux
    port map (
            O => \N__18451\,
            I => \N__18442\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__18448\,
            I => \N__18439\
        );

    \I__1608\ : InMux
    port map (
            O => \N__18445\,
            I => \N__18436\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__18442\,
            I => \N__18433\
        );

    \I__1606\ : Span4Mux_v
    port map (
            O => \N__18439\,
            I => \N__18430\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__18436\,
            I => \N__18427\
        );

    \I__1604\ : Span4Mux_s1_h
    port map (
            O => \N__18433\,
            I => \N__18424\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__18430\,
            I => pwm_duty_input_4
        );

    \I__1602\ : Odrv12
    port map (
            O => \N__18427\,
            I => pwm_duty_input_4
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__18424\,
            I => pwm_duty_input_4
        );

    \I__1600\ : InMux
    port map (
            O => \N__18417\,
            I => \N__18414\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__18414\,
            I => \N__18410\
        );

    \I__1598\ : InMux
    port map (
            O => \N__18413\,
            I => \N__18407\
        );

    \I__1597\ : Span4Mux_v
    port map (
            O => \N__18410\,
            I => \N__18404\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__18407\,
            I => pwm_duty_input_1
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__18404\,
            I => pwm_duty_input_1
        );

    \I__1594\ : InMux
    port map (
            O => \N__18399\,
            I => \N__18396\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__18396\,
            I => \N__18392\
        );

    \I__1592\ : InMux
    port map (
            O => \N__18395\,
            I => \N__18389\
        );

    \I__1591\ : Span4Mux_v
    port map (
            O => \N__18392\,
            I => \N__18386\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__18389\,
            I => pwm_duty_input_2
        );

    \I__1589\ : Odrv4
    port map (
            O => \N__18386\,
            I => pwm_duty_input_2
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__18381\,
            I => \N__18377\
        );

    \I__1587\ : InMux
    port map (
            O => \N__18380\,
            I => \N__18374\
        );

    \I__1586\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18371\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__18374\,
            I => \N__18368\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__18371\,
            I => \N__18363\
        );

    \I__1583\ : Span4Mux_v
    port map (
            O => \N__18368\,
            I => \N__18363\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__18363\,
            I => pwm_duty_input_0
        );

    \I__1581\ : InMux
    port map (
            O => \N__18360\,
            I => \N__18356\
        );

    \I__1580\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18353\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__18356\,
            I => \N__18350\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__18353\,
            I => \N__18346\
        );

    \I__1577\ : Span4Mux_h
    port map (
            O => \N__18350\,
            I => \N__18343\
        );

    \I__1576\ : InMux
    port map (
            O => \N__18349\,
            I => \N__18340\
        );

    \I__1575\ : Odrv12
    port map (
            O => \N__18346\,
            I => pwm_duty_input_3
        );

    \I__1574\ : Odrv4
    port map (
            O => \N__18343\,
            I => pwm_duty_input_3
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__18340\,
            I => pwm_duty_input_3
        );

    \I__1572\ : InMux
    port map (
            O => \N__18333\,
            I => \N__18330\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__18330\,
            I => \current_shift_inst.PI_CTRL.N_19\
        );

    \I__1570\ : InMux
    port map (
            O => \N__18327\,
            I => \N__18318\
        );

    \I__1569\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18318\
        );

    \I__1568\ : InMux
    port map (
            O => \N__18325\,
            I => \N__18318\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__18318\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \I__1566\ : InMux
    port map (
            O => \N__18315\,
            I => \N__18306\
        );

    \I__1565\ : InMux
    port map (
            O => \N__18314\,
            I => \N__18306\
        );

    \I__1564\ : InMux
    port map (
            O => \N__18313\,
            I => \N__18306\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__18306\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1562\ : InMux
    port map (
            O => \N__18303\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19\
        );

    \I__1561\ : InMux
    port map (
            O => \N__18300\,
            I => \N__18297\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__18297\,
            I => \N__18294\
        );

    \I__1559\ : Span4Mux_v
    port map (
            O => \N__18294\,
            I => \N__18290\
        );

    \I__1558\ : InMux
    port map (
            O => \N__18293\,
            I => \N__18287\
        );

    \I__1557\ : Odrv4
    port map (
            O => \N__18290\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__18287\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__18282\,
            I => \N__18279\
        );

    \I__1554\ : InMux
    port map (
            O => \N__18279\,
            I => \N__18276\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__18276\,
            I => \N__18273\
        );

    \I__1552\ : Span4Mux_v
    port map (
            O => \N__18273\,
            I => \N__18270\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__18270\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_16\
        );

    \I__1550\ : InMux
    port map (
            O => \N__18267\,
            I => \N__18261\
        );

    \I__1549\ : InMux
    port map (
            O => \N__18266\,
            I => \N__18261\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__18261\,
            I => \N__18257\
        );

    \I__1547\ : InMux
    port map (
            O => \N__18260\,
            I => \N__18254\
        );

    \I__1546\ : Odrv12
    port map (
            O => \N__18257\,
            I => pwm_duty_input_7
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__18254\,
            I => pwm_duty_input_7
        );

    \I__1544\ : InMux
    port map (
            O => \N__18249\,
            I => \N__18243\
        );

    \I__1543\ : InMux
    port map (
            O => \N__18248\,
            I => \N__18243\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__18243\,
            I => \N__18239\
        );

    \I__1541\ : InMux
    port map (
            O => \N__18242\,
            I => \N__18236\
        );

    \I__1540\ : Odrv12
    port map (
            O => \N__18239\,
            I => pwm_duty_input_5
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__18236\,
            I => pwm_duty_input_5
        );

    \I__1538\ : InMux
    port map (
            O => \N__18231\,
            I => \bfn_1_10_0_\
        );

    \I__1537\ : InMux
    port map (
            O => \N__18228\,
            I => \N__18225\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__18225\,
            I => \N__18222\
        );

    \I__1535\ : Odrv4
    port map (
            O => \N__18222\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1534\ : InMux
    port map (
            O => \N__18219\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0\
        );

    \I__1533\ : InMux
    port map (
            O => \N__18216\,
            I => \N__18213\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__18213\,
            I => \N__18210\
        );

    \I__1531\ : Odrv4
    port map (
            O => \N__18210\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1530\ : InMux
    port map (
            O => \N__18207\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1\
        );

    \I__1529\ : InMux
    port map (
            O => \N__18204\,
            I => \N__18201\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__18201\,
            I => \N__18198\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__18198\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1526\ : InMux
    port map (
            O => \N__18195\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2\
        );

    \I__1525\ : InMux
    port map (
            O => \N__18192\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3\
        );

    \I__1524\ : InMux
    port map (
            O => \N__18189\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4\
        );

    \I__1523\ : InMux
    port map (
            O => \N__18186\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5\
        );

    \I__1522\ : InMux
    port map (
            O => \N__18183\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6\
        );

    \I__1521\ : CascadeMux
    port map (
            O => \N__18180\,
            I => \current_shift_inst.PI_CTRL.m7_2_cascade_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_6\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_14\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_22\,
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_30\,
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_4_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_5_0_\
        );

    \IN_MUX_bfv_4_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_counter_cry_8,
            carryinitout => \bfn_4_6_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_16_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_16_12_0_\
        );

    \IN_MUX_bfv_16_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_16_13_0_\
        );

    \IN_MUX_bfv_18_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_11_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_18_16_0_\
        );

    \IN_MUX_bfv_12_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_7_0_\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_12_8_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_14_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_5_0_\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_5_cry_8\,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_5_cry_16\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_5_cry_24\,
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_3_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_11_0_\
        );

    \IN_MUX_bfv_3_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            carryinitout => \bfn_3_12_0_\
        );

    \IN_MUX_bfv_3_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            carryinitout => \bfn_3_13_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_3_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_8_0_\
        );

    \IN_MUX_bfv_3_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            carryinitout => \bfn_3_9_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_16_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_18_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_16_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_16_20_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_18_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_7_0_\
        );

    \IN_MUX_bfv_18_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_18_8_0_\
        );

    \IN_MUX_bfv_18_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_18_9_0_\
        );

    \IN_MUX_bfv_18_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_18_10_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_cry_7\,
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_cry_15\,
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_10_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_cry_23\,
            carryinitout => \bfn_10_20_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_cry_8\,
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_cry_16\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_cry_24\,
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_12_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_12_21_0_\
        );

    \IN_MUX_bfv_12_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_12_22_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.counter_cry_7\,
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_7_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.counter_cry_15\,
            carryinitout => \bfn_7_21_0_\
        );

    \IN_MUX_bfv_7_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.counter_cry_23\,
            carryinitout => \bfn_7_22_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_7\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_15\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_23\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_4_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryinitout => \bfn_4_15_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryinitout => \bfn_4_16_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryinitout => \bfn_5_13_0_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__33852\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_335_i_g\
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__29022\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_187_i_g\
        );

    \current_shift_inst.timer_phase.running_RNIC90O_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__32373\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_phase.N_188_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__27531\,
            CLKHFEN => \N__27535\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__27556\,
            RGB2PWM => \N__18573\,
            RGB1 => rgb_g_wire,
            CURREN => \N__27595\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__19329\,
            RGB0PWM => \N__46987\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21300\,
            lcout => pwm_duty_input_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47463\,
            ce => \N__24483\,
            sr => \N__46905\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__19026\,
            in1 => \N__18293\,
            in2 => \_gnd_net_\,
            in3 => \N__18535\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18611\,
            in1 => \N__18266\,
            in2 => \N__18594\,
            in3 => \N__18248\,
            lcout => \current_shift_inst.PI_CTRL.m14_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__18249\,
            in1 => \N__18359\,
            in2 => \N__18452\,
            in3 => \N__18612\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.m7_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__18593\,
            in1 => \N__18536\,
            in2 => \N__18180\,
            in3 => \N__18267\,
            lcout => i8_mux,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__18325\,
            in1 => \N__19432\,
            in2 => \N__20592\,
            in3 => \N__18313\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47460\,
            ce => \N__24465\,
            sr => \N__46918\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__18326\,
            in1 => \N__19433\,
            in2 => \N__20898\,
            in3 => \N__18314\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47460\,
            ce => \N__24465\,
            sr => \N__46918\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__18327\,
            in1 => \N__19434\,
            in2 => \N__20871\,
            in3 => \N__18315\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47460\,
            ce => \N__24465\,
            sr => \N__46918\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19841\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18228\,
            in2 => \_gnd_net_\,
            in3 => \N__18219\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18216\,
            in2 => \_gnd_net_\,
            in3 => \N__18207\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18204\,
            in2 => \_gnd_net_\,
            in3 => \N__18195\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18618\,
            in2 => \_gnd_net_\,
            in3 => \N__18192\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27716\,
            in2 => \N__18936\,
            in3 => \N__18189\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18894\,
            in2 => \N__27776\,
            in3 => \N__18186\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18855\,
            in2 => \N__27777\,
            in3 => \N__18183\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18816\,
            in2 => \_gnd_net_\,
            in3 => \N__18231\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18777\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18738\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18699\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19218\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19179\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19152\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19128\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19101\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19077\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19050\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18975\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18303\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18671\,
            in2 => \_gnd_net_\,
            in3 => \N__19948\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000111100"
        )
    port map (
            in0 => \N__18300\,
            in1 => \N__19025\,
            in2 => \N__18282\,
            in3 => \N__18559\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__19399\,
            in1 => \N__21293\,
            in2 => \N__20679\,
            in3 => \N__20300\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47446\,
            ce => \N__24500\,
            sr => \N__46935\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__19401\,
            in1 => \N__19301\,
            in2 => \N__20846\,
            in3 => \N__19420\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47446\,
            ce => \N__24500\,
            sr => \N__46935\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__19397\,
            in1 => \N__21291\,
            in2 => \N__20763\,
            in3 => \N__20298\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47446\,
            ce => \N__24500\,
            sr => \N__46935\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__19398\,
            in1 => \N__21292\,
            in2 => \N__20730\,
            in3 => \N__20299\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47446\,
            ce => \N__24500\,
            sr => \N__46935\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__19400\,
            in1 => \N__21294\,
            in2 => \N__21063\,
            in3 => \N__20301\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47446\,
            ce => \N__24500\,
            sr => \N__46935\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__20297\,
            in1 => \N__19254\,
            in2 => \N__20811\,
            in3 => \N__19350\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47439\,
            ce => \N__24510\,
            sr => \N__46939\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__19382\,
            in1 => \N__21295\,
            in2 => \N__20640\,
            in3 => \N__20296\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47439\,
            ce => \N__24510\,
            sr => \N__46939\
        );

    \current_shift_inst.N_22_i_i_LC_1_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__35073\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46986\,
            lcout => \N_22_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__18333\,
            in1 => \N__18567\,
            in2 => \N__18555\,
            in3 => \N__18453\,
            lcout => \N_28_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__18413\,
            in1 => \N__18395\,
            in2 => \N__18381\,
            in3 => \N__18360\,
            lcout => \current_shift_inst.PI_CTRL.N_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__21296\,
            in1 => \N__19395\,
            in2 => \_gnd_net_\,
            in3 => \N__19272\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000100"
        )
    port map (
            in0 => \N__19396\,
            in1 => \N__19302\,
            in2 => \N__20850\,
            in3 => \N__19431\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19811\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19544\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__20218\,
            in1 => \N__19526\,
            in2 => \N__20199\,
            in3 => \N__19892\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20177\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18689\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_15\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__18690\,
            in1 => \N__20163\,
            in2 => \N__18681\,
            in3 => \N__19893\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20077\,
            in2 => \_gnd_net_\,
            in3 => \N__19739\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__18678\,
            in1 => \N__19952\,
            in2 => \N__19926\,
            in3 => \N__19890\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19775\,
            in2 => \_gnd_net_\,
            in3 => \N__18659\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_13\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__18660\,
            in1 => \N__19761\,
            in2 => \N__18651\,
            in3 => \N__19891\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20117\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19508\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18648\,
            in2 => \N__18633\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18966\,
            in2 => \N__18954\,
            in3 => \N__18927\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18924\,
            in2 => \N__18912\,
            in3 => \N__18888\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18885\,
            in2 => \N__18873\,
            in3 => \N__18849\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18846\,
            in2 => \N__18834\,
            in3 => \N__18810\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18807\,
            in2 => \N__18795\,
            in3 => \N__18771\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18768\,
            in2 => \N__18756\,
            in3 => \N__18732\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18729\,
            in2 => \N__18717\,
            in3 => \N__18693\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19248\,
            in2 => \N__19236\,
            in3 => \N__19212\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19209\,
            in2 => \N__19197\,
            in3 => \N__19173\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19013\,
            in2 => \N__19170\,
            in3 => \N__19146\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19143\,
            in2 => \N__19027\,
            in3 => \N__19122\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19017\,
            in2 => \N__19119\,
            in3 => \N__19095\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19092\,
            in2 => \N__19028\,
            in3 => \N__19071\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19021\,
            in2 => \N__19068\,
            in3 => \N__19044\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19041\,
            in2 => \N__19029\,
            in3 => \N__18969\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19320\,
            in1 => \N__19314\,
            in2 => \_gnd_net_\,
            in3 => \N__19308\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\,
            ltout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__19287\,
            in1 => \N__20133\,
            in2 => \N__19305\,
            in3 => \N__20147\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20809\,
            in2 => \_gnd_net_\,
            in3 => \N__20836\,
            lcout => \current_shift_inst.PI_CTRL.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__21266\,
            in1 => \N__20810\,
            in2 => \_gnd_net_\,
            in3 => \N__19268\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20148\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19286\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20749\,
            in2 => \_gnd_net_\,
            in3 => \N__21059\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__20674\,
            in1 => \N__20722\,
            in2 => \N__19275\,
            in3 => \N__20633\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => \current_shift_inst.PI_CTRL.N_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__21265\,
            in1 => \N__20805\,
            in2 => \N__19257\,
            in3 => \N__19376\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__19440\,
            in1 => \N__19349\,
            in2 => \N__21284\,
            in3 => \N__20275\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIOLF4_14_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20964\,
            in1 => \N__21354\,
            in2 => \N__21330\,
            in3 => \N__21387\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20031\,
            in1 => \N__19335\,
            in2 => \N__19404\,
            in3 => \N__20232\,
            lcout => \current_shift_inst.PI_CTRL.N_178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIV2LD_8_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20626\,
            in2 => \_gnd_net_\,
            in3 => \N__21055\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20675\,
            in1 => \N__20723\,
            in2 => \N__19353\,
            in3 => \N__20756\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_15_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20946\,
            in2 => \_gnd_net_\,
            in3 => \N__21144\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI2QR8_10_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21126\,
            in1 => \N__20334\,
            in2 => \N__19338\,
            in3 => \N__21030\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un7_start_stop_0_a3_LC_2_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35072\,
            in2 => \_gnd_net_\,
            in3 => \N__46985\,
            lcout => un7_start_stop_0_a3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_6_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__20435\,
            in1 => \N__20550\,
            in2 => \N__20499\,
            in3 => \N__19587\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__46892\
        );

    \pwm_generator_inst.threshold_0_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19491\,
            lcout => \pwm_generator_inst.thresholdZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__46892\
        );

    \pwm_generator_inst.threshold_ACC_7_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__20436\,
            in1 => \N__20551\,
            in2 => \N__20500\,
            in3 => \N__19578\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__46892\
        );

    \pwm_generator_inst.threshold_ACC_0_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000001100"
        )
    port map (
            in0 => \N__20434\,
            in1 => \N__19479\,
            in2 => \N__20498\,
            in3 => \N__20549\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__46892\
        );

    \pwm_generator_inst.threshold_ACC_4_LC_3_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__20548\,
            in1 => \N__20482\,
            in2 => \N__20447\,
            in3 => \N__19449\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__46892\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19485\,
            in2 => \N__19911\,
            in3 => \N__19909\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_8_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19827\,
            in2 => \_gnd_net_\,
            in3 => \N__19473\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19533\,
            in2 => \_gnd_net_\,
            in3 => \N__19470\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19467\,
            in3 => \N__19458\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19455\,
            in2 => \_gnd_net_\,
            in3 => \N__19443\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19608\,
            in2 => \_gnd_net_\,
            in3 => \N__19602\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19599\,
            in2 => \_gnd_net_\,
            in3 => \N__19581\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19497\,
            in2 => \_gnd_net_\,
            in3 => \N__19572\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19728\,
            in3 => \N__19569\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_3_9_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__19904\,
            in1 => \N__20040\,
            in2 => \N__19566\,
            in3 => \N__19551\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__19900\,
            in1 => \N__19548\,
            in2 => \N__19791\,
            in3 => \N__19810\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20219\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19527\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__20097\,
            in1 => \N__20116\,
            in2 => \N__19910\,
            in3 => \N__19512\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__19905\,
            in1 => \N__19746\,
            in2 => \N__20081\,
            in3 => \N__20055\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__37410\,
            in1 => \N__40893\,
            in2 => \_gnd_net_\,
            in3 => \N__37680\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47447\,
            ce => \N__30888\,
            sr => \N__46919\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19707\,
            in2 => \_gnd_net_\,
            in3 => \N__19719\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_3_11_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19689\,
            in2 => \_gnd_net_\,
            in3 => \N__19701\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19671\,
            in2 => \_gnd_net_\,
            in3 => \N__19683\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19653\,
            in2 => \_gnd_net_\,
            in3 => \N__19665\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19632\,
            in2 => \_gnd_net_\,
            in3 => \N__19647\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19614\,
            in2 => \_gnd_net_\,
            in3 => \N__19626\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20013\,
            in2 => \_gnd_net_\,
            in3 => \N__20025\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19995\,
            in2 => \_gnd_net_\,
            in3 => \N__20007\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19977\,
            in2 => \_gnd_net_\,
            in3 => \N__19989\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_3_12_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19959\,
            in2 => \_gnd_net_\,
            in3 => \N__19971\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19953\,
            in2 => \_gnd_net_\,
            in3 => \N__19914\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__19865\,
            in1 => \N__19845\,
            in2 => \_gnd_net_\,
            in3 => \N__19818\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19815\,
            in2 => \_gnd_net_\,
            in3 => \N__19779\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19776\,
            in2 => \_gnd_net_\,
            in3 => \N__19749\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20220\,
            in2 => \_gnd_net_\,
            in3 => \N__20184\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20181\,
            in2 => \_gnd_net_\,
            in3 => \N__20151\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20146\,
            in2 => \_gnd_net_\,
            in3 => \N__20127\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_3_13_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20124\,
            in3 => \N__20085\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20082\,
            in2 => \_gnd_net_\,
            in3 => \N__20046\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20043\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIC5B4_11_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20994\,
            in1 => \N__20925\,
            in2 => \N__21009\,
            in3 => \N__20981\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIG72_10_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21323\,
            in2 => \_gnd_net_\,
            in3 => \N__21023\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRKT8_11_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21386\,
            in1 => \N__21005\,
            in2 => \N__20307\,
            in3 => \N__20247\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20241\,
            in1 => \N__20253\,
            in2 => \N__20304\,
            in3 => \N__20259\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3DG5_12_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20993\,
            in1 => \N__20960\,
            in2 => \N__21105\,
            in3 => \N__20226\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIOIC4_15_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21194\,
            in1 => \N__21206\,
            in2 => \N__21125\,
            in3 => \N__20939\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGDF4_20_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21140\,
            in1 => \N__21155\,
            in2 => \N__21350\,
            in3 => \N__21170\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIOJD4_13_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21081\,
            in1 => \N__20924\,
            in2 => \N__20982\,
            in3 => \N__21365\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21207\,
            in2 => \_gnd_net_\,
            in3 => \N__21171\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8JH5_19_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21183\,
            in1 => \N__21366\,
            in2 => \N__20235\,
            in3 => \N__21080\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0U62_19_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21398\,
            in2 => \_gnd_net_\,
            in3 => \N__21182\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMIE4_18_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21399\,
            in1 => \N__21101\,
            in2 => \N__21159\,
            in3 => \N__21195\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_counter_cry_1_c_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21581\,
            in2 => \N__22077\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_5_0_\,
            carryout => un5_counter_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21594\,
            in2 => \_gnd_net_\,
            in3 => \N__20328\,
            lcout => \counterZ0Z_2\,
            ltout => OPEN,
            carryin => un5_counter_cry_1,
            carryout => un5_counter_cry_2,
            clk => \N__47461\,
            ce => 'H',
            sr => \N__46866\
        );

    \counter_3_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21486\,
            in2 => \_gnd_net_\,
            in3 => \N__20325\,
            lcout => \counterZ0Z_3\,
            ltout => OPEN,
            carryin => un5_counter_cry_2,
            carryout => un5_counter_cry_3,
            clk => \N__47461\,
            ce => 'H',
            sr => \N__46866\
        );

    \counter_4_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21513\,
            in2 => \_gnd_net_\,
            in3 => \N__20322\,
            lcout => \counterZ0Z_4\,
            ltout => OPEN,
            carryin => un5_counter_cry_3,
            carryout => un5_counter_cry_4,
            clk => \N__47461\,
            ce => 'H',
            sr => \N__46866\
        );

    \counter_5_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21525\,
            in2 => \_gnd_net_\,
            in3 => \N__20319\,
            lcout => \counterZ0Z_5\,
            ltout => OPEN,
            carryin => un5_counter_cry_4,
            carryout => un5_counter_cry_5,
            clk => \N__47461\,
            ce => 'H',
            sr => \N__46866\
        );

    \counter_6_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21500\,
            in2 => \_gnd_net_\,
            in3 => \N__20316\,
            lcout => \counterZ0Z_6\,
            ltout => OPEN,
            carryin => un5_counter_cry_5,
            carryout => un5_counter_cry_6,
            clk => \N__47461\,
            ce => 'H',
            sr => \N__46866\
        );

    \counter_RNO_0_7_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21219\,
            in2 => \_gnd_net_\,
            in3 => \N__20313\,
            lcout => \counter_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => un5_counter_cry_6,
            carryout => un5_counter_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_8_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21561\,
            in2 => \_gnd_net_\,
            in3 => \N__20310\,
            lcout => \counterZ0Z_8\,
            ltout => OPEN,
            carryin => un5_counter_cry_7,
            carryout => un5_counter_cry_8,
            clk => \N__47461\,
            ce => 'H',
            sr => \N__46866\
        );

    \counter_9_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21537\,
            in2 => \_gnd_net_\,
            in3 => \N__20370\,
            lcout => \counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_4_6_0_\,
            carryout => un5_counter_cry_9,
            clk => \N__47459\,
            ce => 'H',
            sr => \N__46876\
        );

    \counter_RNO_0_10_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21411\,
            in2 => \_gnd_net_\,
            in3 => \N__20367\,
            lcout => \counter_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => un5_counter_cry_9,
            carryout => un5_counter_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_11_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21549\,
            in2 => \_gnd_net_\,
            in3 => \N__20364\,
            lcout => \counterZ0Z_11\,
            ltout => OPEN,
            carryin => un5_counter_cry_10,
            carryout => un5_counter_cry_11,
            clk => \N__47459\,
            ce => 'H',
            sr => \N__46876\
        );

    \counter_RNO_0_12_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21434\,
            in2 => \_gnd_net_\,
            in3 => \N__20361\,
            lcout => \counter_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_2_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__20552\,
            in1 => \N__20490\,
            in2 => \N__20444\,
            in3 => \N__20358\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47453\,
            ce => 'H',
            sr => \N__46885\
        );

    \pwm_generator_inst.threshold_ACC_3_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__20553\,
            in1 => \N__20491\,
            in2 => \N__20445\,
            in3 => \N__20352\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47453\,
            ce => 'H',
            sr => \N__46885\
        );

    \pwm_generator_inst.threshold_ACC_1_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111001010"
        )
    port map (
            in0 => \N__20489\,
            in1 => \N__20424\,
            in2 => \N__20563\,
            in3 => \N__20346\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47453\,
            ce => 'H',
            sr => \N__46885\
        );

    \pwm_generator_inst.threshold_ACC_5_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__20554\,
            in1 => \N__20492\,
            in2 => \N__20446\,
            in3 => \N__20340\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47453\,
            ce => 'H',
            sr => \N__46885\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25344\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47451\,
            ce => \N__24466\,
            sr => \N__46893\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25284\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47451\,
            ce => \N__24466\,
            sr => \N__46893\
        );

    \pwm_generator_inst.threshold_ACC_8_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__20501\,
            in1 => \N__20565\,
            in2 => \N__20574\,
            in3 => \N__20440\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__46906\
        );

    \pwm_generator_inst.threshold_ACC_9_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__20564\,
            in1 => \N__20502\,
            in2 => \N__20448\,
            in3 => \N__20382\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__46906\
        );

    \pwm_generator_inst.threshold_9_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20376\,
            lcout => \pwm_generator_inst.thresholdZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__46906\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011010000"
        )
    port map (
            in0 => \N__24653\,
            in1 => \N__21672\,
            in2 => \N__24885\,
            in3 => \N__24977\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47440\,
            ce => \N__24485\,
            sr => \N__46912\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110100001101"
        )
    port map (
            in0 => \N__24978\,
            in1 => \N__21663\,
            in2 => \N__24890\,
            in3 => \N__24654\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47440\,
            ce => \N__24485\,
            sr => \N__46912\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110010001111"
        )
    port map (
            in0 => \N__24655\,
            in1 => \N__21654\,
            in2 => \N__24886\,
            in3 => \N__24979\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47440\,
            ce => \N__24485\,
            sr => \N__46912\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110100001101"
        )
    port map (
            in0 => \N__24980\,
            in1 => \N__21645\,
            in2 => \N__24891\,
            in3 => \N__24656\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47440\,
            ce => \N__24485\,
            sr => \N__46912\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110010001111"
        )
    port map (
            in0 => \N__24657\,
            in1 => \N__21834\,
            in2 => \N__24887\,
            in3 => \N__24981\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47440\,
            ce => \N__24485\,
            sr => \N__46912\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000100110001"
        )
    port map (
            in0 => \N__24982\,
            in1 => \N__24840\,
            in2 => \N__21825\,
            in3 => \N__24658\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47440\,
            ce => \N__24485\,
            sr => \N__46912\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24257\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47440\,
            ce => \N__24485\,
            sr => \N__46912\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011111"
        )
    port map (
            in0 => \N__21698\,
            in1 => \N__21721\,
            in2 => \N__22528\,
            in3 => \N__21745\,
            lcout => \current_shift_inst.PI_CTRL.N_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__21942\,
            in1 => \N__24659\,
            in2 => \N__24892\,
            in3 => \N__25023\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47431\,
            ce => \N__24492\,
            sr => \N__46920\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011010000"
        )
    port map (
            in0 => \N__24662\,
            in1 => \N__21861\,
            in2 => \N__24889\,
            in3 => \N__25026\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47424\,
            ce => \N__24468\,
            sr => \N__46924\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24282\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47424\,
            ce => \N__24468\,
            sr => \N__46924\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011010000"
        )
    port map (
            in0 => \N__24660\,
            in1 => \N__21882\,
            in2 => \N__24888\,
            in3 => \N__25024\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47424\,
            ce => \N__24468\,
            sr => \N__46924\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011101100"
        )
    port map (
            in0 => \N__25025\,
            in1 => \N__24850\,
            in2 => \N__21873\,
            in3 => \N__24661\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47424\,
            ce => \N__24468\,
            sr => \N__46924\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011101100"
        )
    port map (
            in0 => \N__25027\,
            in1 => \N__24851\,
            in2 => \N__21852\,
            in3 => \N__24663\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47424\,
            ce => \N__24468\,
            sr => \N__46924\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24234\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47424\,
            ce => \N__24468\,
            sr => \N__46924\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21753\,
            in2 => \N__20604\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            clk => \N__47416\,
            ce => \N__24502\,
            sr => \N__46927\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21729\,
            in2 => \N__20910\,
            in3 => \N__20880\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \N__47416\,
            ce => \N__24502\,
            sr => \N__46927\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20877\,
            in2 => \N__21702\,
            in3 => \N__20853\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__47416\,
            ce => \N__24502\,
            sr => \N__46927\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22533\,
            in2 => \N__22152\,
            in3 => \N__20814\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__47416\,
            ce => \N__24502\,
            sr => \N__46927\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22566\,
            in2 => \N__22881\,
            in3 => \N__20775\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__47416\,
            ce => \N__24502\,
            sr => \N__46927\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20772\,
            in2 => \N__22374\,
            in3 => \N__20733\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__47416\,
            ce => \N__24502\,
            sr => \N__46927\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22404\,
            in2 => \N__21909\,
            in3 => \N__20697\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__47416\,
            ce => \N__24502\,
            sr => \N__46927\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22433\,
            in2 => \N__20694\,
            in3 => \N__20643\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__47416\,
            ce => \N__24502\,
            sr => \N__46927\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22491\,
            in2 => \N__22128\,
            in3 => \N__20607\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__47408\,
            ce => \N__24507\,
            sr => \N__46931\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21606\,
            in2 => \N__22464\,
            in3 => \N__21033\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__47408\,
            ce => \N__24507\,
            sr => \N__46931\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22038\,
            in2 => \N__25077\,
            in3 => \N__21012\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__47408\,
            ce => \N__24507\,
            sr => \N__46931\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23145\,
            in2 => \N__22113\,
            in3 => \N__20997\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__47408\,
            ce => \N__24507\,
            sr => \N__46931\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22697\,
            in2 => \N__22023\,
            in3 => \N__20985\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__47408\,
            ce => \N__24507\,
            sr => \N__46931\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23226\,
            in2 => \N__22032\,
            in3 => \N__20967\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__47408\,
            ce => \N__24507\,
            sr => \N__46931\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23250\,
            in2 => \N__21921\,
            in3 => \N__20949\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__47408\,
            ce => \N__24507\,
            sr => \N__46931\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22617\,
            in2 => \N__22008\,
            in3 => \N__20928\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__47408\,
            ce => \N__24507\,
            sr => \N__46931\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21999\,
            in2 => \N__23190\,
            in3 => \N__20913\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_4_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__47399\,
            ce => \N__24508\,
            sr => \N__46936\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24540\,
            in2 => \N__21981\,
            in3 => \N__21198\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__47399\,
            ce => \N__24508\,
            sr => \N__46936\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23964\,
            in2 => \N__21993\,
            in3 => \N__21186\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__47399\,
            ce => \N__24508\,
            sr => \N__46936\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23106\,
            in2 => \N__22137\,
            in3 => \N__21174\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__47399\,
            ce => \N__24508\,
            sr => \N__46936\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23074\,
            in2 => \N__21960\,
            in3 => \N__21162\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__47399\,
            ce => \N__24508\,
            sr => \N__46936\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23822\,
            in2 => \N__25110\,
            in3 => \N__21147\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__47399\,
            ce => \N__24508\,
            sr => \N__46936\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23045\,
            in2 => \N__22101\,
            in3 => \N__21129\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__47399\,
            ce => \N__24508\,
            sr => \N__46936\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22083\,
            in2 => \N__22647\,
            in3 => \N__21108\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__47399\,
            ce => \N__24508\,
            sr => \N__46936\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23859\,
            in2 => \N__22092\,
            in3 => \N__21084\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_4_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__47389\,
            ce => \N__24509\,
            sr => \N__46940\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22917\,
            in2 => \N__23904\,
            in3 => \N__21066\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__47389\,
            ce => \N__24509\,
            sr => \N__46940\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22925\,
            in2 => \N__23787\,
            in3 => \N__21390\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__47389\,
            ce => \N__24509\,
            sr => \N__46940\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22856\,
            in2 => \N__22934\,
            in3 => \N__21369\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__47389\,
            ce => \N__24509\,
            sr => \N__46940\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22736\,
            in2 => \N__22932\,
            in3 => \N__21357\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__47389\,
            ce => \N__24509\,
            sr => \N__46940\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23292\,
            in2 => \N__22935\,
            in3 => \N__21333\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__47389\,
            ce => \N__24509\,
            sr => \N__46940\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22983\,
            in2 => \N__22933\,
            in3 => \N__21306\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__47389\,
            ce => \N__24509\,
            sr => \N__46940\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24867\,
            in1 => \N__22924\,
            in2 => \_gnd_net_\,
            in3 => \N__21303\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47389\,
            ce => \N__24509\,
            sr => \N__46940\
        );

    \counter_7_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__22314\,
            in1 => \N__22272\,
            in2 => \N__21228\,
            in3 => \N__22227\,
            lcout => \counterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47462\,
            ce => 'H',
            sr => \N__46848\
        );

    \counter_1_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21582\,
            in2 => \_gnd_net_\,
            in3 => \N__22072\,
            lcout => \counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47462\,
            ce => 'H',
            sr => \N__46848\
        );

    \counter_RNI800G_7_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21410\,
            in2 => \_gnd_net_\,
            in3 => \N__21218\,
            lcout => OPEN,
            ltout => \un2_counter_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI3BSP_1_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21593\,
            in1 => \N__21580\,
            in2 => \N__21564\,
            in3 => \N__22073\,
            lcout => un2_counter_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIM6001_12_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21560\,
            in1 => \N__21548\,
            in2 => \N__21435\,
            in3 => \N__21536\,
            lcout => un2_counter_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNII76D_3_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21524\,
            in1 => \N__21512\,
            in2 => \N__21501\,
            in3 => \N__21485\,
            lcout => un2_counter_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_4_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21474\,
            lcout => \pwm_generator_inst.thresholdZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47454\,
            ce => 'H',
            sr => \N__46867\
        );

    \pwm_generator_inst.threshold_2_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21462\,
            lcout => \pwm_generator_inst.thresholdZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47454\,
            ce => 'H',
            sr => \N__46867\
        );

    \pwm_generator_inst.threshold_6_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21456\,
            lcout => \pwm_generator_inst.thresholdZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47454\,
            ce => 'H',
            sr => \N__46867\
        );

    \counter_12_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__22313\,
            in1 => \N__22271\,
            in2 => \N__21444\,
            in3 => \N__22226\,
            lcout => \counterZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47454\,
            ce => 'H',
            sr => \N__46867\
        );

    \counter_10_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__22312\,
            in1 => \N__22270\,
            in2 => \N__21420\,
            in3 => \N__22225\,
            lcout => \counterZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47454\,
            ce => 'H',
            sr => \N__46867\
        );

    \pwm_generator_inst.threshold_8_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21636\,
            lcout => \pwm_generator_inst.thresholdZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47452\,
            ce => 'H',
            sr => \N__46877\
        );

    \pwm_generator_inst.threshold_3_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21627\,
            lcout => \pwm_generator_inst.thresholdZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47452\,
            ce => 'H',
            sr => \N__46877\
        );

    \pwm_generator_inst.threshold_7_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21621\,
            lcout => \pwm_generator_inst.thresholdZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47452\,
            ce => 'H',
            sr => \N__46877\
        );

    \pwm_generator_inst.threshold_5_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21612\,
            lcout => \pwm_generator_inst.thresholdZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47452\,
            ce => 'H',
            sr => \N__46877\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25224\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47449\,
            ce => \N__24407\,
            sr => \N__46886\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011010000"
        )
    port map (
            in0 => \N__24605\,
            in1 => \N__21894\,
            in2 => \N__24897\,
            in3 => \N__25005\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47441\,
            ce => \N__24475\,
            sr => \N__46894\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011010000"
        )
    port map (
            in0 => \N__24604\,
            in1 => \N__21765\,
            in2 => \N__24896\,
            in3 => \N__25004\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47441\,
            ce => \N__24475\,
            sr => \N__46894\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011010000"
        )
    port map (
            in0 => \N__24601\,
            in1 => \N__21810\,
            in2 => \N__24894\,
            in3 => \N__25001\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47441\,
            ce => \N__24475\,
            sr => \N__46894\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011010000"
        )
    port map (
            in0 => \N__24602\,
            in1 => \N__21798\,
            in2 => \N__24895\,
            in3 => \N__25002\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47441\,
            ce => \N__24475\,
            sr => \N__46894\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011101100"
        )
    port map (
            in0 => \N__25003\,
            in1 => \N__24872\,
            in2 => \N__21786\,
            in3 => \N__24603\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47441\,
            ce => \N__24475\,
            sr => \N__46894\
        );

    \current_shift_inst.PI_CTRL.integrator_0_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21746\,
            in2 => \N__24281\,
            in3 => \N__22802\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\,
            clk => \N__47432\,
            ce => \N__24484\,
            sr => \N__46907\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__22800\,
            in1 => \N__21722\,
            in2 => \N__24258\,
            in3 => \N__21705\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \N__47432\,
            ce => \N__24484\,
            sr => \N__46907\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__22803\,
            in1 => \N__21697\,
            in2 => \N__24233\,
            in3 => \N__21678\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \N__47432\,
            ce => \N__24484\,
            sr => \N__46907\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__22801\,
            in1 => \N__22527\,
            in2 => \N__24207\,
            in3 => \N__21675\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \N__47432\,
            ce => \N__24484\,
            sr => \N__46907\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22560\,
            in2 => \N__25368\,
            in3 => \N__21666\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22357\,
            in2 => \N__25343\,
            in3 => \N__21657\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22398\,
            in2 => \N__25311\,
            in3 => \N__21648\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22425\,
            in2 => \N__25283\,
            in3 => \N__21639\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22485\,
            in2 => \N__25254\,
            in3 => \N__21828\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22455\,
            in2 => \N__25223\,
            in3 => \N__21816\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25191\,
            in2 => \N__25076\,
            in3 => \N__21813\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25166\,
            in2 => \N__23144\,
            in3 => \N__21801\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25595\,
            in2 => \N__22696\,
            in3 => \N__21789\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23220\,
            in2 => \N__25575\,
            in3 => \N__21774\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23257\,
            in2 => \N__25551\,
            in3 => \N__21771\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22613\,
            in2 => \N__25527\,
            in3 => \N__21768\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23175\,
            in2 => \N__25503\,
            in3 => \N__21756\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24536\,
            in2 => \N__25476\,
            in3 => \N__21897\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23944\,
            in2 => \N__25449\,
            in3 => \N__21885\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23100\,
            in2 => \N__25419\,
            in3 => \N__21876\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23073\,
            in2 => \N__25392\,
            in3 => \N__21864\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23808\,
            in2 => \N__25737\,
            in3 => \N__21855\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23037\,
            in2 => \N__25710\,
            in3 => \N__21843\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22643\,
            in2 => \N__25683\,
            in3 => \N__21840\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23855\,
            in2 => \N__25656\,
            in3 => \N__21837\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27221\,
            in2 => \N__23898\,
            in3 => \N__21951\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23779\,
            in2 => \N__27237\,
            in3 => \N__21948\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27225\,
            in2 => \N__22857\,
            in3 => \N__21945\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22735\,
            in2 => \N__27238\,
            in3 => \N__21933\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23288\,
            in2 => \N__27243\,
            in3 => \N__21930\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22978\,
            in2 => \N__27239\,
            in3 => \N__21927\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24782\,
            in1 => \N__27232\,
            in2 => \_gnd_net_\,
            in3 => \N__21924\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25550\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47400\,
            ce => \N__24506\,
            sr => \N__46928\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25310\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47400\,
            ce => \N__24506\,
            sr => \N__46928\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25190\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47400\,
            ce => \N__24506\,
            sr => \N__46928\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25574\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47400\,
            ce => \N__24506\,
            sr => \N__46928\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25596\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47400\,
            ce => \N__24506\,
            sr => \N__46928\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__22014\,
            in1 => \N__24671\,
            in2 => \N__24871\,
            in3 => \N__25034\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47400\,
            ce => \N__24506\,
            sr => \N__46928\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25526\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47400\,
            ce => \N__24506\,
            sr => \N__46928\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25499\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47390\,
            ce => \N__24499\,
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25442\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47390\,
            ce => \N__24499\,
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25472\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47390\,
            ce => \N__24499\,
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__21969\,
            in1 => \N__24672\,
            in2 => \N__24893\,
            in3 => \N__25035\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47390\,
            ce => \N__24499\,
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25388\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47390\,
            ce => \N__24499\,
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24206\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47390\,
            ce => \N__24499\,
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25415\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47390\,
            ce => \N__24499\,
            sr => \N__46932\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25253\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47381\,
            ce => \N__24501\,
            sr => \N__46937\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25167\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47381\,
            ce => \N__24501\,
            sr => \N__46937\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25709\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47381\,
            ce => \N__24501\,
            sr => \N__46937\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25652\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47381\,
            ce => \N__24501\,
            sr => \N__46937\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25682\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47381\,
            ce => \N__24501\,
            sr => \N__46937\
        );

    \counter_0_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__22236\,
            in1 => \N__22329\,
            in2 => \N__22071\,
            in3 => \N__22283\,
            lcout => \counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47455\,
            ce => 'H',
            sr => \N__46836\
        );

    \clk_10khz_RNIIENA2_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__22321\,
            in1 => \N__22273\,
            in2 => \N__22194\,
            in3 => \N__22228\,
            lcout => \clk_10khz_RNIIENAZ0Z2\,
            ltout => \clk_10khz_RNIIENAZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__35047\,
            in1 => \_gnd_net_\,
            in2 => \N__22338\,
            in3 => \N__22191\,
            lcout => \N_655_g\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.phase_valid_RNISLOR2_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__28998\,
            in1 => \N__22192\,
            in2 => \N__35059\,
            in3 => \N__22335\,
            lcout => \current_shift_inst.phase_valid_RNISLORZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_10khz_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__22328\,
            in1 => \N__22193\,
            in2 => \N__22284\,
            in3 => \N__22235\,
            lcout => clk_10khz_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47450\,
            ce => 'H',
            sr => \N__46849\
        );

    \pwm_generator_inst.threshold_1_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22173\,
            lcout => \pwm_generator_inst.thresholdZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47442\,
            ce => 'H',
            sr => \N__46857\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23605\,
            in2 => \_gnd_net_\,
            in3 => \N__23653\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__24178\,
            in1 => \N__23584\,
            in2 => \N__22164\,
            in3 => \N__23632\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__22158\,
            in1 => \N__24131\,
            in2 => \N__22161\,
            in3 => \N__24155\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__24079\,
            in1 => \N__24010\,
            in2 => \_gnd_net_\,
            in3 => \N__24106\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22779\,
            in1 => \N__22584\,
            in2 => \N__22770\,
            in3 => \N__22656\,
            lcout => \current_shift_inst.PI_CTRL.N_46_21\,
            ltout => \current_shift_inst.PI_CTRL.N_46_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23016\,
            in1 => \N__23961\,
            in2 => \N__22587\,
            in3 => \N__22500\,
            lcout => \current_shift_inst.PI_CTRL.N_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23262\,
            in1 => \N__23224\,
            in2 => \N__23188\,
            in3 => \N__23142\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFCK44_4_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__22565\,
            in1 => \N__22578\,
            in2 => \_gnd_net_\,
            in3 => \N__22344\,
            lcout => \current_shift_inst.PI_CTRL.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22457\,
            in1 => \N__22402\,
            in2 => \N__22434\,
            in3 => \N__22367\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__22490\,
            in1 => \N__22564\,
            in2 => \N__22536\,
            in3 => \N__22529\,
            lcout => \current_shift_inst.PI_CTRL.N_44\,
            ltout => \current_shift_inst.PI_CTRL.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24823\,
            in1 => \N__23951\,
            in2 => \N__22494\,
            in3 => \N__23015\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__22489\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22456\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__22432\,
            in1 => \N__22403\,
            in2 => \N__22377\,
            in3 => \N__22366\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__23993\,
            in1 => \N__24824\,
            in2 => \N__23962\,
            in3 => \N__25121\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__22818\,
            in1 => \N__22812\,
            in2 => \N__22806\,
            in3 => \N__23975\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22734\,
            in1 => \N__22846\,
            in2 => \N__22982\,
            in3 => \N__22698\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23902\,
            in1 => \N__23854\,
            in2 => \N__23783\,
            in3 => \N__23818\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__22758\,
            in1 => \N__24641\,
            in2 => \N__24828\,
            in3 => \N__24949\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47409\,
            ce => \N__24411\,
            sr => \N__46895\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000001100"
        )
    port map (
            in0 => \N__24950\,
            in1 => \N__24778\,
            in2 => \N__24670\,
            in3 => \N__22749\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47409\,
            ce => \N__24411\,
            sr => \N__46895\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22737\,
            in1 => \N__22842\,
            in2 => \N__22974\,
            in3 => \N__22695\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25056\,
            in1 => \N__23280\,
            in2 => \N__22612\,
            in3 => \N__22631\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22630\,
            in1 => \N__22602\,
            in2 => \N__23287\,
            in3 => \N__25057\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23258\,
            in1 => \N__23225\,
            in2 => \N__23189\,
            in3 => \N__23143\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24535\,
            in1 => \N__23044\,
            in2 => \N__23079\,
            in3 => \N__23105\,
            lcout => \current_shift_inst.PI_CTRL.N_47_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23104\,
            in1 => \N__23075\,
            in2 => \N__23046\,
            in3 => \N__24534\,
            lcout => \current_shift_inst.PI_CTRL.N_46_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011000100"
        )
    port map (
            in0 => \N__24649\,
            in1 => \N__24752\,
            in2 => \N__22998\,
            in3 => \N__24975\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47391\,
            ce => \N__24476\,
            sr => \N__46913\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__24972\,
            in1 => \N__22944\,
            in2 => \N__24819\,
            in3 => \N__24646\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47391\,
            ce => \N__24476\,
            sr => \N__46913\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27233\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47391\,
            ce => \N__24476\,
            sr => \N__46913\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__24971\,
            in1 => \N__22890\,
            in2 => \N__24818\,
            in3 => \N__24645\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47391\,
            ce => \N__24476\,
            sr => \N__46913\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25361\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47391\,
            ce => \N__24476\,
            sr => \N__46913\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__24973\,
            in1 => \N__22866\,
            in2 => \N__24820\,
            in3 => \N__24647\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47391\,
            ce => \N__24476\,
            sr => \N__46913\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011000100"
        )
    port map (
            in0 => \N__24650\,
            in1 => \N__24753\,
            in2 => \N__23316\,
            in3 => \N__24976\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47391\,
            ce => \N__24476\,
            sr => \N__46913\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__24974\,
            in1 => \N__23301\,
            in2 => \N__24821\,
            in3 => \N__24648\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47391\,
            ce => \N__24476\,
            sr => \N__46913\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__28048\,
            in1 => \N__28414\,
            in2 => \N__29529\,
            in3 => \N__29482\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27304\,
            in2 => \_gnd_net_\,
            in3 => \N__29635\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29605\,
            in2 => \_gnd_net_\,
            in3 => \N__28262\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNILORI_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__27336\,
            in1 => \N__27305\,
            in2 => \N__29673\,
            in3 => \N__29636\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29668\,
            in2 => \_gnd_net_\,
            in3 => \N__27335\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__28261\,
            in1 => \N__29637\,
            in2 => \N__29607\,
            in3 => \N__27306\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__27334\,
            in1 => \N__28159\,
            in2 => \N__29718\,
            in3 => \N__29672\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \N__29832\,
            in1 => \N__27408\,
            in2 => \N__27381\,
            in3 => \N__29801\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIDR081_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27406\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29831\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27379\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29800\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__27407\,
            in1 => \N__27437\,
            in2 => \N__29865\,
            in3 => \N__29830\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPC571_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27438\,
            in3 => \N__29860\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__27380\,
            in1 => \N__30346\,
            in2 => \N__29805\,
            in3 => \N__30289\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__30290\,
            in1 => \_gnd_net_\,
            in2 => \N__30351\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIR32K_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__29861\,
            in1 => \N__27471\,
            in2 => \N__29907\,
            in3 => \N__27433\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIE6961_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__27466\,
            in1 => \N__29902\,
            in2 => \N__29949\,
            in3 => \N__28345\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIH6661_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__29903\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27467\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111000011"
        )
    port map (
            in0 => \N__30402\,
            in1 => \N__27940\,
            in2 => \N__30203\,
            in3 => \N__30441\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27945\,
            in3 => \N__30196\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__27913\,
            in1 => \N__27944\,
            in2 => \N__30204\,
            in3 => \N__30166\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINKG81_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__30167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27914\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111000011"
        )
    port map (
            in0 => \N__27915\,
            in1 => \N__30137\,
            in2 => \N__27888\,
            in3 => \N__30168\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__30138\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27887\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__26969\,
            in1 => \N__30524\,
            in2 => \_gnd_net_\,
            in3 => \N__30477\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.counter_0_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26585\,
            in1 => \N__28648\,
            in2 => \_gnd_net_\,
            in3 => \N__23325\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_0\,
            clk => \N__47345\,
            ce => \N__33641\,
            sr => \N__46941\
        );

    \current_shift_inst.timer_phase.counter_1_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26580\,
            in1 => \N__28687\,
            in2 => \_gnd_net_\,
            in3 => \N__23322\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_0\,
            carryout => \current_shift_inst.timer_phase.counter_cry_1\,
            clk => \N__47345\,
            ce => \N__33641\,
            sr => \N__46941\
        );

    \current_shift_inst.timer_phase.counter_2_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26586\,
            in1 => \N__25615\,
            in2 => \_gnd_net_\,
            in3 => \N__23319\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_1\,
            carryout => \current_shift_inst.timer_phase.counter_cry_2\,
            clk => \N__47345\,
            ce => \N__33641\,
            sr => \N__46941\
        );

    \current_shift_inst.timer_phase.counter_3_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26581\,
            in1 => \N__25975\,
            in2 => \_gnd_net_\,
            in3 => \N__23352\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_2\,
            carryout => \current_shift_inst.timer_phase.counter_cry_3\,
            clk => \N__47345\,
            ce => \N__33641\,
            sr => \N__46941\
        );

    \current_shift_inst.timer_phase.counter_4_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26587\,
            in1 => \N__25949\,
            in2 => \_gnd_net_\,
            in3 => \N__23349\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_3\,
            carryout => \current_shift_inst.timer_phase.counter_cry_4\,
            clk => \N__47345\,
            ce => \N__33641\,
            sr => \N__46941\
        );

    \current_shift_inst.timer_phase.counter_5_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26582\,
            in1 => \N__25930\,
            in2 => \_gnd_net_\,
            in3 => \N__23346\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_4\,
            carryout => \current_shift_inst.timer_phase.counter_cry_5\,
            clk => \N__47345\,
            ce => \N__33641\,
            sr => \N__46941\
        );

    \current_shift_inst.timer_phase.counter_6_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26584\,
            in1 => \N__25898\,
            in2 => \_gnd_net_\,
            in3 => \N__23343\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_5\,
            carryout => \current_shift_inst.timer_phase.counter_cry_6\,
            clk => \N__47345\,
            ce => \N__33641\,
            sr => \N__46941\
        );

    \current_shift_inst.timer_phase.counter_7_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26583\,
            in1 => \N__25868\,
            in2 => \_gnd_net_\,
            in3 => \N__23340\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_6\,
            carryout => \current_shift_inst.timer_phase.counter_cry_7\,
            clk => \N__47345\,
            ce => \N__33641\,
            sr => \N__46941\
        );

    \current_shift_inst.timer_phase.counter_8_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26591\,
            in1 => \N__25843\,
            in2 => \_gnd_net_\,
            in3 => \N__23337\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_20_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_8\,
            clk => \N__47337\,
            ce => \N__33645\,
            sr => \N__46943\
        );

    \current_shift_inst.timer_phase.counter_9_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26595\,
            in1 => \N__25813\,
            in2 => \_gnd_net_\,
            in3 => \N__23334\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_8\,
            carryout => \current_shift_inst.timer_phase.counter_cry_9\,
            clk => \N__47337\,
            ce => \N__33645\,
            sr => \N__46943\
        );

    \current_shift_inst.timer_phase.counter_10_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26588\,
            in1 => \N__25783\,
            in2 => \_gnd_net_\,
            in3 => \N__23331\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_9\,
            carryout => \current_shift_inst.timer_phase.counter_cry_10\,
            clk => \N__47337\,
            ce => \N__33645\,
            sr => \N__46943\
        );

    \current_shift_inst.timer_phase.counter_11_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26592\,
            in1 => \N__25756\,
            in2 => \_gnd_net_\,
            in3 => \N__23328\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_10\,
            carryout => \current_shift_inst.timer_phase.counter_cry_11\,
            clk => \N__47337\,
            ce => \N__33645\,
            sr => \N__46943\
        );

    \current_shift_inst.timer_phase.counter_12_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26589\,
            in1 => \N__26182\,
            in2 => \_gnd_net_\,
            in3 => \N__23379\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_11\,
            carryout => \current_shift_inst.timer_phase.counter_cry_12\,
            clk => \N__47337\,
            ce => \N__33645\,
            sr => \N__46943\
        );

    \current_shift_inst.timer_phase.counter_13_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26593\,
            in1 => \N__26152\,
            in2 => \_gnd_net_\,
            in3 => \N__23376\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_12\,
            carryout => \current_shift_inst.timer_phase.counter_cry_13\,
            clk => \N__47337\,
            ce => \N__33645\,
            sr => \N__46943\
        );

    \current_shift_inst.timer_phase.counter_14_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26590\,
            in1 => \N__26131\,
            in2 => \_gnd_net_\,
            in3 => \N__23373\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_13\,
            carryout => \current_shift_inst.timer_phase.counter_cry_14\,
            clk => \N__47337\,
            ce => \N__33645\,
            sr => \N__46943\
        );

    \current_shift_inst.timer_phase.counter_15_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26594\,
            in1 => \N__26110\,
            in2 => \_gnd_net_\,
            in3 => \N__23370\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_14\,
            carryout => \current_shift_inst.timer_phase.counter_cry_15\,
            clk => \N__47337\,
            ce => \N__33645\,
            sr => \N__46943\
        );

    \current_shift_inst.timer_phase.counter_16_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26536\,
            in1 => \N__26086\,
            in2 => \_gnd_net_\,
            in3 => \N__23367\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_7_21_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_16\,
            clk => \N__47331\,
            ce => \N__33640\,
            sr => \N__46944\
        );

    \current_shift_inst.timer_phase.counter_17_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26540\,
            in1 => \N__26059\,
            in2 => \_gnd_net_\,
            in3 => \N__23364\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_16\,
            carryout => \current_shift_inst.timer_phase.counter_cry_17\,
            clk => \N__47331\,
            ce => \N__33640\,
            sr => \N__46944\
        );

    \current_shift_inst.timer_phase.counter_18_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26537\,
            in1 => \N__26029\,
            in2 => \_gnd_net_\,
            in3 => \N__23361\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_17\,
            carryout => \current_shift_inst.timer_phase.counter_cry_18\,
            clk => \N__47331\,
            ce => \N__33640\,
            sr => \N__46944\
        );

    \current_shift_inst.timer_phase.counter_19_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26541\,
            in1 => \N__26002\,
            in2 => \_gnd_net_\,
            in3 => \N__23358\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_18\,
            carryout => \current_shift_inst.timer_phase.counter_cry_19\,
            clk => \N__47331\,
            ce => \N__33640\,
            sr => \N__46944\
        );

    \current_shift_inst.timer_phase.counter_20_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26538\,
            in1 => \N__26428\,
            in2 => \_gnd_net_\,
            in3 => \N__23355\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_19\,
            carryout => \current_shift_inst.timer_phase.counter_cry_20\,
            clk => \N__47331\,
            ce => \N__33640\,
            sr => \N__46944\
        );

    \current_shift_inst.timer_phase.counter_21_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26542\,
            in1 => \N__26398\,
            in2 => \_gnd_net_\,
            in3 => \N__23418\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_20\,
            carryout => \current_shift_inst.timer_phase.counter_cry_21\,
            clk => \N__47331\,
            ce => \N__33640\,
            sr => \N__46944\
        );

    \current_shift_inst.timer_phase.counter_22_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26539\,
            in1 => \N__26377\,
            in2 => \_gnd_net_\,
            in3 => \N__23415\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_21\,
            carryout => \current_shift_inst.timer_phase.counter_cry_22\,
            clk => \N__47331\,
            ce => \N__33640\,
            sr => \N__46944\
        );

    \current_shift_inst.timer_phase.counter_23_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26543\,
            in1 => \N__26356\,
            in2 => \_gnd_net_\,
            in3 => \N__23412\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_22\,
            carryout => \current_shift_inst.timer_phase.counter_cry_23\,
            clk => \N__47331\,
            ce => \N__33640\,
            sr => \N__46944\
        );

    \current_shift_inst.timer_phase.counter_24_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26530\,
            in1 => \N__26332\,
            in2 => \_gnd_net_\,
            in3 => \N__23409\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_7_22_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_24\,
            clk => \N__47326\,
            ce => \N__33639\,
            sr => \N__46946\
        );

    \current_shift_inst.timer_phase.counter_25_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26534\,
            in1 => \N__26305\,
            in2 => \_gnd_net_\,
            in3 => \N__23406\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_24\,
            carryout => \current_shift_inst.timer_phase.counter_cry_25\,
            clk => \N__47326\,
            ce => \N__33639\,
            sr => \N__46946\
        );

    \current_shift_inst.timer_phase.counter_26_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26531\,
            in1 => \N__26257\,
            in2 => \_gnd_net_\,
            in3 => \N__23403\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_25\,
            carryout => \current_shift_inst.timer_phase.counter_cry_26\,
            clk => \N__47326\,
            ce => \N__33639\,
            sr => \N__46946\
        );

    \current_shift_inst.timer_phase.counter_27_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26535\,
            in1 => \N__26212\,
            in2 => \_gnd_net_\,
            in3 => \N__23400\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_26\,
            carryout => \current_shift_inst.timer_phase.counter_cry_27\,
            clk => \N__47326\,
            ce => \N__33639\,
            sr => \N__46946\
        );

    \current_shift_inst.timer_phase.counter_28_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26532\,
            in1 => \N__26279\,
            in2 => \_gnd_net_\,
            in3 => \N__23397\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_27\,
            carryout => \current_shift_inst.timer_phase.counter_cry_28\,
            clk => \N__47326\,
            ce => \N__33639\,
            sr => \N__46946\
        );

    \current_shift_inst.timer_phase.counter_29_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__26234\,
            in1 => \N__26533\,
            in2 => \_gnd_net_\,
            in3 => \N__23394\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47326\,
            ce => \N__33639\,
            sr => \N__46946\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23391\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47456\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23562\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47456\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23535\,
            in2 => \N__23553\,
            in3 => \N__23658\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23520\,
            in2 => \N__23529\,
            in3 => \N__23634\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23502\,
            in2 => \N__23514\,
            in3 => \N__23610\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23496\,
            in2 => \N__23484\,
            in3 => \N__23586\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23463\,
            in2 => \N__23475\,
            in3 => \N__24180\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24156\,
            in1 => \N__23442\,
            in2 => \N__23457\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23424\,
            in2 => \N__23436\,
            in3 => \N__24132\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24108\,
            in1 => \N__23745\,
            in2 => \N__23733\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23712\,
            in2 => \N__23724\,
            in3 => \N__24084\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23691\,
            in2 => \N__23706\,
            in3 => \N__24015\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23685\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47433\,
            ce => 'H',
            sr => \N__46850\
        );

    \pwm_generator_inst.counter_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24057\,
            in1 => \N__23657\,
            in2 => \_gnd_net_\,
            in3 => \N__23637\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__47425\,
            ce => 'H',
            sr => \N__46858\
        );

    \pwm_generator_inst.counter_1_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24042\,
            in1 => \N__23633\,
            in2 => \_gnd_net_\,
            in3 => \N__23613\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__47425\,
            ce => 'H',
            sr => \N__46858\
        );

    \pwm_generator_inst.counter_2_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24058\,
            in1 => \N__23609\,
            in2 => \_gnd_net_\,
            in3 => \N__23589\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__47425\,
            ce => 'H',
            sr => \N__46858\
        );

    \pwm_generator_inst.counter_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24043\,
            in1 => \N__23585\,
            in2 => \_gnd_net_\,
            in3 => \N__23565\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__47425\,
            ce => 'H',
            sr => \N__46858\
        );

    \pwm_generator_inst.counter_4_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24059\,
            in1 => \N__24179\,
            in2 => \_gnd_net_\,
            in3 => \N__24159\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__47425\,
            ce => 'H',
            sr => \N__46858\
        );

    \pwm_generator_inst.counter_5_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24044\,
            in1 => \N__24154\,
            in2 => \_gnd_net_\,
            in3 => \N__24135\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__47425\,
            ce => 'H',
            sr => \N__46858\
        );

    \pwm_generator_inst.counter_6_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24060\,
            in1 => \N__24130\,
            in2 => \_gnd_net_\,
            in3 => \N__24111\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__47425\,
            ce => 'H',
            sr => \N__46858\
        );

    \pwm_generator_inst.counter_7_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24045\,
            in1 => \N__24107\,
            in2 => \_gnd_net_\,
            in3 => \N__24087\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__47425\,
            ce => 'H',
            sr => \N__46858\
        );

    \pwm_generator_inst.counter_8_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24047\,
            in1 => \N__24083\,
            in2 => \_gnd_net_\,
            in3 => \N__24063\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__47417\,
            ce => 'H',
            sr => \N__46868\
        );

    \pwm_generator_inst.counter_9_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__24014\,
            in1 => \N__24046\,
            in2 => \_gnd_net_\,
            in3 => \N__24018\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47417\,
            ce => 'H',
            sr => \N__46868\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23994\,
            in1 => \N__23976\,
            in2 => \N__23963\,
            in3 => \N__25122\,
            lcout => \current_shift_inst.PI_CTRL.N_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23903\,
            in1 => \N__23853\,
            in2 => \N__23823\,
            in3 => \N__23775\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25143\,
            in1 => \N__25137\,
            in2 => \N__25131\,
            in3 => \N__25128\,
            lcout => \current_shift_inst.PI_CTRL.N_47_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25733\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47392\,
            ce => \N__24467\,
            sr => \N__46896\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011000100"
        )
    port map (
            in0 => \N__24651\,
            in1 => \N__24766\,
            in2 => \N__25092\,
            in3 => \N__24969\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47392\,
            ce => \N__24467\,
            sr => \N__46896\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__24970\,
            in1 => \N__24906\,
            in2 => \N__24822\,
            in3 => \N__24652\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47392\,
            ce => \N__24467\,
            sr => \N__46896\
        );

    \current_shift_inst.control_input_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26613\,
            in2 => \N__30708\,
            in3 => \N__30707\,
            lcout => \current_shift_inst.control_inputZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \current_shift_inst.control_input_1_cry_0\,
            clk => \N__47382\,
            ce => \N__27162\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26604\,
            in2 => \_gnd_net_\,
            in3 => \N__24237\,
            lcout => \current_shift_inst.control_inputZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_0\,
            carryout => \current_shift_inst.control_input_1_cry_1\,
            clk => \N__47382\,
            ce => \N__27162\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26772\,
            in2 => \_gnd_net_\,
            in3 => \N__24210\,
            lcout => \current_shift_inst.control_inputZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_1\,
            carryout => \current_shift_inst.control_input_1_cry_2\,
            clk => \N__47382\,
            ce => \N__27162\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_3_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26754\,
            in2 => \_gnd_net_\,
            in3 => \N__24183\,
            lcout => \current_shift_inst.control_inputZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_2\,
            carryout => \current_shift_inst.control_input_1_cry_3\,
            clk => \N__47382\,
            ce => \N__27162\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_4_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26721\,
            in2 => \_gnd_net_\,
            in3 => \N__25347\,
            lcout => \current_shift_inst.control_inputZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_3\,
            carryout => \current_shift_inst.control_input_1_cry_4\,
            clk => \N__47382\,
            ce => \N__27162\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_5_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26688\,
            in2 => \_gnd_net_\,
            in3 => \N__25314\,
            lcout => \current_shift_inst.control_inputZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_4\,
            carryout => \current_shift_inst.control_input_1_cry_5\,
            clk => \N__47382\,
            ce => \N__27162\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_6_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26667\,
            in2 => \_gnd_net_\,
            in3 => \N__25287\,
            lcout => \current_shift_inst.control_inputZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_5\,
            carryout => \current_shift_inst.control_input_1_cry_6\,
            clk => \N__47382\,
            ce => \N__27162\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_7_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26658\,
            in2 => \_gnd_net_\,
            in3 => \N__25257\,
            lcout => \current_shift_inst.control_inputZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_6\,
            carryout => \current_shift_inst.control_input_1_cry_7\,
            clk => \N__47382\,
            ce => \N__27162\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_8_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26637\,
            in2 => \_gnd_net_\,
            in3 => \N__25227\,
            lcout => \current_shift_inst.control_inputZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \current_shift_inst.control_input_1_cry_8\,
            clk => \N__47376\,
            ce => \N__27174\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_9_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26946\,
            in2 => \_gnd_net_\,
            in3 => \N__25194\,
            lcout => \current_shift_inst.control_inputZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_8\,
            carryout => \current_shift_inst.control_input_1_cry_9\,
            clk => \N__47376\,
            ce => \N__27174\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_10_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26937\,
            in2 => \_gnd_net_\,
            in3 => \N__25170\,
            lcout => \current_shift_inst.control_inputZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_9\,
            carryout => \current_shift_inst.control_input_1_cry_10\,
            clk => \N__47376\,
            ce => \N__27174\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_11_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26928\,
            in2 => \_gnd_net_\,
            in3 => \N__25146\,
            lcout => \current_shift_inst.control_inputZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_10\,
            carryout => \current_shift_inst.control_input_1_cry_11\,
            clk => \N__47376\,
            ce => \N__27174\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_12_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26907\,
            in2 => \_gnd_net_\,
            in3 => \N__25578\,
            lcout => \current_shift_inst.control_inputZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_11\,
            carryout => \current_shift_inst.control_input_1_cry_12\,
            clk => \N__47376\,
            ce => \N__27174\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_13_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26874\,
            in2 => \_gnd_net_\,
            in3 => \N__25554\,
            lcout => \current_shift_inst.control_inputZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_12\,
            carryout => \current_shift_inst.control_input_1_cry_13\,
            clk => \N__47376\,
            ce => \N__27174\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_14_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26844\,
            in2 => \_gnd_net_\,
            in3 => \N__25530\,
            lcout => \current_shift_inst.control_inputZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_13\,
            carryout => \current_shift_inst.control_input_1_cry_14\,
            clk => \N__47376\,
            ce => \N__27174\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_15_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26814\,
            in2 => \_gnd_net_\,
            in3 => \N__25506\,
            lcout => \current_shift_inst.control_inputZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_14\,
            carryout => \current_shift_inst.control_input_1_cry_15\,
            clk => \N__47376\,
            ce => \N__27174\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_16_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26784\,
            in2 => \_gnd_net_\,
            in3 => \N__25479\,
            lcout => \current_shift_inst.control_inputZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \current_shift_inst.control_input_1_cry_16\,
            clk => \N__47369\,
            ce => \N__27184\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_17_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27099\,
            in2 => \_gnd_net_\,
            in3 => \N__25452\,
            lcout => \current_shift_inst.control_inputZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_16\,
            carryout => \current_shift_inst.control_input_1_cry_17\,
            clk => \N__47369\,
            ce => \N__27184\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_18_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27090\,
            in2 => \_gnd_net_\,
            in3 => \N__25422\,
            lcout => \current_shift_inst.control_inputZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_17\,
            carryout => \current_shift_inst.control_input_1_cry_18\,
            clk => \N__47369\,
            ce => \N__27184\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_19_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27081\,
            in2 => \_gnd_net_\,
            in3 => \N__25395\,
            lcout => \current_shift_inst.control_inputZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_18\,
            carryout => \current_shift_inst.control_input_1_cry_19\,
            clk => \N__47369\,
            ce => \N__27184\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_20_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27072\,
            in2 => \_gnd_net_\,
            in3 => \N__25371\,
            lcout => \current_shift_inst.control_inputZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_19\,
            carryout => \current_shift_inst.control_input_1_cry_20\,
            clk => \N__47369\,
            ce => \N__27184\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_21_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27054\,
            in2 => \_gnd_net_\,
            in3 => \N__25713\,
            lcout => \current_shift_inst.control_inputZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_20\,
            carryout => \current_shift_inst.control_input_1_cry_21\,
            clk => \N__47369\,
            ce => \N__27184\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_22_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27024\,
            in2 => \_gnd_net_\,
            in3 => \N__25686\,
            lcout => \current_shift_inst.control_inputZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_21\,
            carryout => \current_shift_inst.control_input_1_cry_22\,
            clk => \N__47369\,
            ce => \N__27184\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_23_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26994\,
            in2 => \_gnd_net_\,
            in3 => \N__25659\,
            lcout => \current_shift_inst.control_inputZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_22\,
            carryout => \current_shift_inst.control_input_1_cry_23\,
            clk => \N__47369\,
            ce => \N__27184\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_24_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26955\,
            in2 => \_gnd_net_\,
            in3 => \N__25632\,
            lcout => \current_shift_inst.control_inputZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \current_shift_inst.control_input_1_cry_24\,
            clk => \N__47362\,
            ce => \N__27186\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25629\,
            lcout => \current_shift_inst.control_input_1_cry_24_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28655\,
            in2 => \N__25622\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_3\,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\,
            clk => \N__47355\,
            ce => \N__28632\,
            sr => \N__46929\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28700\,
            in2 => \N__25982\,
            in3 => \N__25626\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\,
            clk => \N__47355\,
            ce => \N__28632\,
            sr => \N__46929\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25955\,
            in2 => \N__25623\,
            in3 => \N__25599\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\,
            clk => \N__47355\,
            ce => \N__28632\,
            sr => \N__46929\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25931\,
            in2 => \N__25983\,
            in3 => \N__25959\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\,
            clk => \N__47355\,
            ce => \N__28632\,
            sr => \N__46929\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25956\,
            in2 => \N__25910\,
            in3 => \N__25935\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\,
            clk => \N__47355\,
            ce => \N__28632\,
            sr => \N__46929\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25932\,
            in2 => \N__25880\,
            in3 => \N__25914\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\,
            clk => \N__47355\,
            ce => \N__28632\,
            sr => \N__46929\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25851\,
            in2 => \N__25911\,
            in3 => \N__25884\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\,
            clk => \N__47355\,
            ce => \N__28632\,
            sr => \N__46929\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25821\,
            in2 => \N__25881\,
            in3 => \N__25854\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9\,
            clk => \N__47355\,
            ce => \N__28632\,
            sr => \N__46929\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25850\,
            in2 => \N__25790\,
            in3 => \N__25824\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_11\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\,
            clk => \N__47346\,
            ce => \N__28631\,
            sr => \N__46933\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25820\,
            in2 => \N__25763\,
            in3 => \N__25794\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\,
            clk => \N__47346\,
            ce => \N__28631\,
            sr => \N__46933\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26189\,
            in2 => \N__25791\,
            in3 => \N__25767\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\,
            clk => \N__47346\,
            ce => \N__28631\,
            sr => \N__46933\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26159\,
            in2 => \N__25764\,
            in3 => \N__25740\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\,
            clk => \N__47346\,
            ce => \N__28631\,
            sr => \N__46933\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26132\,
            in2 => \N__26193\,
            in3 => \N__26166\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\,
            clk => \N__47346\,
            ce => \N__28631\,
            sr => \N__46933\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26111\,
            in2 => \N__26163\,
            in3 => \N__26136\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\,
            clk => \N__47346\,
            ce => \N__28631\,
            sr => \N__46933\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26133\,
            in2 => \N__26091\,
            in3 => \N__26115\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\,
            clk => \N__47346\,
            ce => \N__28631\,
            sr => \N__46933\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26112\,
            in2 => \N__26064\,
            in3 => \N__26094\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17\,
            clk => \N__47346\,
            ce => \N__28631\,
            sr => \N__46933\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26090\,
            in2 => \N__26036\,
            in3 => \N__26067\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_19\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\,
            clk => \N__47338\,
            ce => \N__28629\,
            sr => \N__46938\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26063\,
            in2 => \N__26009\,
            in3 => \N__26040\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\,
            clk => \N__47338\,
            ce => \N__28629\,
            sr => \N__46938\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26435\,
            in2 => \N__26037\,
            in3 => \N__26013\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\,
            clk => \N__47338\,
            ce => \N__28629\,
            sr => \N__46938\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26405\,
            in2 => \N__26010\,
            in3 => \N__25986\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\,
            clk => \N__47338\,
            ce => \N__28629\,
            sr => \N__46938\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26378\,
            in2 => \N__26439\,
            in3 => \N__26412\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\,
            clk => \N__47338\,
            ce => \N__28629\,
            sr => \N__46938\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26357\,
            in2 => \N__26409\,
            in3 => \N__26382\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\,
            clk => \N__47338\,
            ce => \N__28629\,
            sr => \N__46938\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26379\,
            in2 => \N__26337\,
            in3 => \N__26361\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\,
            clk => \N__47338\,
            ce => \N__28629\,
            sr => \N__46938\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26358\,
            in2 => \N__26310\,
            in3 => \N__26340\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25\,
            clk => \N__47338\,
            ce => \N__28629\,
            sr => \N__46938\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26336\,
            in2 => \N__26264\,
            in3 => \N__26313\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_27\,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\,
            clk => \N__47332\,
            ce => \N__28628\,
            sr => \N__46942\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26309\,
            in2 => \N__26219\,
            in3 => \N__26286\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\,
            clk => \N__47332\,
            ce => \N__28628\,
            sr => \N__46942\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26283\,
            in2 => \N__26265\,
            in3 => \N__26241\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\,
            clk => \N__47332\,
            ce => \N__28628\,
            sr => \N__46942\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26238\,
            in2 => \N__26220\,
            in3 => \N__26196\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29\,
            clk => \N__47332\,
            ce => \N__28628\,
            sr => \N__46942\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26598\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47332\,
            ce => \N__28628\,
            sr => \N__46942\
        );

    \current_shift_inst.timer_phase.running_RNIB31B_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33674\,
            lcout => \current_shift_inst.timer_phase.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26469\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001100"
        )
    port map (
            in0 => \N__36508\,
            in1 => \N__37329\,
            in2 => \N__37869\,
            in3 => \N__34368\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47410\,
            ce => \N__30883\,
            sr => \N__46859\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000000010000"
        )
    port map (
            in0 => \N__34369\,
            in1 => \N__37844\,
            in2 => \N__37366\,
            in3 => \N__34430\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47410\,
            ce => \N__30883\,
            sr => \N__46859\
        );

    \current_shift_inst.stop_timer_s1_RNO_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28982\,
            in1 => \N__31322\,
            in2 => \N__33156\,
            in3 => \N__31371\,
            lcout => \current_shift_inst.N_199\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_sync0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32924\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.S1_syncZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_rise_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26445\,
            in2 => \_gnd_net_\,
            in3 => \N__26453\,
            lcout => \current_shift_inst.S1_riseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_sync1_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26460\,
            lcout => \current_shift_inst.S1_syncZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_sync_prev_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26454\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.S1_sync_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30581\,
            in2 => \N__30592\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26628\,
            in2 => \N__29418\,
            in3 => \N__30729\,
            lcout => \current_shift_inst.z_i_0_31\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO\,
            carryout => \current_shift_inst.un38_control_input_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_1_c_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29388\,
            in2 => \N__28230\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_0\,
            carryout => \current_shift_inst.un38_control_input_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_2_c_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29352\,
            in2 => \N__28611\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_1\,
            carryout => \current_shift_inst.un38_control_input_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29319\,
            in2 => \N__26622\,
            in3 => \N__28671\,
            lcout => \current_shift_inst.un38_control_input_0_cry_3_c_invZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_2\,
            carryout => \current_shift_inst.un38_control_input_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_4_c_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28527\,
            in2 => \N__28545\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_3\,
            carryout => \current_shift_inst.un38_control_input_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28125\,
            in2 => \N__28482\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_4\,
            carryout => \current_shift_inst.un38_control_input_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29076\,
            in2 => \N__28215\,
            in3 => \N__26607\,
            lcout => \current_shift_inst.control_input_1_axb_0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_5\,
            carryout => \current_shift_inst.un38_control_input_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28011\,
            in2 => \N__28005\,
            in3 => \N__26775\,
            lcout => \current_shift_inst.control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28170\,
            in2 => \N__27993\,
            in3 => \N__26766\,
            lcout => \current_shift_inst.control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_7\,
            carryout => \current_shift_inst.un38_control_input_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26763\,
            in2 => \N__28134\,
            in3 => \N__26748\,
            lcout => \current_shift_inst.control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_8\,
            carryout => \current_shift_inst.un38_control_input_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26745\,
            in2 => \N__26736\,
            in3 => \N__26715\,
            lcout => \current_shift_inst.control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_9\,
            carryout => \current_shift_inst.un38_control_input_0_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26712\,
            in2 => \N__26703\,
            in3 => \N__26682\,
            lcout => \current_shift_inst.control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_10\,
            carryout => \current_shift_inst.un38_control_input_0_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28236\,
            in2 => \N__26679\,
            in3 => \N__26661\,
            lcout => \current_shift_inst.control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_11\,
            carryout => \current_shift_inst.un38_control_input_0_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28203\,
            in2 => \N__28065\,
            in3 => \N__26652\,
            lcout => \current_shift_inst.control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_12\,
            carryout => \current_shift_inst.un38_control_input_0_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28020\,
            in2 => \N__26649\,
            in3 => \N__26631\,
            lcout => \current_shift_inst.control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_13\,
            carryout => \current_shift_inst.un38_control_input_0_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28071\,
            in2 => \N__28386\,
            in3 => \N__26940\,
            lcout => \current_shift_inst.control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28119\,
            in2 => \N__28113\,
            in3 => \N__26931\,
            lcout => \current_shift_inst.control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_15\,
            carryout => \current_shift_inst.un38_control_input_0_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28353\,
            in2 => \N__28104\,
            in3 => \N__26922\,
            lcout => \current_shift_inst.control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_16\,
            carryout => \current_shift_inst.un38_control_input_0_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26919\,
            in2 => \N__28311\,
            in3 => \N__26901\,
            lcout => \current_shift_inst.control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_17\,
            carryout => \current_shift_inst.un38_control_input_0_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26898\,
            in2 => \N__26889\,
            in3 => \N__26868\,
            lcout => \current_shift_inst.control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_18\,
            carryout => \current_shift_inst.un38_control_input_0_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26865\,
            in2 => \N__26856\,
            in3 => \N__26838\,
            lcout => \current_shift_inst.control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_19\,
            carryout => \current_shift_inst.un38_control_input_0_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26835\,
            in2 => \N__26826\,
            in3 => \N__26808\,
            lcout => \current_shift_inst.control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_20\,
            carryout => \current_shift_inst.un38_control_input_0_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26805\,
            in2 => \N__26796\,
            in3 => \N__26778\,
            lcout => \current_shift_inst.control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_21\,
            carryout => \current_shift_inst.un38_control_input_0_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30228\,
            in2 => \N__27114\,
            in3 => \N__27093\,
            lcout => \current_shift_inst.control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30621\,
            in2 => \N__30609\,
            in3 => \N__27084\,
            lcout => \current_shift_inst.control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_23\,
            carryout => \current_shift_inst.un38_control_input_0_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30027\,
            in2 => \N__30744\,
            in3 => \N__27075\,
            lcout => \current_shift_inst.control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_24\,
            carryout => \current_shift_inst.un38_control_input_0_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30111\,
            in2 => \N__29151\,
            in3 => \N__27066\,
            lcout => \current_shift_inst.control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_25\,
            carryout => \current_shift_inst.un38_control_input_0_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27063\,
            in2 => \N__30369\,
            in3 => \N__27048\,
            lcout => \current_shift_inst.control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_26\,
            carryout => \current_shift_inst.un38_control_input_0_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27045\,
            in2 => \N__27036\,
            in3 => \N__27018\,
            lcout => \current_shift_inst.control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_27\,
            carryout => \current_shift_inst.un38_control_input_0_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27015\,
            in2 => \N__27006\,
            in3 => \N__26988\,
            lcout => \current_shift_inst.control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_28\,
            carryout => \current_shift_inst.un38_control_input_0_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26985\,
            in2 => \N__26973\,
            in3 => \N__26949\,
            lcout => \current_shift_inst.control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_29\,
            carryout => \current_shift_inst.un38_control_input_0_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_25_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30453\,
            in2 => \N__27255\,
            in3 => \N__27246\,
            lcout => \current_shift_inst.control_inputZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47347\,
            ce => \N__27185\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28458\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \current_shift_inst.z_5_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28571\,
            in2 => \N__27772\,
            in3 => \N__27135\,
            lcout => \current_shift_inst.z_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_1\,
            carryout => \current_shift_inst.z_5_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27698\,
            in2 => \N__28589\,
            in3 => \N__27132\,
            lcout => \current_shift_inst.z_5_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_2\,
            carryout => \current_shift_inst.z_5_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28493\,
            in2 => \N__27773\,
            in3 => \N__27129\,
            lcout => \current_shift_inst.z_5_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_3\,
            carryout => \current_shift_inst.z_5_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29087\,
            in2 => \N__27861\,
            in3 => \N__27126\,
            lcout => \current_shift_inst.z_5_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_4\,
            carryout => \current_shift_inst.z_5_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29117\,
            in2 => \N__27774\,
            in3 => \N__27123\,
            lcout => \current_shift_inst.z_5_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_5\,
            carryout => \current_shift_inst.z_5_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27705\,
            in2 => \N__28187\,
            in3 => \N__27120\,
            lcout => \current_shift_inst.z_5_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_6\,
            carryout => \current_shift_inst.z_5_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28147\,
            in2 => \N__27775\,
            in3 => \N__27117\,
            lcout => \current_shift_inst.z_5_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_7\,
            carryout => \current_shift_inst.z_5_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27326\,
            in2 => \N__27860\,
            in3 => \N__27309\,
            lcout => \current_shift_inst.z_5_9\,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \current_shift_inst.z_5_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27296\,
            in2 => \N__27838\,
            in3 => \N__27279\,
            lcout => \current_shift_inst.z_5_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_9\,
            carryout => \current_shift_inst.z_5_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28247\,
            in2 => \N__27857\,
            in3 => \N__27276\,
            lcout => \current_shift_inst.z_5_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_10\,
            carryout => \current_shift_inst.z_5_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28280\,
            in2 => \N__27839\,
            in3 => \N__27273\,
            lcout => \current_shift_inst.z_5_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_11\,
            carryout => \current_shift_inst.z_5_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28031\,
            in2 => \N__27858\,
            in3 => \N__27270\,
            lcout => \current_shift_inst.z_5_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_12\,
            carryout => \current_shift_inst.z_5_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28399\,
            in2 => \N__27840\,
            in3 => \N__27267\,
            lcout => \current_shift_inst.z_5_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_13\,
            carryout => \current_shift_inst.z_5_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28082\,
            in2 => \N__27859\,
            in3 => \N__27264\,
            lcout => \current_shift_inst.z_5_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_14\,
            carryout => \current_shift_inst.z_5_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28364\,
            in2 => \N__27841\,
            in3 => \N__27261\,
            lcout => \current_shift_inst.z_5_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_15\,
            carryout => \current_shift_inst.z_5_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28330\,
            in2 => \N__27798\,
            in3 => \N__27258\,
            lcout => \current_shift_inst.z_5_17\,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \current_shift_inst.z_5_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27465\,
            in2 => \N__27826\,
            in3 => \N__27441\,
            lcout => \current_shift_inst.z_5_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_17\,
            carryout => \current_shift_inst.z_5_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27422\,
            in2 => \N__27799\,
            in3 => \N__27411\,
            lcout => \current_shift_inst.z_5_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_18\,
            carryout => \current_shift_inst.z_5_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27395\,
            in2 => \N__27827\,
            in3 => \N__27384\,
            lcout => \current_shift_inst.z_5_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_19\,
            carryout => \current_shift_inst.z_5_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27362\,
            in2 => \N__27800\,
            in3 => \N__27351\,
            lcout => \current_shift_inst.z_5_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_20\,
            carryout => \current_shift_inst.z_5_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30331\,
            in2 => \N__27828\,
            in3 => \N__27348\,
            lcout => \current_shift_inst.z_5_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_21\,
            carryout => \current_shift_inst.z_5_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30239\,
            in2 => \N__27801\,
            in3 => \N__27345\,
            lcout => \current_shift_inst.z_5_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_22\,
            carryout => \current_shift_inst.z_5_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30664\,
            in2 => \N__27829\,
            in3 => \N__27342\,
            lcout => \current_shift_inst.z_5_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_23\,
            carryout => \current_shift_inst.z_5_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30057\,
            in2 => \N__27666\,
            in3 => \N__27339\,
            lcout => \current_shift_inst.z_5_25\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \current_shift_inst.z_5_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30432\,
            in2 => \N__27669\,
            in3 => \N__27948\,
            lcout => \current_shift_inst.z_5_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_25\,
            carryout => \current_shift_inst.z_5_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27929\,
            in2 => \N__27667\,
            in3 => \N__27918\,
            lcout => \current_shift_inst.z_5_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_26\,
            carryout => \current_shift_inst.z_5_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27902\,
            in2 => \N__27670\,
            in3 => \N__27891\,
            lcout => \current_shift_inst.z_5_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_27\,
            carryout => \current_shift_inst.z_5_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27875\,
            in2 => \N__27668\,
            in3 => \N__27864\,
            lcout => \current_shift_inst.z_5_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_28\,
            carryout => \current_shift_inst.z_5_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30517\,
            in2 => \N__27671\,
            in3 => \N__27489\,
            lcout => \current_shift_inst.z_5_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_29\,
            carryout => \current_shift_inst.z_5_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27486\,
            lcout => \current_shift_inst.z_5_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27483\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__36752\,
            in1 => \N__37374\,
            in2 => \_gnd_net_\,
            in3 => \N__37698\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47418\,
            ce => \N__30881\,
            sr => \N__46826\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37349\,
            in1 => \N__37160\,
            in2 => \N__37242\,
            in3 => \N__37474\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47411\,
            ce => \N__30885\,
            sr => \N__46831\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__37852\,
            in1 => \N__36831\,
            in2 => \_gnd_net_\,
            in3 => \N__37695\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47411\,
            ce => \N__30885\,
            sr => \N__46831\
        );

    \delay_measurement_inst.delay_hc_reg_22_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__41895\,
            in1 => \N__40800\,
            in2 => \N__27969\,
            in3 => \N__39040\,
            lcout => measured_delay_hc_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47402\,
            ce => 'H',
            sr => \N__46840\
        );

    \delay_measurement_inst.delay_hc_reg_20_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__28958\,
            in1 => \N__40799\,
            in2 => \N__41901\,
            in3 => \N__39039\,
            lcout => measured_delay_hc_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47402\,
            ce => 'H',
            sr => \N__46840\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_5_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36562\,
            in2 => \_gnd_net_\,
            in3 => \N__37038\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__27964\,
            in1 => \N__28897\,
            in2 => \N__27984\,
            in3 => \N__31212\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto31_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__37842\,
            in1 => \N__29028\,
            in2 => \N__27981\,
            in3 => \N__29052\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27978\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__28898\,
            in1 => \N__27965\,
            in2 => \N__28959\,
            in3 => \N__29051\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto30_2\,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto30_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto31_c_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27951\,
            in3 => \N__37843\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.target_time_11_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37485\,
            in1 => \N__36655\,
            in2 => \N__37367\,
            in3 => \N__37141\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47384\,
            ce => \N__37107\,
            sr => \N__46851\
        );

    \current_shift_inst.meas_state_0_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110101010"
        )
    port map (
            in0 => \N__31373\,
            in1 => \N__28987\,
            in2 => \N__33155\,
            in3 => \N__31334\,
            lcout => \current_shift_inst.meas_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47377\,
            ce => 'H',
            sr => \N__46860\
        );

    \current_shift_inst.phase_valid_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100011111000"
        )
    port map (
            in0 => \N__31333\,
            in1 => \N__31425\,
            in2 => \N__28994\,
            in3 => \N__31372\,
            lcout => \current_shift_inst.phase_validZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47377\,
            ce => 'H',
            sr => \N__46860\
        );

    \delay_measurement_inst.delay_hc_reg_23_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__29067\,
            in1 => \N__40801\,
            in2 => \N__41852\,
            in3 => \N__39037\,
            lcout => measured_delay_hc_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47377\,
            ce => 'H',
            sr => \N__46860\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__29522\,
            in1 => \N__28049\,
            in2 => \N__29571\,
            in3 => \N__28302\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28053\,
            in3 => \N__29521\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_27_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__29172\,
            in1 => \N__40802\,
            in2 => \N__41900\,
            in3 => \N__39038\,
            lcout => measured_delay_hc_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47371\,
            ce => 'H',
            sr => \N__46872\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__29217\,
            in1 => \N__28195\,
            in2 => \N__29136\,
            in3 => \N__29759\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29132\,
            in2 => \_gnd_net_\,
            in3 => \N__29216\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28196\,
            in2 => \_gnd_net_\,
            in3 => \N__29758\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29101\,
            in2 => \_gnd_net_\,
            in3 => \N__29249\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIER9V_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28300\,
            in2 => \_gnd_net_\,
            in3 => \N__29567\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111000011"
        )
    port map (
            in0 => \N__28197\,
            in1 => \N__28160\,
            in2 => \N__29717\,
            in3 => \N__29760\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28164\,
            in3 => \N__29710\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__28515\,
            in1 => \N__29248\,
            in2 => \N__29292\,
            in3 => \N__29102\,
            lcout => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__28095\,
            in1 => \N__28375\,
            in2 => \N__30015\,
            in3 => \N__29978\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5M161_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28094\,
            in2 => \_gnd_net_\,
            in3 => \N__30010\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI190J_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28376\,
            in2 => \_gnd_net_\,
            in3 => \N__29977\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__28416\,
            in1 => \N__28093\,
            in2 => \N__29487\,
            in3 => \N__30011\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28415\,
            in2 => \_gnd_net_\,
            in3 => \N__29483\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__28377\,
            in1 => \N__28346\,
            in2 => \N__29982\,
            in3 => \N__29942\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIBU361_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29941\,
            in2 => \_gnd_net_\,
            in3 => \N__28347\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__29606\,
            in1 => \N__28301\,
            in2 => \N__28269\,
            in3 => \N__29563\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31869\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47349\,
            ce => \N__31694\,
            sr => \N__46900\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31836\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47349\,
            ce => \N__31694\,
            sr => \N__46900\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31673\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47349\,
            ce => \N__31694\,
            sr => \N__46900\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31674\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47349\,
            ce => \N__31694\,
            sr => \N__46900\
        );

    \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__30560\,
            in1 => \N__28451\,
            in2 => \_gnd_net_\,
            in3 => \N__29384\,
            lcout => \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28701\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47340\,
            ce => \N__28630\,
            sr => \N__46908\
        );

    \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100101"
        )
    port map (
            in0 => \N__28595\,
            in1 => \N__28566\,
            in2 => \N__30579\,
            in3 => \N__28450\,
            lcout => \current_shift_inst.N_1633_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28659\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47340\,
            ce => \N__28630\,
            sr => \N__46908\
        );

    \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101010011010"
        )
    port map (
            in0 => \N__28570\,
            in1 => \N__28452\,
            in2 => \N__30580\,
            in3 => \N__29348\,
            lcout => \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__28453\,
            in1 => \N__28596\,
            in2 => \N__28572\,
            in3 => \N__30564\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3\,
            ltout => \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28507\,
            in2 => \N__28530\,
            in3 => \N__29280\,
            lcout => \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__29281\,
            in1 => \_gnd_net_\,
            in2 => \N__28514\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29442\,
            in1 => \N__29408\,
            in2 => \N__28467\,
            in3 => \_gnd_net_\,
            lcout => \G_406\,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \current_shift_inst.z_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29380\,
            in2 => \N__28425\,
            in3 => \N__28457\,
            lcout => \G_405\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_0\,
            carryout => \current_shift_inst.z_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_2_c_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29344\,
            in2 => \N__28764\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_1\,
            carryout => \current_shift_inst.z_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_3_c_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29312\,
            in2 => \N__28755\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_2\,
            carryout => \current_shift_inst.z_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_4_c_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28746\,
            in2 => \N__29285\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_3\,
            carryout => \current_shift_inst.z_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_5_c_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29239\,
            in2 => \N__28740\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_4\,
            carryout => \current_shift_inst.z_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_6_c_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29203\,
            in2 => \N__28731\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_5\,
            carryout => \current_shift_inst.z_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_7_c_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28722\,
            in2 => \N__29749\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_6\,
            carryout => \current_shift_inst.z_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_8_c_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28716\,
            in2 => \N__29701\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \current_shift_inst.z_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_9_c_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28707\,
            in2 => \N__29659\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_8\,
            carryout => \current_shift_inst.z_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_10_c_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28821\,
            in2 => \N__29627\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_9\,
            carryout => \current_shift_inst.z_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_11_c_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28815\,
            in2 => \N__29593\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_10\,
            carryout => \current_shift_inst.z_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_12_c_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28809\,
            in2 => \N__29559\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_11\,
            carryout => \current_shift_inst.z_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_13_c_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28803\,
            in2 => \N__29512\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_12\,
            carryout => \current_shift_inst.z_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_14_c_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28797\,
            in2 => \N__29473\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_13\,
            carryout => \current_shift_inst.z_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_15_c_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28791\,
            in2 => \N__30002\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_14\,
            carryout => \current_shift_inst.z_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_16_c_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28785\,
            in2 => \N__29969\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_19_0_\,
            carryout => \current_shift_inst.z_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_17_c_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28776\,
            in2 => \N__29931\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_16\,
            carryout => \current_shift_inst.z_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_18_c_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28770\,
            in2 => \N__29893\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_17\,
            carryout => \current_shift_inst.z_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_19_c_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28875\,
            in2 => \N__29852\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_18\,
            carryout => \current_shift_inst.z_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_20_c_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29819\,
            in2 => \N__28869\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_19\,
            carryout => \current_shift_inst.z_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_21_c_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28860\,
            in2 => \N__29792\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_20\,
            carryout => \current_shift_inst.z_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_22_c_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28854\,
            in2 => \N__30280\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_21\,
            carryout => \current_shift_inst.z_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_23_c_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28848\,
            in2 => \N__30312\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_22\,
            carryout => \current_shift_inst.z_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_24_c_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28842\,
            in2 => \N__30647\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_20_0_\,
            carryout => \current_shift_inst.z_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_25_c_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30093\,
            in2 => \N__28836\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_24\,
            carryout => \current_shift_inst.z_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_26_c_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28827\,
            in2 => \N__30398\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_25\,
            carryout => \current_shift_inst.z_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_27_c_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28938\,
            in2 => \N__30188\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_26\,
            carryout => \current_shift_inst.z_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_28_c_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28932\,
            in2 => \N__30158\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_27\,
            carryout => \current_shift_inst.z_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_29_c_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30128\,
            in2 => \N__28926\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_28\,
            carryout => \current_shift_inst.z_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_30_c_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30469\,
            in2 => \N__28917\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_29\,
            carryout => \current_shift_inst.z_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_s_31_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30593\,
            in1 => \N__28908\,
            in2 => \N__30500\,
            in3 => \N__28902\,
            lcout => \current_shift_inst.z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__37848\,
            in1 => \N__37751\,
            in2 => \_gnd_net_\,
            in3 => \N__37689\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47419\,
            ce => \N__30887\,
            sr => \N__46816\
        );

    \delay_measurement_inst.delay_hc_reg_21_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__41880\,
            in1 => \N__40759\,
            in2 => \N__28899\,
            in3 => \N__39042\,
            lcout => measured_delay_hc_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47412\,
            ce => 'H',
            sr => \N__46821\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto31_d_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110111"
        )
    port map (
            in0 => \N__40554\,
            in1 => \N__31191\,
            in2 => \N__37870\,
            in3 => \N__31443\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0\,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_0_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37361\,
            in1 => \N__37161\,
            in2 => \N__28878\,
            in3 => \N__36992\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47403\,
            ce => \N__30882\,
            sr => \N__46827\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37162\,
            in1 => \N__36606\,
            in2 => \N__37409\,
            in3 => \N__37469\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47403\,
            ce => \N__30882\,
            sr => \N__46827\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37471\,
            in1 => \N__37323\,
            in2 => \N__36660\,
            in3 => \N__37155\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47394\,
            ce => \N__30856\,
            sr => \N__46832\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37322\,
            in1 => \N__37154\,
            in2 => \N__40563\,
            in3 => \N__37473\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47394\,
            ce => \N__30856\,
            sr => \N__46832\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37472\,
            in1 => \N__37324\,
            in2 => \N__37566\,
            in3 => \N__37156\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47394\,
            ce => \N__30856\,
            sr => \N__46832\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36702\,
            in1 => \N__37153\,
            in2 => \N__37365\,
            in3 => \N__37470\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47394\,
            ce => \N__30856\,
            sr => \N__46832\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__37651\,
            in1 => \N__36792\,
            in2 => \_gnd_net_\,
            in3 => \N__37328\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47394\,
            ce => \N__30856\,
            sr => \N__46832\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__37321\,
            in1 => \N__37047\,
            in2 => \_gnd_net_\,
            in3 => \N__37652\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47394\,
            ce => \N__30856\,
            sr => \N__46832\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__36230\,
            in1 => \N__32735\,
            in2 => \_gnd_net_\,
            in3 => \N__32813\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__28954\,
            in1 => \N__40541\,
            in2 => \_gnd_net_\,
            in3 => \N__36827\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36563\,
            in1 => \N__36791\,
            in2 => \N__36512\,
            in3 => \N__34422\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_14_3_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32949\,
            in2 => \_gnd_net_\,
            in3 => \N__29066\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_14_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__32966\,
            in1 => \N__32895\,
            in2 => \N__29055\,
            in3 => \N__29160\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36784\,
            in1 => \N__36751\,
            in2 => \N__36516\,
            in3 => \N__37561\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__36241\,
            in1 => \N__32803\,
            in2 => \_gnd_net_\,
            in3 => \N__32760\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto3_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__36875\,
            in1 => \N__36915\,
            in2 => \_gnd_net_\,
            in3 => \N__40886\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlt30_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_14_6_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__29043\,
            in1 => \N__31203\,
            in2 => \N__29037\,
            in3 => \N__29034\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33370\,
            in2 => \_gnd_net_\,
            in3 => \N__33114\,
            lcout => \current_shift_inst.timer_s1.N_187_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.start_timer_s1_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111111001100"
        )
    port map (
            in0 => \N__28986\,
            in1 => \N__33141\,
            in2 => \N__31344\,
            in3 => \N__31392\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47372\,
            ce => \N__34786\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__33140\,
            in1 => \N__33371\,
            in2 => \_gnd_net_\,
            in3 => \N__33115\,
            lcout => \current_shift_inst.timer_s1.N_191_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_phase_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111000000"
        )
    port map (
            in0 => \N__31393\,
            in1 => \N__31342\,
            in2 => \N__31421\,
            in3 => \N__33729\,
            lcout => \current_shift_inst.stop_timer_phaseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47372\,
            ce => \N__34786\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33095\,
            in1 => \N__33068\,
            in2 => \N__46988\,
            in3 => \N__34291\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47364\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_14_4_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31286\,
            in1 => \N__31301\,
            in2 => \N__31275\,
            in3 => \N__29171\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30072\,
            in2 => \_gnd_net_\,
            in3 => \N__30099\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__29250\,
            in1 => \N__29131\,
            in2 => \N__29106\,
            in3 => \N__29210\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_0_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__45673\,
            in1 => \N__45379\,
            in2 => \N__45599\,
            in3 => \N__41089\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47350\,
            ce => \N__34793\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_1_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__41090\,
            in1 => \N__45590\,
            in2 => \N__45413\,
            in3 => \N__45674\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47350\,
            ce => \N__34793\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_state_0_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__36302\,
            in1 => \N__35119\,
            in2 => \_gnd_net_\,
            in3 => \N__35106\,
            lcout => \delay_measurement_inst.tr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47350\,
            ce => \N__34793\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.hc_state_0_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__33096\,
            in1 => \N__33061\,
            in2 => \_gnd_net_\,
            in3 => \N__34293\,
            lcout => \delay_measurement_inst.hc_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47350\,
            ce => \N__34793\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29184\,
            lcout => \current_shift_inst.un4_control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29178\,
            lcout => \current_shift_inst.un4_control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31260\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__37697\,
            in1 => \N__37885\,
            in2 => \_gnd_net_\,
            in3 => \N__37941\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47341\,
            ce => \N__30886\,
            sr => \N__46887\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__37884\,
            in1 => \N__36564\,
            in2 => \_gnd_net_\,
            in3 => \N__37696\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47341\,
            ce => \N__30886\,
            sr => \N__46887\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31503\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31494\,
            lcout => \current_shift_inst.un4_control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31485\,
            lcout => \current_shift_inst.un4_control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31476\,
            lcout => \current_shift_inst.un4_control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31467\,
            lcout => \current_shift_inst.un4_control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31458\,
            lcout => \current_shift_inst.un4_control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29451\,
            in2 => \N__29441\,
            in3 => \N__29440\,
            lcout => \current_shift_inst.un38_control_input_0\,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29397\,
            in2 => \_gnd_net_\,
            in3 => \N__29364\,
            lcout => \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_1\,
            carryout => \current_shift_inst.un4_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29361\,
            in2 => \_gnd_net_\,
            in3 => \N__29328\,
            lcout => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_2\,
            carryout => \current_shift_inst.un4_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29325\,
            in2 => \_gnd_net_\,
            in3 => \N__29301\,
            lcout => \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_3\,
            carryout => \current_shift_inst.un4_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29298\,
            in2 => \_gnd_net_\,
            in3 => \N__29259\,
            lcout => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_4\,
            carryout => \current_shift_inst.un4_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29256\,
            in2 => \_gnd_net_\,
            in3 => \N__29226\,
            lcout => \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_5\,
            carryout => \current_shift_inst.un4_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29223\,
            in2 => \_gnd_net_\,
            in3 => \N__29187\,
            lcout => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_6\,
            carryout => \current_shift_inst.un4_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29766\,
            in2 => \_gnd_net_\,
            in3 => \N__29730\,
            lcout => \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_7\,
            carryout => \current_shift_inst.un4_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29727\,
            in2 => \_gnd_net_\,
            in3 => \N__29676\,
            lcout => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33186\,
            in2 => \_gnd_net_\,
            in3 => \N__29640\,
            lcout => \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_9\,
            carryout => \current_shift_inst.un4_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33168\,
            in2 => \_gnd_net_\,
            in3 => \N__29610\,
            lcout => \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_10\,
            carryout => \current_shift_inst.un4_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33504\,
            in2 => \_gnd_net_\,
            in3 => \N__29574\,
            lcout => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_11\,
            carryout => \current_shift_inst.un4_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33468\,
            in2 => \_gnd_net_\,
            in3 => \N__29532\,
            lcout => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_12\,
            carryout => \current_shift_inst.un4_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33450\,
            in2 => \_gnd_net_\,
            in3 => \N__29490\,
            lcout => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_13\,
            carryout => \current_shift_inst.un4_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33420\,
            in2 => \_gnd_net_\,
            in3 => \N__29454\,
            lcout => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_14\,
            carryout => \current_shift_inst.un4_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33402\,
            in2 => \_gnd_net_\,
            in3 => \N__29985\,
            lcout => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_15\,
            carryout => \current_shift_inst.un4_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33384\,
            in2 => \_gnd_net_\,
            in3 => \N__29952\,
            lcout => \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33486\,
            in2 => \_gnd_net_\,
            in3 => \N__29910\,
            lcout => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_17\,
            carryout => \current_shift_inst.un4_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31593\,
            in3 => \N__29868\,
            lcout => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_18\,
            carryout => \current_shift_inst.un4_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31623\,
            in2 => \_gnd_net_\,
            in3 => \N__29835\,
            lcout => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_19\,
            carryout => \current_shift_inst.un4_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33204\,
            in2 => \_gnd_net_\,
            in3 => \N__29808\,
            lcout => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_20\,
            carryout => \current_shift_inst.un4_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31875\,
            in2 => \_gnd_net_\,
            in3 => \N__29775\,
            lcout => \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_21\,
            carryout => \current_shift_inst.un4_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33432\,
            in2 => \_gnd_net_\,
            in3 => \N__29772\,
            lcout => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_22\,
            carryout => \current_shift_inst.un4_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32985\,
            in2 => \_gnd_net_\,
            in3 => \N__29769\,
            lcout => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_23\,
            carryout => \current_shift_inst.un4_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31890\,
            in2 => \_gnd_net_\,
            in3 => \N__30213\,
            lcout => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31575\,
            in2 => \_gnd_net_\,
            in3 => \N__30210\,
            lcout => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_25\,
            carryout => \current_shift_inst.un4_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31563\,
            in2 => \_gnd_net_\,
            in3 => \N__30207\,
            lcout => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_26\,
            carryout => \current_shift_inst.un4_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31638\,
            in2 => \_gnd_net_\,
            in3 => \N__30171\,
            lcout => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_27\,
            carryout => \current_shift_inst.un4_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31653\,
            in2 => \_gnd_net_\,
            in3 => \N__30141\,
            lcout => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_28\,
            carryout => \current_shift_inst.un4_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31611\,
            in3 => \N__30117\,
            lcout => \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_29\,
            carryout => \current_shift_inst.un4_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__30585\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30114\,
            lcout => \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30098\,
            in1 => \N__30439\,
            in2 => \N__30071\,
            in3 => \N__30394\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30646\,
            in1 => \N__30094\,
            in2 => \N__30684\,
            in3 => \N__30070\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5S981_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__30645\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30679\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_i_31_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30722\,
            lcout => \current_shift_inst.z_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__30683\,
            in1 => \N__30315\,
            in2 => \N__30648\,
            in3 => \N__30254\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__30314\,
            in1 => \_gnd_net_\,
            in2 => \N__30255\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIU73K_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_0_25_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__30594\,
            in1 => \N__30525\,
            in2 => \N__30501\,
            in3 => \N__30473\,
            lcout => \current_shift_inst.un38_control_input_0_axb_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30440\,
            in2 => \_gnd_net_\,
            in3 => \N__30393\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30350\,
            in1 => \N__30313\,
            in2 => \N__30291\,
            in3 => \N__30250\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPB581_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.running_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__33705\,
            in1 => \N__33673\,
            in2 => \_gnd_net_\,
            in3 => \N__33743\,
            lcout => \current_shift_inst.timer_phase.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47310\,
            ce => 'H',
            sr => \N__46934\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30900\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto9_c_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__37936\,
            in1 => \N__37234\,
            in2 => \_gnd_net_\,
            in3 => \N__37046\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto9_cZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto14_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__36753\,
            in1 => \N__34305\,
            in2 => \N__30891\,
            in3 => \N__34323\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111111"
        )
    port map (
            in0 => \N__37668\,
            in1 => \N__36871\,
            in2 => \_gnd_net_\,
            in3 => \N__37373\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47401\,
            ce => \N__30884\,
            sr => \N__46817\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__37667\,
            in1 => \N__37372\,
            in2 => \_gnd_net_\,
            in3 => \N__36913\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47401\,
            ce => \N__30884\,
            sr => \N__46817\
        );

    \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010101010"
        )
    port map (
            in0 => \N__37371\,
            in1 => \_gnd_net_\,
            in2 => \N__36955\,
            in3 => \N__37666\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47401\,
            ce => \N__30884\,
            sr => \N__46817\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30795\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30774\,
            in2 => \N__30786\,
            in3 => \N__33820\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30750\,
            in2 => \N__30768\,
            in3 => \N__33803\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31038\,
            in2 => \N__31050\,
            in3 => \N__33767\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31020\,
            in2 => \N__31032\,
            in3 => \N__34070\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30999\,
            in2 => \N__31014\,
            in3 => \N__34049\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30978\,
            in2 => \N__30993\,
            in3 => \N__34028\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30960\,
            in2 => \N__30972\,
            in3 => \N__34004\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30939\,
            in2 => \N__30954\,
            in3 => \N__33980\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30924\,
            in2 => \N__30933\,
            in3 => \N__33953\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33932\,
            in1 => \N__30906\,
            in2 => \N__30918\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31161\,
            in2 => \N__31173\,
            in3 => \N__34253\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31146\,
            in2 => \N__31155\,
            in3 => \N__34229\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31128\,
            in2 => \N__31140\,
            in3 => \N__34208\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31107\,
            in2 => \N__31122\,
            in3 => \N__34187\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31089\,
            in2 => \N__31101\,
            in3 => \N__34166\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31074\,
            in2 => \N__31083\,
            in3 => \N__34143\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34115\,
            in1 => \N__31056\,
            in2 => \N__31068\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31242\,
            in2 => \N__31254\,
            in3 => \N__34094\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31221\,
            in2 => \N__31236\,
            in3 => \N__34346\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31215\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37223\,
            in1 => \N__36609\,
            in2 => \N__37940\,
            in3 => \N__36656\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34634\,
            in1 => \N__33824\,
            in2 => \_gnd_net_\,
            in3 => \N__34582\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32796\,
            in2 => \_gnd_net_\,
            in3 => \N__32682\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36951\,
            in1 => \N__36701\,
            in2 => \N__34431\,
            in3 => \N__37752\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_sync_prev_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33012\,
            lcout => \current_shift_inst.S3_sync_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_rise_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__33011\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31197\,
            lcout => \current_shift_inst.S3_riseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto19_3_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001001100"
        )
    port map (
            in0 => \N__40555\,
            in1 => \N__34381\,
            in2 => \N__31190\,
            in3 => \N__31442\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt31_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.start_timer_phase_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110101001100"
        )
    port map (
            in0 => \N__31335\,
            in1 => \N__33689\,
            in2 => \N__31420\,
            in3 => \N__31394\,
            lcout => \current_shift_inst.start_timer_phaseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47363\,
            ce => \N__34785\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_1_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001100010"
        )
    port map (
            in0 => \N__32750\,
            in1 => \N__32812\,
            in2 => \N__36246\,
            in3 => \N__34589\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47363\,
            ce => \N__34785\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_s1_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111001100"
        )
    port map (
            in0 => \N__31395\,
            in1 => \N__31353\,
            in2 => \N__31343\,
            in3 => \N__33117\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47363\,
            ce => \N__34785\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.prev_hc_sig_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34292\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.prev_hc_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47356\,
            ce => 'H',
            sr => \N__46852\
        );

    \delay_measurement_inst.delay_hc_reg_28_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__31302\,
            in1 => \N__40834\,
            in2 => \N__41892\,
            in3 => \N__39027\,
            lcout => measured_delay_hc_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47356\,
            ce => 'H',
            sr => \N__46852\
        );

    \delay_measurement_inst.delay_hc_reg_29_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__39028\,
            in1 => \N__41869\,
            in2 => \N__31290\,
            in3 => \N__40836\,
            lcout => measured_delay_hc_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47356\,
            ce => 'H',
            sr => \N__46852\
        );

    \delay_measurement_inst.delay_hc_reg_30_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__31274\,
            in1 => \N__40835\,
            in2 => \N__41893\,
            in3 => \N__39029\,
            lcout => measured_delay_hc_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47356\,
            ce => 'H',
            sr => \N__46852\
        );

    \phase_controller_inst1.T01_er_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34458\,
            lcout => shift_flag_start,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47348\,
            ce => \N__33024\,
            sr => \N__46861\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31802\,
            in2 => \N__31868\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__47339\,
            ce => \N__31698\,
            sr => \N__46873\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31781\,
            in2 => \N__31835\,
            in3 => \N__31497\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__47339\,
            ce => \N__31698\,
            sr => \N__46873\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31803\,
            in2 => \N__31761\,
            in3 => \N__31488\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__47339\,
            ce => \N__31698\,
            sr => \N__46873\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31782\,
            in2 => \N__31731\,
            in3 => \N__31479\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__47339\,
            ce => \N__31698\,
            sr => \N__46873\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31757\,
            in2 => \N__32138\,
            in3 => \N__31470\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__47339\,
            ce => \N__31698\,
            sr => \N__46873\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31727\,
            in2 => \N__32111\,
            in3 => \N__31461\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__47339\,
            ce => \N__31698\,
            sr => \N__46873\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32081\,
            in2 => \N__32139\,
            in3 => \N__31452\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__47339\,
            ce => \N__31698\,
            sr => \N__46873\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32054\,
            in2 => \N__32112\,
            in3 => \N__31449\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__47339\,
            ce => \N__31698\,
            sr => \N__46873\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32082\,
            in2 => \N__32030\,
            in3 => \N__31446\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__47333\,
            ce => \N__31697\,
            sr => \N__46881\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32055\,
            in2 => \N__32003\,
            in3 => \N__31530\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__47333\,
            ce => \N__31697\,
            sr => \N__46881\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31976\,
            in2 => \N__32031\,
            in3 => \N__31527\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__47333\,
            ce => \N__31697\,
            sr => \N__46881\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31955\,
            in2 => \N__32004\,
            in3 => \N__31524\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__47333\,
            ce => \N__31697\,
            sr => \N__46881\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31977\,
            in2 => \N__31932\,
            in3 => \N__31521\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__47333\,
            ce => \N__31697\,
            sr => \N__46881\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31956\,
            in2 => \N__32357\,
            in3 => \N__31518\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__47333\,
            ce => \N__31697\,
            sr => \N__46881\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31928\,
            in2 => \N__32328\,
            in3 => \N__31515\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__47333\,
            ce => \N__31697\,
            sr => \N__46881\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32297\,
            in2 => \N__32358\,
            in3 => \N__31512\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__47333\,
            ce => \N__31697\,
            sr => \N__46881\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32327\,
            in2 => \N__32270\,
            in3 => \N__31509\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__47327\,
            ce => \N__31696\,
            sr => \N__46888\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32298\,
            in2 => \N__32240\,
            in3 => \N__31506\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__47327\,
            ce => \N__31696\,
            sr => \N__46888\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32210\,
            in2 => \N__32271\,
            in3 => \N__31557\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__47327\,
            ce => \N__31696\,
            sr => \N__46888\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32186\,
            in2 => \N__32241\,
            in3 => \N__31554\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__47327\,
            ce => \N__31696\,
            sr => \N__46888\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32211\,
            in2 => \N__32165\,
            in3 => \N__31551\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__47327\,
            ce => \N__31696\,
            sr => \N__46888\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32187\,
            in2 => \N__32591\,
            in3 => \N__31548\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__47327\,
            ce => \N__31696\,
            sr => \N__46888\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32561\,
            in2 => \N__32166\,
            in3 => \N__31545\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__47327\,
            ce => \N__31696\,
            sr => \N__46888\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32531\,
            in2 => \N__32592\,
            in3 => \N__31542\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__47327\,
            ce => \N__31696\,
            sr => \N__46888\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32562\,
            in2 => \N__32504\,
            in3 => \N__31539\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__47322\,
            ce => \N__31695\,
            sr => \N__46901\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32474\,
            in2 => \N__32535\,
            in3 => \N__31536\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__47322\,
            ce => \N__31695\,
            sr => \N__46901\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32454\,
            in2 => \N__32505\,
            in3 => \N__31533\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__47322\,
            ce => \N__31695\,
            sr => \N__46901\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32475\,
            in2 => \N__32430\,
            in3 => \N__31701\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__47322\,
            ce => \N__31695\,
            sr => \N__46901\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31677\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31659\,
            lcout => \current_shift_inst.un4_control_input_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31644\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31632\,
            lcout => \current_shift_inst.un4_control_input_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31617\,
            lcout => \current_shift_inst.un4_control_input_axb_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31602\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31584\,
            lcout => \current_shift_inst.un4_control_input_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31569\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31899\,
            lcout => \current_shift_inst.un4_control_input_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31884\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33315\,
            in1 => \N__31858\,
            in2 => \_gnd_net_\,
            in3 => \N__31839\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_12_19_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__47315\,
            ce => \N__32403\,
            sr => \N__46914\
        );

    \current_shift_inst.timer_s1.counter_1_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33307\,
            in1 => \N__31825\,
            in2 => \_gnd_net_\,
            in3 => \N__31806\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__47315\,
            ce => \N__32403\,
            sr => \N__46914\
        );

    \current_shift_inst.timer_s1.counter_2_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33316\,
            in1 => \N__31801\,
            in2 => \_gnd_net_\,
            in3 => \N__31785\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__47315\,
            ce => \N__32403\,
            sr => \N__46914\
        );

    \current_shift_inst.timer_s1.counter_3_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33308\,
            in1 => \N__31780\,
            in2 => \_gnd_net_\,
            in3 => \N__31764\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__47315\,
            ce => \N__32403\,
            sr => \N__46914\
        );

    \current_shift_inst.timer_s1.counter_4_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33317\,
            in1 => \N__31753\,
            in2 => \_gnd_net_\,
            in3 => \N__31734\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__47315\,
            ce => \N__32403\,
            sr => \N__46914\
        );

    \current_shift_inst.timer_s1.counter_5_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33309\,
            in1 => \N__31723\,
            in2 => \_gnd_net_\,
            in3 => \N__31704\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__47315\,
            ce => \N__32403\,
            sr => \N__46914\
        );

    \current_shift_inst.timer_s1.counter_6_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33318\,
            in1 => \N__32131\,
            in2 => \_gnd_net_\,
            in3 => \N__32115\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__47315\,
            ce => \N__32403\,
            sr => \N__46914\
        );

    \current_shift_inst.timer_s1.counter_7_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33310\,
            in1 => \N__32099\,
            in2 => \_gnd_net_\,
            in3 => \N__32085\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__47315\,
            ce => \N__32403\,
            sr => \N__46914\
        );

    \current_shift_inst.timer_s1.counter_8_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33335\,
            in1 => \N__32074\,
            in2 => \_gnd_net_\,
            in3 => \N__32058\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__47312\,
            ce => \N__32411\,
            sr => \N__46921\
        );

    \current_shift_inst.timer_s1.counter_9_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33322\,
            in1 => \N__32053\,
            in2 => \_gnd_net_\,
            in3 => \N__32034\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__47312\,
            ce => \N__32411\,
            sr => \N__46921\
        );

    \current_shift_inst.timer_s1.counter_10_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33332\,
            in1 => \N__32023\,
            in2 => \_gnd_net_\,
            in3 => \N__32007\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__47312\,
            ce => \N__32411\,
            sr => \N__46921\
        );

    \current_shift_inst.timer_s1.counter_11_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33319\,
            in1 => \N__31996\,
            in2 => \_gnd_net_\,
            in3 => \N__31980\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__47312\,
            ce => \N__32411\,
            sr => \N__46921\
        );

    \current_shift_inst.timer_s1.counter_12_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33333\,
            in1 => \N__31975\,
            in2 => \_gnd_net_\,
            in3 => \N__31959\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__47312\,
            ce => \N__32411\,
            sr => \N__46921\
        );

    \current_shift_inst.timer_s1.counter_13_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33320\,
            in1 => \N__31949\,
            in2 => \_gnd_net_\,
            in3 => \N__31935\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__47312\,
            ce => \N__32411\,
            sr => \N__46921\
        );

    \current_shift_inst.timer_s1.counter_14_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33334\,
            in1 => \N__31924\,
            in2 => \_gnd_net_\,
            in3 => \N__31902\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__47312\,
            ce => \N__32411\,
            sr => \N__46921\
        );

    \current_shift_inst.timer_s1.counter_15_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33321\,
            in1 => \N__32345\,
            in2 => \_gnd_net_\,
            in3 => \N__32331\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__47312\,
            ce => \N__32411\,
            sr => \N__46921\
        );

    \current_shift_inst.timer_s1.counter_16_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33311\,
            in1 => \N__32317\,
            in2 => \_gnd_net_\,
            in3 => \N__32301\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_12_21_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__47309\,
            ce => \N__32404\,
            sr => \N__46925\
        );

    \current_shift_inst.timer_s1.counter_17_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33342\,
            in1 => \N__32290\,
            in2 => \_gnd_net_\,
            in3 => \N__32274\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__47309\,
            ce => \N__32404\,
            sr => \N__46925\
        );

    \current_shift_inst.timer_s1.counter_18_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33312\,
            in1 => \N__32258\,
            in2 => \_gnd_net_\,
            in3 => \N__32244\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__47309\,
            ce => \N__32404\,
            sr => \N__46925\
        );

    \current_shift_inst.timer_s1.counter_19_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33343\,
            in1 => \N__32228\,
            in2 => \_gnd_net_\,
            in3 => \N__32214\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__47309\,
            ce => \N__32404\,
            sr => \N__46925\
        );

    \current_shift_inst.timer_s1.counter_20_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33313\,
            in1 => \N__32204\,
            in2 => \_gnd_net_\,
            in3 => \N__32190\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__47309\,
            ce => \N__32404\,
            sr => \N__46925\
        );

    \current_shift_inst.timer_s1.counter_21_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33344\,
            in1 => \N__32185\,
            in2 => \_gnd_net_\,
            in3 => \N__32169\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__47309\,
            ce => \N__32404\,
            sr => \N__46925\
        );

    \current_shift_inst.timer_s1.counter_22_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33314\,
            in1 => \N__32158\,
            in2 => \_gnd_net_\,
            in3 => \N__32142\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__47309\,
            ce => \N__32404\,
            sr => \N__46925\
        );

    \current_shift_inst.timer_s1.counter_23_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33345\,
            in1 => \N__32579\,
            in2 => \_gnd_net_\,
            in3 => \N__32565\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__47309\,
            ce => \N__32404\,
            sr => \N__46925\
        );

    \current_shift_inst.timer_s1.counter_24_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33336\,
            in1 => \N__32554\,
            in2 => \_gnd_net_\,
            in3 => \N__32538\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_12_22_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__47308\,
            ce => \N__32412\,
            sr => \N__46930\
        );

    \current_shift_inst.timer_s1.counter_25_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33340\,
            in1 => \N__32524\,
            in2 => \_gnd_net_\,
            in3 => \N__32508\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__47308\,
            ce => \N__32412\,
            sr => \N__46930\
        );

    \current_shift_inst.timer_s1.counter_26_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33337\,
            in1 => \N__32492\,
            in2 => \_gnd_net_\,
            in3 => \N__32478\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__47308\,
            ce => \N__32412\,
            sr => \N__46930\
        );

    \current_shift_inst.timer_s1.counter_27_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33341\,
            in1 => \N__32473\,
            in2 => \_gnd_net_\,
            in3 => \N__32457\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__47308\,
            ce => \N__32412\,
            sr => \N__46930\
        );

    \current_shift_inst.timer_s1.counter_28_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33338\,
            in1 => \N__32450\,
            in2 => \_gnd_net_\,
            in3 => \N__32436\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__47308\,
            ce => \N__32412\,
            sr => \N__46930\
        );

    \current_shift_inst.timer_s1.counter_29_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__32426\,
            in1 => \N__33339\,
            in2 => \_gnd_net_\,
            in3 => \N__32433\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47308\,
            ce => \N__32412\,
            sr => \N__46930\
        );

    \current_shift_inst.timer_phase.running_RNIC90O_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33666\,
            in2 => \_gnd_net_\,
            in3 => \N__33744\,
            lcout => \current_shift_inst.timer_phase.N_188_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_12_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32640\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32616\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32598\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47420\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__32745\,
            in1 => \N__36229\,
            in2 => \N__34017\,
            in3 => \N__32867\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47413\,
            ce => 'H',
            sr => \N__46813\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__32864\,
            in1 => \N__32749\,
            in2 => \N__36245\,
            in3 => \N__33993\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47413\,
            ce => 'H',
            sr => \N__46813\
        );

    \delay_measurement_inst.delay_hc_reg_31_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__41879\,
            in1 => \N__40798\,
            in2 => \N__37841\,
            in3 => \N__39041\,
            lcout => measured_delay_hc_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47413\,
            ce => 'H',
            sr => \N__46813\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__32861\,
            in1 => \N__32746\,
            in2 => \N__36242\,
            in3 => \N__33792\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47413\,
            ce => 'H',
            sr => \N__46813\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__32744\,
            in1 => \N__36228\,
            in2 => \N__33756\,
            in3 => \N__32866\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47413\,
            ce => 'H',
            sr => \N__46813\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__32862\,
            in1 => \N__32747\,
            in2 => \N__36243\,
            in3 => \N__34059\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47413\,
            ce => 'H',
            sr => \N__46813\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__32743\,
            in1 => \N__36227\,
            in2 => \N__34128\,
            in3 => \N__32865\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47413\,
            ce => 'H',
            sr => \N__46813\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__32863\,
            in1 => \N__32748\,
            in2 => \N__36244\,
            in3 => \N__34038\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47413\,
            ce => 'H',
            sr => \N__46813\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__32736\,
            in1 => \N__32871\,
            in2 => \N__36234\,
            in3 => \N__34218\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47404\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__32868\,
            in1 => \N__36197\,
            in2 => \N__33921\,
            in3 => \N__32740\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47404\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__32737\,
            in1 => \N__32872\,
            in2 => \N__36235\,
            in3 => \N__34197\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47404\,
            ce => 'H',
            sr => \N__46818\
        );

    \delay_measurement_inst.delay_hc_reg_6_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__40808\,
            in1 => \N__41259\,
            in2 => \N__36956\,
            in3 => \N__40916\,
            lcout => measured_delay_hc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47404\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__32739\,
            in1 => \N__32874\,
            in2 => \N__36237\,
            in3 => \N__33942\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47404\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__32869\,
            in1 => \N__36198\,
            in2 => \N__34242\,
            in3 => \N__32741\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47404\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__32738\,
            in1 => \N__32873\,
            in2 => \N__36236\,
            in3 => \N__34176\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47404\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__32870\,
            in1 => \N__36199\,
            in2 => \N__34155\,
            in3 => \N__32742\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47404\,
            ce => 'H',
            sr => \N__46818\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100010001100"
        )
    port map (
            in0 => \N__32730\,
            in1 => \N__34083\,
            in2 => \N__36239\,
            in3 => \N__32860\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47395\,
            ce => 'H',
            sr => \N__46822\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__32856\,
            in1 => \N__36200\,
            in2 => \N__32761\,
            in3 => \N__34332\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47395\,
            ce => 'H',
            sr => \N__46822\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__32857\,
            in1 => \N__36201\,
            in2 => \N__32762\,
            in3 => \N__32901\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47395\,
            ce => 'H',
            sr => \N__46822\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__32729\,
            in1 => \N__32859\,
            in2 => \N__36238\,
            in3 => \N__34104\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47395\,
            ce => 'H',
            sr => \N__46822\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__32858\,
            in1 => \N__36202\,
            in2 => \N__32763\,
            in3 => \N__33969\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47395\,
            ce => 'H',
            sr => \N__46822\
        );

    \delay_measurement_inst.delay_hc_reg_25_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__41637\,
            in1 => \N__40822\,
            in2 => \N__32894\,
            in3 => \N__40622\,
            lcout => measured_delay_hc_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47395\,
            ce => 'H',
            sr => \N__46822\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_0_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__32855\,
            in1 => \N__32731\,
            in2 => \N__36240\,
            in3 => \N__34581\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47385\,
            ce => \N__34781\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34626\,
            in2 => \_gnd_net_\,
            in3 => \N__34579\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34580\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34627\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__47686\,
            in1 => \N__47514\,
            in2 => \N__47940\,
            in3 => \N__45968\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47385\,
            ce => \N__34781\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_1_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__45969\,
            in1 => \N__47932\,
            in2 => \N__47535\,
            in3 => \N__47687\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47385\,
            ce => \N__34781\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__44819\,
            in1 => \N__44622\,
            in2 => \N__42231\,
            in3 => \N__44696\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47385\,
            ce => \N__34781\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__44621\,
            in1 => \N__42226\,
            in2 => \N__44729\,
            in3 => \N__44820\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47385\,
            ce => \N__34781\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_26_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__41961\,
            in1 => \N__40821\,
            in2 => \N__32967\,
            in3 => \N__40639\,
            lcout => measured_delay_hc_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47378\,
            ce => 'H',
            sr => \N__46833\
        );

    \phase_controller_inst1.state_3_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__34553\,
            in1 => \N__34656\,
            in2 => \N__34522\,
            in3 => \N__42029\,
            lcout => \phase_controller_inst1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47378\,
            ce => 'H',
            sr => \N__46833\
        );

    \delay_measurement_inst.delay_hc_reg_7_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__40640\,
            in1 => \N__40823\,
            in2 => \N__37233\,
            in3 => \N__41220\,
            lcout => measured_delay_hc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47378\,
            ce => 'H',
            sr => \N__46833\
        );

    \phase_controller_inst1.state_4_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35037\,
            in2 => \_gnd_net_\,
            in3 => \N__42055\,
            lcout => \phase_controller_inst1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47378\,
            ce => 'H',
            sr => \N__46833\
        );

    \delay_measurement_inst.delay_hc_reg_24_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__32948\,
            in1 => \N__40820\,
            in2 => \N__41894\,
            in3 => \N__39015\,
            lcout => measured_delay_hc_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47378\,
            ce => 'H',
            sr => \N__46833\
        );

    \phase_controller_inst1.S1_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34514\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47373\,
            ce => 'H',
            sr => \N__46841\
        );

    \phase_controller_inst1.state_0_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__42009\,
            in1 => \N__34683\,
            in2 => \N__34730\,
            in3 => \N__33044\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47373\,
            ce => 'H',
            sr => \N__46841\
        );

    \current_shift_inst.timer_s1.running_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__33154\,
            in1 => \N__33369\,
            in2 => \_gnd_net_\,
            in3 => \N__33116\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47373\,
            ce => 'H',
            sr => \N__46841\
        );

    \delay_measurement_inst.start_timer_hc_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__33088\,
            in1 => \N__33072\,
            in2 => \_gnd_net_\,
            in3 => \N__34287\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47365\,
            ce => 'H',
            sr => \N__46844\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42007\,
            in2 => \_gnd_net_\,
            in3 => \N__33040\,
            lcout => \phase_controller_inst1.N_231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.T01_sbtinv_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__42008\,
            in1 => \N__34729\,
            in2 => \N__34526\,
            in3 => \N__33045\,
            lcout => \phase_controller_inst1.N_221_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_sync1_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33000\,
            lcout => \current_shift_inst.S3_syncZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__42115\,
            in1 => \N__44821\,
            in2 => \_gnd_net_\,
            in3 => \N__44707\,
            lcout => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_hc_RNO_0_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34876\,
            in2 => \_gnd_net_\,
            in3 => \N__34857\,
            lcout => \phase_controller_slave.N_214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_sync0_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34819\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.S3_syncZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32994\,
            lcout => \current_shift_inst.un4_control_input_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32973\,
            lcout => \current_shift_inst.un4_control_input_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33408\,
            lcout => \current_shift_inst.un4_control_input_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33390\,
            lcout => \current_shift_inst.un4_control_input_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33372\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33213\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45660\,
            in2 => \_gnd_net_\,
            in3 => \N__45363\,
            lcout => \phase_controller_slave.stoper_tr.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__47900\,
            in1 => \N__47725\,
            in2 => \_gnd_net_\,
            in3 => \N__47542\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33192\,
            lcout => \current_shift_inst.un4_control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33174\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33510\,
            lcout => \current_shift_inst.un4_control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33492\,
            lcout => \current_shift_inst.un4_control_input_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__42680\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43156\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47334\,
            ce => \N__43046\,
            sr => \N__46882\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43157\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42647\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47334\,
            ce => \N__43046\,
            sr => \N__46882\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43158\,
            in2 => \_gnd_net_\,
            in3 => \N__42611\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47334\,
            ce => \N__43046\,
            sr => \N__46882\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33474\,
            lcout => \current_shift_inst.un4_control_input_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33456\,
            lcout => \current_shift_inst.un4_control_input_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33438\,
            lcout => \current_shift_inst.un4_control_input_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46984\,
            in2 => \_gnd_net_\,
            in3 => \N__39602\,
            lcout => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__35627\,
            in1 => \N__33525\,
            in2 => \N__38075\,
            in3 => \N__33584\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_15_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__39669\,
            in1 => \N__33900\,
            in2 => \N__33540\,
            in3 => \N__35237\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_321_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__35238\,
            in1 => \N__36433\,
            in2 => \N__33537\,
            in3 => \N__33531\,
            lcout => \delay_measurement_inst.un3_elapsed_time_tr_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__33585\,
            in1 => \N__35942\,
            in2 => \N__33519\,
            in3 => \N__35970\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI61PC3_6_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__33555\,
            in1 => \N__35750\,
            in2 => \N__33534\,
            in3 => \N__35820\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110100"
        )
    port map (
            in0 => \N__33901\,
            in1 => \N__39670\,
            in2 => \N__35295\,
            in3 => \N__36434\,
            lcout => \delay_measurement_inst.N_284_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__35741\,
            in1 => \N__35639\,
            in2 => \N__35459\,
            in3 => \N__35817\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__38289\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47323\,
            ce => \N__36365\,
            sr => \N__46902\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38262\,
            lcout => \delay_measurement_inst.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47323\,
            ce => \N__36365\,
            sr => \N__46902\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__35906\,
            in1 => \N__35452\,
            in2 => \N__35883\,
            in3 => \N__35626\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35837\,
            in2 => \_gnd_net_\,
            in3 => \N__35435\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_320_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__35966\,
            in1 => \N__35882\,
            in2 => \N__35943\,
            in3 => \N__35907\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_9_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000110001"
        )
    port map (
            in0 => \N__33572\,
            in1 => \N__33870\,
            in2 => \N__35749\,
            in3 => \N__36439\,
            lcout => measured_delay_tr_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47319\,
            ce => \N__35508\,
            sr => \N__46909\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__33554\,
            in1 => \N__33902\,
            in2 => \_gnd_net_\,
            in3 => \N__35290\,
            lcout => \delay_measurement_inst.N_305_1\,
            ltout => \delay_measurement_inst.N_305_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_10_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36437\,
            in2 => \N__33576\,
            in3 => \N__35703\,
            lcout => measured_delay_tr_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47319\,
            ce => \N__35508\,
            sr => \N__46909\
        );

    \delay_measurement_inst.delay_tr_reg_esr_11_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010101000"
        )
    port map (
            in0 => \N__35688\,
            in1 => \N__33567\,
            in2 => \N__36454\,
            in3 => \_gnd_net_\,
            lcout => measured_delay_tr_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47319\,
            ce => \N__35508\,
            sr => \N__46909\
        );

    \delay_measurement_inst.delay_tr_reg_esr_12_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36438\,
            in2 => \N__33573\,
            in3 => \N__35667\,
            lcout => measured_delay_tr_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47319\,
            ce => \N__35508\,
            sr => \N__46909\
        );

    \delay_measurement_inst.delay_tr_reg_esr_13_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010101000"
        )
    port map (
            in0 => \N__36003\,
            in1 => \N__33571\,
            in2 => \N__36455\,
            in3 => \_gnd_net_\,
            lcout => measured_delay_tr_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47319\,
            ce => \N__35508\,
            sr => \N__46909\
        );

    \delay_measurement_inst.delay_tr_reg_esr_19_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__36432\,
            in1 => \N__35878\,
            in2 => \_gnd_net_\,
            in3 => \N__35288\,
            lcout => measured_delay_tr_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47316\,
            ce => \N__35507\,
            sr => \N__46915\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUIS_14_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39643\,
            in2 => \_gnd_net_\,
            in3 => \N__38056\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33591\,
            in1 => \N__33597\,
            in2 => \N__35856\,
            in3 => \N__33879\,
            lcout => \delay_measurement_inst.N_358\,
            ltout => \delay_measurement_inst.N_358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_16_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36430\,
            in2 => \N__33747\,
            in3 => \N__35965\,
            lcout => measured_delay_tr_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47313\,
            ce => \N__35509\,
            sr => \N__46922\
        );

    \delay_measurement_inst.delay_tr_reg_esr_17_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__36429\,
            in1 => \N__35932\,
            in2 => \_gnd_net_\,
            in3 => \N__35287\,
            lcout => measured_delay_tr_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47313\,
            ce => \N__35509\,
            sr => \N__46922\
        );

    \delay_measurement_inst.delay_tr_reg_esr_18_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__35286\,
            in1 => \N__36431\,
            in2 => \_gnd_net_\,
            in3 => \N__35900\,
            lcout => measured_delay_tr_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47313\,
            ce => \N__35509\,
            sr => \N__46922\
        );

    \current_shift_inst.timer_phase.running_RNIL91O_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__33742\,
            in1 => \N__33701\,
            in2 => \_gnd_net_\,
            in3 => \N__33675\,
            lcout => \current_shift_inst.timer_phase.N_192_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36033\,
            in1 => \N__36042\,
            in2 => \N__36024\,
            in3 => \N__36051\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35343\,
            in2 => \_gnd_net_\,
            in3 => \N__39981\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_337_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36072\,
            in1 => \N__36081\,
            in2 => \N__36063\,
            in3 => \N__35844\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_14_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__35745\,
            in1 => \N__38062\,
            in2 => \_gnd_net_\,
            in3 => \N__35591\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_293_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2EEG9_15_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011100"
        )
    port map (
            in0 => \N__39653\,
            in1 => \N__33909\,
            in2 => \N__33882\,
            in3 => \N__35285\,
            lcout => \delay_measurement_inst.N_324\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36468\,
            in2 => \_gnd_net_\,
            in3 => \N__36012\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__35592\,
            in1 => \N__39671\,
            in2 => \N__35751\,
            in3 => \N__35294\,
            lcout => \delay_measurement_inst.N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S2_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34734\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47307\,
            ce => 'H',
            sr => \N__46945\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40954\,
            in2 => \_gnd_net_\,
            in3 => \N__43000\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_335_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34527\,
            in2 => \_gnd_net_\,
            in3 => \N__34546\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33840\,
            in2 => \N__33828\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_5_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33804\,
            in2 => \_gnd_net_\,
            in3 => \N__33786\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33783\,
            in2 => \N__33771\,
            in3 => \N__34074\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34071\,
            in2 => \_gnd_net_\,
            in3 => \N__34053\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34050\,
            in2 => \_gnd_net_\,
            in3 => \N__34032\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34029\,
            in2 => \_gnd_net_\,
            in3 => \N__34008\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34005\,
            in2 => \_gnd_net_\,
            in3 => \N__33987\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33984\,
            in2 => \_gnd_net_\,
            in3 => \N__33957\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33954\,
            in2 => \_gnd_net_\,
            in3 => \N__33936\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33933\,
            in2 => \_gnd_net_\,
            in3 => \N__33912\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34254\,
            in2 => \_gnd_net_\,
            in3 => \N__34233\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34230\,
            in2 => \_gnd_net_\,
            in3 => \N__34212\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34209\,
            in2 => \_gnd_net_\,
            in3 => \N__34191\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34188\,
            in2 => \_gnd_net_\,
            in3 => \N__34170\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34167\,
            in2 => \_gnd_net_\,
            in3 => \N__34146\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34142\,
            in2 => \_gnd_net_\,
            in3 => \N__34119\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34116\,
            in2 => \_gnd_net_\,
            in3 => \N__34098\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34095\,
            in2 => \_gnd_net_\,
            in3 => \N__34077\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34347\,
            in2 => \_gnd_net_\,
            in3 => \N__34335\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m2_e_2_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36857\,
            in2 => \_gnd_net_\,
            in3 => \N__40878\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m3_0_a3_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__37037\,
            in1 => \N__36938\,
            in2 => \N__34326\,
            in3 => \N__34311\,
            lcout => \phase_controller_inst1.stoper_hc.un1_N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__39006\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41824\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto31_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m2_e_3_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36826\,
            in1 => \N__36899\,
            in2 => \N__37739\,
            in3 => \N__36978\,
            lcout => \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34473\,
            in2 => \_gnd_net_\,
            in3 => \N__34449\,
            lcout => \phase_controller_inst1.N_228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m3_0_1_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36590\,
            in1 => \N__36630\,
            in2 => \N__37550\,
            in3 => \N__36683\,
            lcout => \phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC2_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41004\,
            lcout => delay_hc_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47405\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41853\,
            in2 => \_gnd_net_\,
            in3 => \N__39005\,
            lcout => \delay_measurement_inst.delay_hc_reg3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_1_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__34681\,
            in1 => \N__34451\,
            in2 => \N__34725\,
            in3 => \N__34476\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47396\,
            ce => 'H',
            sr => \N__46823\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__34475\,
            in1 => \N__34638\,
            in2 => \N__34605\,
            in3 => \N__34590\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47396\,
            ce => 'H',
            sr => \N__46823\
        );

    \delay_measurement_inst.delay_hc_reg_14_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111010111010"
        )
    port map (
            in0 => \N__40618\,
            in1 => \N__40811\,
            in2 => \N__36750\,
            in3 => \N__41496\,
            lcout => measured_delay_hc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47396\,
            ce => 'H',
            sr => \N__46823\
        );

    \delay_measurement_inst.delay_hc_reg_13_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__40809\,
            in1 => \N__41523\,
            in2 => \N__37560\,
            in3 => \N__40617\,
            lcout => measured_delay_hc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47396\,
            ce => 'H',
            sr => \N__46823\
        );

    \delay_measurement_inst.prev_tr_sig_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36303\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.prev_tr_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47396\,
            ce => 'H',
            sr => \N__46823\
        );

    \delay_measurement_inst.delay_hc_reg_18_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__40810\,
            in1 => \N__41730\,
            in2 => \N__34426\,
            in3 => \N__40619\,
            lcout => measured_delay_hc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47396\,
            ce => 'H',
            sr => \N__46823\
        );

    \phase_controller_inst1.state_2_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__34554\,
            in1 => \N__34450\,
            in2 => \N__34521\,
            in3 => \N__34474\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47396\,
            ce => 'H',
            sr => \N__46823\
        );

    \phase_controller_slave.stoper_hc.target_time_18_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000000010000"
        )
    port map (
            in0 => \N__34383\,
            in1 => \N__37865\,
            in2 => \N__37439\,
            in3 => \N__34415\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47386\,
            ce => \N__37091\,
            sr => \N__46828\
        );

    \phase_controller_slave.stoper_hc.target_time_12_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36607\,
            in1 => \N__37186\,
            in2 => \N__37440\,
            in3 => \N__37495\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47386\,
            ce => \N__37091\,
            sr => \N__46828\
        );

    \phase_controller_slave.stoper_hc.target_time_17_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001100"
        )
    port map (
            in0 => \N__36500\,
            in1 => \N__37429\,
            in2 => \N__37883\,
            in3 => \N__34382\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47386\,
            ce => \N__37091\,
            sr => \N__46828\
        );

    \reset_ibuf_gb_io_RNI79U7_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46977\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => red_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34718\,
            in2 => \_gnd_net_\,
            in3 => \N__34682\,
            lcout => \phase_controller_inst1.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__42130\,
            in1 => \N__44822\,
            in2 => \_gnd_net_\,
            in3 => \N__44708\,
            lcout => \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_RNO_0_3_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35054\,
            in2 => \_gnd_net_\,
            in3 => \N__42054\,
            lcout => \phase_controller_inst1.N_232\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.target_time_9_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__37411\,
            in1 => \N__37042\,
            in2 => \_gnd_net_\,
            in3 => \N__37690\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47374\,
            ce => \N__37099\,
            sr => \N__46842\
        );

    \phase_controller_slave.stoper_hc.target_time_19_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__37691\,
            in1 => \N__37881\,
            in2 => \_gnd_net_\,
            in3 => \N__36558\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47374\,
            ce => \N__37099\,
            sr => \N__46842\
        );

    \phase_controller_slave.start_timer_hc_RNO_1_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35161\,
            in2 => \_gnd_net_\,
            in3 => \N__35197\,
            lcout => \phase_controller_slave.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.state_2_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__35198\,
            in1 => \N__34877\,
            in2 => \N__35166\,
            in3 => \N__34858\,
            lcout => \phase_controller_slave.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47366\,
            ce => 'H',
            sr => \N__46845\
        );

    \phase_controller_slave.stoper_hc.time_passed_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__34859\,
            in1 => \N__44649\,
            in2 => \N__34650\,
            in3 => \N__44620\,
            lcout => \phase_controller_slave.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47366\,
            ce => 'H',
            sr => \N__46845\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_13_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__44873\,
            in1 => \N__42129\,
            in2 => \N__44772\,
            in3 => \N__44406\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47366\,
            ce => 'H',
            sr => \N__46845\
        );

    \phase_controller_slave.start_timer_hc_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__34942\,
            in1 => \N__34914\,
            in2 => \N__42192\,
            in3 => \N__34908\,
            lcout => \phase_controller_slave.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47358\,
            ce => 'H',
            sr => \N__46853\
        );

    \phase_controller_slave.S2_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__34974\,
            in1 => \N__35157\,
            in2 => \N__34895\,
            in3 => \N__35406\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47358\,
            ce => 'H',
            sr => \N__46853\
        );

    \phase_controller_slave.state_1_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__35385\,
            in1 => \N__34878\,
            in2 => \N__35412\,
            in3 => \N__34860\,
            lcout => \phase_controller_slave.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47358\,
            ce => 'H',
            sr => \N__46853\
        );

    \phase_controller_slave.S1_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__34973\,
            in1 => \_gnd_net_\,
            in2 => \N__34823\,
            in3 => \N__35156\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47358\,
            ce => 'H',
            sr => \N__46853\
        );

    \phase_controller_slave.state_4_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__35055\,
            in1 => \N__34972\,
            in2 => \_gnd_net_\,
            in3 => \N__34941\,
            lcout => \phase_controller_slave.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47358\,
            ce => 'H',
            sr => \N__46853\
        );

    \delay_measurement_inst.start_timer_tr_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__36291\,
            in1 => \N__35132\,
            in2 => \_gnd_net_\,
            in3 => \N__35101\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47358\,
            ce => 'H',
            sr => \N__46853\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__35339\,
            in1 => \N__35312\,
            in2 => \_gnd_net_\,
            in3 => \N__39976\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47358\,
            ce => 'H',
            sr => \N__46853\
        );

    \phase_controller_slave.state_RNIVDE2_0_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35218\,
            in2 => \_gnd_net_\,
            in3 => \N__35207\,
            lcout => \phase_controller_slave.N_211\,
            ltout => \phase_controller_slave.N_211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_tr_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__45533\,
            in1 => \N__35352\,
            in2 => \N__34800\,
            in3 => \N__34943\,
            lcout => \phase_controller_slave.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47351\,
            ce => 'H',
            sr => \N__46862\
        );

    \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__45495\,
            in1 => \N__45730\,
            in2 => \_gnd_net_\,
            in3 => \N__45411\,
            lcout => OPEN,
            ltout => \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.time_passed_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__35222\,
            in1 => \N__39528\,
            in2 => \N__35226\,
            in3 => \N__41091\,
            lcout => \phase_controller_slave.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47351\,
            ce => 'H',
            sr => \N__46862\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_16_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45723\,
            in1 => \N__45412\,
            in2 => \N__45534\,
            in3 => \N__37980\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47351\,
            ce => 'H',
            sr => \N__46862\
        );

    \phase_controller_slave.state_0_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__35208\,
            in1 => \N__35410\,
            in2 => \N__35223\,
            in3 => \N__35384\,
            lcout => \phase_controller_slave.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47351\,
            ce => 'H',
            sr => \N__46862\
        );

    \phase_controller_slave.state_3_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__34920\,
            in1 => \N__35199\,
            in2 => \N__35165\,
            in3 => \N__35172\,
            lcout => \phase_controller_slave.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47351\,
            ce => 'H',
            sr => \N__46862\
        );

    \delay_measurement_inst.stop_timer_tr_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__36301\,
            in1 => \N__35133\,
            in2 => \N__46989\,
            in3 => \N__35102\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.state_RNO_0_3_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__35065\,
            in1 => \N__34971\,
            in2 => \_gnd_net_\,
            in3 => \N__34944\,
            lcout => \phase_controller_slave.N_213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__43259\,
            in1 => \N__46214\,
            in2 => \_gnd_net_\,
            in3 => \N__46174\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43328\,
            in2 => \N__35415\,
            in3 => \N__42739\,
            lcout => \phase_controller_inst1.stoper_tr.N_20_li\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_tr_RNO_0_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35411\,
            in2 => \_gnd_net_\,
            in3 => \N__35383\,
            lcout => \phase_controller_slave.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__35332\,
            in1 => \N__35313\,
            in2 => \_gnd_net_\,
            in3 => \N__39972\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_338_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42646\,
            in1 => \N__42679\,
            in2 => \N__42612\,
            in3 => \N__43105\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110101"
        )
    port map (
            in0 => \N__42893\,
            in1 => \N__46255\,
            in2 => \N__35298\,
            in3 => \N__43258\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_5_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__35607\,
            in1 => \N__36448\,
            in2 => \N__35563\,
            in3 => \N__35838\,
            lcout => measured_delay_tr_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47328\,
            ce => \N__35510\,
            sr => \N__46889\
        );

    \delay_measurement_inst.delay_tr_reg_ess_3_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__36447\,
            in1 => \N__35610\,
            in2 => \N__35460\,
            in3 => \N__35557\,
            lcout => measured_delay_tr_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47328\,
            ce => \N__35510\,
            sr => \N__46889\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__35790\,
            in1 => \N__35576\,
            in2 => \N__35772\,
            in3 => \N__35289\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_331\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI80KG7_6_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39665\,
            in2 => \N__35229\,
            in3 => \N__35818\,
            lcout => \delay_measurement_inst.N_333\,
            ltout => \delay_measurement_inst.N_333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_4_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__35549\,
            in1 => \N__35436\,
            in2 => \N__35643\,
            in3 => \N__36452\,
            lcout => measured_delay_tr_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47328\,
            ce => \N__35510\,
            sr => \N__46889\
        );

    \delay_measurement_inst.delay_tr_reg_esr_6_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000001"
        )
    port map (
            in0 => \N__36446\,
            in1 => \N__35608\,
            in2 => \N__35565\,
            in3 => \N__35819\,
            lcout => measured_delay_tr_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47328\,
            ce => \N__35510\,
            sr => \N__46889\
        );

    \delay_measurement_inst.delay_tr_reg_ess_1_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__35609\,
            in1 => \N__35640\,
            in2 => \N__35564\,
            in3 => \N__36453\,
            lcout => measured_delay_tr_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47328\,
            ce => \N__35510\,
            sr => \N__46889\
        );

    \delay_measurement_inst.delay_tr_reg_esr_2_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__35628\,
            in1 => \N__35550\,
            in2 => \N__36456\,
            in3 => \N__35606\,
            lcout => measured_delay_tr_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47328\,
            ce => \N__35510\,
            sr => \N__46889\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35663\,
            in1 => \N__35687\,
            in2 => \N__36002\,
            in3 => \N__35702\,
            lcout => \delay_measurement_inst.N_328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_7_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__36435\,
            in1 => \N__35561\,
            in2 => \_gnd_net_\,
            in3 => \N__35789\,
            lcout => measured_delay_tr_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47324\,
            ce => \N__35511\,
            sr => \N__46903\
        );

    \delay_measurement_inst.delay_tr_reg_esr_8_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__36436\,
            in1 => \N__35562\,
            in2 => \_gnd_net_\,
            in3 => \N__35768\,
            lcout => measured_delay_tr_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47324\,
            ce => \N__35511\,
            sr => \N__46903\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__39574\,
            in1 => \N__42493\,
            in2 => \_gnd_net_\,
            in3 => \N__42844\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38282\,
            in2 => \N__38235\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__47320\,
            ce => \N__36366\,
            sr => \N__46910\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38255\,
            in2 => \N__38211\,
            in3 => \N__35418\,
            lcout => \delay_measurement_inst.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__47320\,
            ce => \N__36366\,
            sr => \N__46910\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38234\,
            in2 => \N__38187\,
            in3 => \N__35823\,
            lcout => \delay_measurement_inst.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__47320\,
            ce => \N__36366\,
            sr => \N__46910\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38210\,
            in2 => \N__38163\,
            in3 => \N__35793\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__47320\,
            ce => \N__36366\,
            sr => \N__46910\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38186\,
            in2 => \N__38139\,
            in3 => \N__35775\,
            lcout => \delay_measurement_inst.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__47320\,
            ce => \N__36366\,
            sr => \N__46910\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38162\,
            in2 => \N__38505\,
            in3 => \N__35754\,
            lcout => \delay_measurement_inst.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__47320\,
            ce => \N__36366\,
            sr => \N__46910\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38138\,
            in2 => \N__38481\,
            in3 => \N__35706\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__47320\,
            ce => \N__36366\,
            sr => \N__46910\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38504\,
            in2 => \N__38457\,
            in3 => \N__35691\,
            lcout => \delay_measurement_inst.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__47320\,
            ce => \N__36366\,
            sr => \N__46910\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38480\,
            in2 => \N__38433\,
            in3 => \N__35670\,
            lcout => \delay_measurement_inst.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__47317\,
            ce => \N__36347\,
            sr => \N__46916\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38456\,
            in2 => \N__38409\,
            in3 => \N__35646\,
            lcout => \delay_measurement_inst.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__47317\,
            ce => \N__36347\,
            sr => \N__46916\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38432\,
            in2 => \N__38385\,
            in3 => \N__35979\,
            lcout => \delay_measurement_inst.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__47317\,
            ce => \N__36347\,
            sr => \N__46916\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38408\,
            in2 => \N__38361\,
            in3 => \N__35976\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__47317\,
            ce => \N__36347\,
            sr => \N__46916\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38384\,
            in2 => \N__38337\,
            in3 => \N__35973\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__47317\,
            ce => \N__36347\,
            sr => \N__46916\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38360\,
            in2 => \N__38313\,
            in3 => \N__35946\,
            lcout => \delay_measurement_inst.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__47317\,
            ce => \N__36347\,
            sr => \N__46916\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38336\,
            in2 => \N__38697\,
            in3 => \N__35910\,
            lcout => \delay_measurement_inst.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__47317\,
            ce => \N__36347\,
            sr => \N__46916\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38312\,
            in2 => \N__38673\,
            in3 => \N__35886\,
            lcout => \delay_measurement_inst.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__47317\,
            ce => \N__36347\,
            sr => \N__46916\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38696\,
            in2 => \N__38649\,
            in3 => \N__35859\,
            lcout => \delay_measurement_inst.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__47314\,
            ce => \N__36355\,
            sr => \N__46923\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38672\,
            in2 => \N__38625\,
            in3 => \N__35847\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__47314\,
            ce => \N__36355\,
            sr => \N__46923\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38648\,
            in2 => \N__38601\,
            in3 => \N__36084\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__47314\,
            ce => \N__36355\,
            sr => \N__46923\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38624\,
            in2 => \N__38577\,
            in3 => \N__36075\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__47314\,
            ce => \N__36355\,
            sr => \N__46923\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38600\,
            in2 => \N__38553\,
            in3 => \N__36066\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__47314\,
            ce => \N__36355\,
            sr => \N__46923\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38576\,
            in2 => \N__38529\,
            in3 => \N__36054\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__47314\,
            ce => \N__36355\,
            sr => \N__46923\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38552\,
            in2 => \N__38871\,
            in3 => \N__36045\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__47314\,
            ce => \N__36355\,
            sr => \N__46923\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38528\,
            in2 => \N__38847\,
            in3 => \N__36036\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__47314\,
            ce => \N__36355\,
            sr => \N__46923\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38870\,
            in2 => \N__38823\,
            in3 => \N__36027\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__47311\,
            ce => \N__36348\,
            sr => \N__46926\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38846\,
            in2 => \N__38799\,
            in3 => \N__36015\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__47311\,
            ce => \N__36348\,
            sr => \N__46926\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38822\,
            in2 => \N__38775\,
            in3 => \N__36006\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__47311\,
            ce => \N__36348\,
            sr => \N__46926\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38798\,
            in2 => \N__38754\,
            in3 => \N__36462\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__47311\,
            ce => \N__36348\,
            sr => \N__46926\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36459\,
            lcout => \delay_measurement_inst.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47311\,
            ce => \N__36348\,
            sr => \N__46926\
        );

    \SB_DFF_inst_DELAY_TR1_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36318\,
            lcout => delay_tr_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47443\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR2_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36309\,
            lcout => delay_tr_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47443\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__36261\,
            in1 => \N__42072\,
            in2 => \N__36178\,
            in3 => \N__36255\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47436\,
            ce => 'H',
            sr => \N__46804\
        );

    \delay_measurement_inst.delay_hc_reg_0_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__40784\,
            in1 => \N__36985\,
            in2 => \N__41899\,
            in3 => \N__39030\,
            lcout => measured_delay_hc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47428\,
            ce => 'H',
            sr => \N__46807\
        );

    \delay_measurement_inst.delay_hc_reg_3_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__36867\,
            in1 => \N__40786\,
            in2 => \N__41346\,
            in3 => \N__40912\,
            lcout => measured_delay_hc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47428\,
            ce => 'H',
            sr => \N__46807\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__40989\,
            in1 => \N__40958\,
            in2 => \_gnd_net_\,
            in3 => \N__42999\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47428\,
            ce => 'H',
            sr => \N__46807\
        );

    \delay_measurement_inst.delay_hc_reg_1_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__36909\,
            in1 => \N__40785\,
            in2 => \N__41388\,
            in3 => \N__40911\,
            lcout => measured_delay_hc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47428\,
            ce => 'H',
            sr => \N__46807\
        );

    \delay_measurement_inst.delay_hc_reg_5_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__40743\,
            in1 => \N__41289\,
            in2 => \N__37747\,
            in3 => \N__40630\,
            lcout => measured_delay_hc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47421\,
            ce => 'H',
            sr => \N__46810\
        );

    \delay_measurement_inst.delay_hc_reg_11_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__40742\,
            in1 => \N__41583\,
            in2 => \N__36648\,
            in3 => \N__40628\,
            lcout => measured_delay_hc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47421\,
            ce => 'H',
            sr => \N__46810\
        );

    \delay_measurement_inst.delay_hc_reg_12_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__40629\,
            in1 => \N__40744\,
            in2 => \N__36608\,
            in3 => \N__41553\,
            lcout => measured_delay_hc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47421\,
            ce => 'H',
            sr => \N__46810\
        );

    \delay_measurement_inst.delay_hc_reg_19_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__40775\,
            in1 => \N__41709\,
            in2 => \N__36551\,
            in3 => \N__40620\,
            lcout => measured_delay_hc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47414\,
            ce => 'H',
            sr => \N__46814\
        );

    \delay_measurement_inst.delay_hc_reg_8_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__40621\,
            in1 => \N__40776\,
            in2 => \N__37932\,
            in3 => \N__41187\,
            lcout => measured_delay_hc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47414\,
            ce => 'H',
            sr => \N__46814\
        );

    \delay_measurement_inst.delay_hc_reg_4_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__36825\,
            in1 => \N__40777\,
            in2 => \N__41319\,
            in3 => \N__40626\,
            lcout => measured_delay_hc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47406\,
            ce => 'H',
            sr => \N__46819\
        );

    \delay_measurement_inst.delay_hc_reg_17_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111010101110"
        )
    port map (
            in0 => \N__40625\,
            in1 => \N__36501\,
            in2 => \N__40819\,
            in3 => \N__41409\,
            lcout => measured_delay_hc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47406\,
            ce => 'H',
            sr => \N__46819\
        );

    \delay_measurement_inst.delay_hc_reg_10_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__36693\,
            in1 => \N__41613\,
            in2 => \N__40832\,
            in3 => \N__40623\,
            lcout => measured_delay_hc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47406\,
            ce => 'H',
            sr => \N__46819\
        );

    \delay_measurement_inst.delay_hc_reg_16_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111010101110"
        )
    port map (
            in0 => \N__40624\,
            in1 => \N__36775\,
            in2 => \N__40818\,
            in3 => \N__41433\,
            lcout => measured_delay_hc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47406\,
            ce => 'H',
            sr => \N__46819\
        );

    \delay_measurement_inst.delay_hc_reg_9_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001010"
        )
    port map (
            in0 => \N__37036\,
            in1 => \N__41154\,
            in2 => \N__40833\,
            in3 => \N__40627\,
            lcout => measured_delay_hc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47406\,
            ce => 'H',
            sr => \N__46819\
        );

    \phase_controller_slave.stoper_hc.target_time_0_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37187\,
            in1 => \N__37508\,
            in2 => \N__36993\,
            in3 => \N__37428\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47397\,
            ce => \N__37106\,
            sr => \N__46824\
        );

    \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__37421\,
            in1 => \N__36957\,
            in2 => \_gnd_net_\,
            in3 => \N__37645\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47397\,
            ce => \N__37106\,
            sr => \N__46824\
        );

    \phase_controller_slave.stoper_hc.target_time_1_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__37647\,
            in1 => \N__37423\,
            in2 => \_gnd_net_\,
            in3 => \N__36914\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47397\,
            ce => \N__37106\,
            sr => \N__46824\
        );

    \phase_controller_slave.stoper_hc.target_time_2_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__40885\,
            in1 => \_gnd_net_\,
            in2 => \N__37438\,
            in3 => \N__37648\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47397\,
            ce => \N__37106\,
            sr => \N__46824\
        );

    \phase_controller_slave.stoper_hc.target_time_3_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__37649\,
            in1 => \N__37424\,
            in2 => \_gnd_net_\,
            in3 => \N__36876\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47397\,
            ce => \N__37106\,
            sr => \N__46824\
        );

    \phase_controller_slave.stoper_hc.target_time_4_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__37882\,
            in1 => \N__36824\,
            in2 => \_gnd_net_\,
            in3 => \N__37650\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47397\,
            ce => \N__37106\,
            sr => \N__46824\
        );

    \phase_controller_slave.stoper_hc.target_time_16_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__37422\,
            in1 => \N__36774\,
            in2 => \_gnd_net_\,
            in3 => \N__37646\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47397\,
            ce => \N__37106\,
            sr => \N__46824\
        );

    \phase_controller_slave.stoper_hc.target_time_14_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__36749\,
            in1 => \_gnd_net_\,
            in2 => \N__37436\,
            in3 => \N__37681\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47387\,
            ce => \N__37092\,
            sr => \N__46829\
        );

    \phase_controller_slave.stoper_hc.target_time_10_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36697\,
            in1 => \N__37188\,
            in2 => \N__37437\,
            in3 => \N__37509\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47387\,
            ce => \N__37092\,
            sr => \N__46829\
        );

    \phase_controller_slave.stoper_hc.target_time_8_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__37683\,
            in1 => \N__37887\,
            in2 => \_gnd_net_\,
            in3 => \N__37928\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47387\,
            ce => \N__37092\,
            sr => \N__46829\
        );

    \phase_controller_slave.stoper_hc.target_time_5_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__37886\,
            in1 => \N__37743\,
            in2 => \_gnd_net_\,
            in3 => \N__37682\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47387\,
            ce => \N__37092\,
            sr => \N__46829\
        );

    \phase_controller_slave.stoper_hc.target_time_13_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37510\,
            in1 => \N__37416\,
            in2 => \N__37562\,
            in3 => \N__37190\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47387\,
            ce => \N__37092\,
            sr => \N__46829\
        );

    \phase_controller_slave.stoper_hc.target_time_15_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37412\,
            in1 => \N__37189\,
            in2 => \N__40562\,
            in3 => \N__37511\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47387\,
            ce => \N__37092\,
            sr => \N__46829\
        );

    \phase_controller_slave.stoper_hc.target_time_7_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37512\,
            in1 => \N__37417\,
            in2 => \N__37241\,
            in3 => \N__37191\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47387\,
            ce => \N__37092\,
            sr => \N__46829\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__47721\,
            in1 => \N__47570\,
            in2 => \N__47939\,
            in3 => \N__45060\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47379\,
            ce => 'H',
            sr => \N__46834\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__47569\,
            in1 => \N__47926\,
            in2 => \N__47741\,
            in3 => \N__45021\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47379\,
            ce => 'H',
            sr => \N__46834\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_1_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__44891\,
            in1 => \N__44751\,
            in2 => \N__42230\,
            in3 => \N__39378\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47379\,
            ce => 'H',
            sr => \N__46834\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_11_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__44750\,
            in1 => \N__44892\,
            in2 => \N__44469\,
            in3 => \N__42217\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47379\,
            ce => 'H',
            sr => \N__46834\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39540\,
            in2 => \N__39801\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39762\,
            in2 => \_gnd_net_\,
            in3 => \N__37965\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39504\,
            in2 => \N__39738\,
            in3 => \N__37962\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40296\,
            in2 => \_gnd_net_\,
            in3 => \N__37959\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45315\,
            in2 => \_gnd_net_\,
            in3 => \N__37956\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40257\,
            in2 => \_gnd_net_\,
            in3 => \N__37953\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40232\,
            in2 => \_gnd_net_\,
            in3 => \N__37950\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40196\,
            in2 => \_gnd_net_\,
            in3 => \N__37947\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40175\,
            in2 => \_gnd_net_\,
            in3 => \N__37944\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40154\,
            in2 => \_gnd_net_\,
            in3 => \N__37998\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40133\,
            in2 => \_gnd_net_\,
            in3 => \N__37995\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40484\,
            in2 => \_gnd_net_\,
            in3 => \N__37992\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40464\,
            in2 => \_gnd_net_\,
            in3 => \N__37989\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40431\,
            in2 => \_gnd_net_\,
            in3 => \N__37986\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40395\,
            in2 => \_gnd_net_\,
            in3 => \N__37983\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40367\,
            in2 => \_gnd_net_\,
            in3 => \N__37974\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40340\,
            in2 => \_gnd_net_\,
            in3 => \N__37971\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40316\,
            in2 => \_gnd_net_\,
            in3 => \N__37968\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41114\,
            in2 => \_gnd_net_\,
            in3 => \N__38085\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45738\,
            in1 => \N__45416\,
            in2 => \N__45558\,
            in3 => \N__38082\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47352\,
            ce => 'H',
            sr => \N__46863\
        );

    \delay_measurement_inst.delay_tr_reg_14_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__39698\,
            in1 => \N__38076\,
            in2 => \N__42902\,
            in3 => \N__39614\,
            lcout => measured_delay_tr_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47352\,
            ce => 'H',
            sr => \N__46863\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45739\,
            in1 => \N__45417\,
            in2 => \N__45559\,
            in3 => \N__38040\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47352\,
            ce => 'H',
            sr => \N__46863\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_2_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__45414\,
            in1 => \N__45513\,
            in2 => \N__45752\,
            in3 => \N__38034\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47352\,
            ce => 'H',
            sr => \N__46863\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_3_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__45740\,
            in1 => \N__38025\,
            in2 => \N__45560\,
            in3 => \N__45419\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47352\,
            ce => 'H',
            sr => \N__46863\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_4_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__45415\,
            in1 => \N__45517\,
            in2 => \N__45753\,
            in3 => \N__38016\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47352\,
            ce => 'H',
            sr => \N__46863\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_6_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45741\,
            in1 => \N__45418\,
            in2 => \N__45561\,
            in3 => \N__38007\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47352\,
            ce => 'H',
            sr => \N__46863\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__39534\,
            in1 => \N__39797\,
            in2 => \_gnd_net_\,
            in3 => \N__41074\,
            lcout => OPEN,
            ltout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__45443\,
            in1 => \N__45569\,
            in2 => \N__38115\,
            in3 => \N__45734\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47343\,
            ce => 'H',
            sr => \N__46874\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45732\,
            in1 => \N__45444\,
            in2 => \N__45591\,
            in3 => \N__38112\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47343\,
            ce => 'H',
            sr => \N__46874\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__45442\,
            in1 => \N__45565\,
            in2 => \N__45751\,
            in3 => \N__38103\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47343\,
            ce => 'H',
            sr => \N__46874\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45733\,
            in1 => \N__45445\,
            in2 => \N__45592\,
            in3 => \N__38094\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47343\,
            ce => 'H',
            sr => \N__46874\
        );

    \phase_controller_slave.stoper_tr.target_time_5_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__42799\,
            in1 => \N__43340\,
            in2 => \N__46336\,
            in3 => \N__42752\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47335\,
            ce => \N__43380\,
            sr => \N__46883\
        );

    \phase_controller_slave.stoper_tr.target_time_8_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__42751\,
            in1 => \N__39575\,
            in2 => \_gnd_net_\,
            in3 => \N__43341\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47335\,
            ce => \N__43380\,
            sr => \N__46883\
        );

    \phase_controller_slave.stoper_tr.target_time_3_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__40047\,
            in1 => \N__40010\,
            in2 => \_gnd_net_\,
            in3 => \N__46157\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47335\,
            ce => \N__43380\,
            sr => \N__46883\
        );

    \phase_controller_slave.stoper_tr.target_time_15_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43251\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43342\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47335\,
            ce => \N__43380\,
            sr => \N__46883\
        );

    \phase_controller_slave.stoper_tr.target_time_14_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__43339\,
            in1 => \N__43252\,
            in2 => \_gnd_net_\,
            in3 => \N__42901\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47335\,
            ce => \N__43380\,
            sr => \N__46883\
        );

    \phase_controller_slave.stoper_tr.target_time_1_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__46158\,
            in1 => \N__40083\,
            in2 => \N__40073\,
            in3 => \N__40045\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47335\,
            ce => \N__43380\,
            sr => \N__46883\
        );

    \phase_controller_slave.stoper_tr.target_time_2_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000010001000"
        )
    port map (
            in0 => \N__40046\,
            in1 => \N__40102\,
            in2 => \N__40019\,
            in3 => \N__46156\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47335\,
            ce => \N__43380\,
            sr => \N__46883\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39939\,
            in1 => \N__38281\,
            in2 => \_gnd_net_\,
            in3 => \N__38265\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__47329\,
            ce => \N__38732\,
            sr => \N__46890\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39935\,
            in1 => \N__38254\,
            in2 => \_gnd_net_\,
            in3 => \N__38238\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__47329\,
            ce => \N__38732\,
            sr => \N__46890\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39940\,
            in1 => \N__38233\,
            in2 => \_gnd_net_\,
            in3 => \N__38214\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__47329\,
            ce => \N__38732\,
            sr => \N__46890\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39936\,
            in1 => \N__38209\,
            in2 => \_gnd_net_\,
            in3 => \N__38190\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__47329\,
            ce => \N__38732\,
            sr => \N__46890\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39941\,
            in1 => \N__38185\,
            in2 => \_gnd_net_\,
            in3 => \N__38166\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__47329\,
            ce => \N__38732\,
            sr => \N__46890\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39937\,
            in1 => \N__38161\,
            in2 => \_gnd_net_\,
            in3 => \N__38142\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__47329\,
            ce => \N__38732\,
            sr => \N__46890\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39942\,
            in1 => \N__38137\,
            in2 => \_gnd_net_\,
            in3 => \N__38118\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__47329\,
            ce => \N__38732\,
            sr => \N__46890\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39938\,
            in1 => \N__38503\,
            in2 => \_gnd_net_\,
            in3 => \N__38484\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__47329\,
            ce => \N__38732\,
            sr => \N__46890\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39930\,
            in1 => \N__38479\,
            in2 => \_gnd_net_\,
            in3 => \N__38460\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__47325\,
            ce => \N__38724\,
            sr => \N__46904\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39889\,
            in1 => \N__38455\,
            in2 => \_gnd_net_\,
            in3 => \N__38436\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__47325\,
            ce => \N__38724\,
            sr => \N__46904\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39927\,
            in1 => \N__38431\,
            in2 => \_gnd_net_\,
            in3 => \N__38412\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__47325\,
            ce => \N__38724\,
            sr => \N__46904\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39886\,
            in1 => \N__38407\,
            in2 => \_gnd_net_\,
            in3 => \N__38388\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__47325\,
            ce => \N__38724\,
            sr => \N__46904\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39928\,
            in1 => \N__38383\,
            in2 => \_gnd_net_\,
            in3 => \N__38364\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__47325\,
            ce => \N__38724\,
            sr => \N__46904\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39887\,
            in1 => \N__38359\,
            in2 => \_gnd_net_\,
            in3 => \N__38340\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__47325\,
            ce => \N__38724\,
            sr => \N__46904\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39929\,
            in1 => \N__38335\,
            in2 => \_gnd_net_\,
            in3 => \N__38316\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__47325\,
            ce => \N__38724\,
            sr => \N__46904\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39888\,
            in1 => \N__38311\,
            in2 => \_gnd_net_\,
            in3 => \N__38292\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__47325\,
            ce => \N__38724\,
            sr => \N__46904\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39931\,
            in1 => \N__38695\,
            in2 => \_gnd_net_\,
            in3 => \N__38676\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__47321\,
            ce => \N__38739\,
            sr => \N__46911\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39923\,
            in1 => \N__38671\,
            in2 => \_gnd_net_\,
            in3 => \N__38652\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__47321\,
            ce => \N__38739\,
            sr => \N__46911\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39932\,
            in1 => \N__38647\,
            in2 => \_gnd_net_\,
            in3 => \N__38628\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__47321\,
            ce => \N__38739\,
            sr => \N__46911\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39924\,
            in1 => \N__38623\,
            in2 => \_gnd_net_\,
            in3 => \N__38604\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__47321\,
            ce => \N__38739\,
            sr => \N__46911\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39933\,
            in1 => \N__38599\,
            in2 => \_gnd_net_\,
            in3 => \N__38580\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__47321\,
            ce => \N__38739\,
            sr => \N__46911\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39925\,
            in1 => \N__38575\,
            in2 => \_gnd_net_\,
            in3 => \N__38556\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__47321\,
            ce => \N__38739\,
            sr => \N__46911\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39934\,
            in1 => \N__38551\,
            in2 => \_gnd_net_\,
            in3 => \N__38532\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__47321\,
            ce => \N__38739\,
            sr => \N__46911\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39926\,
            in1 => \N__38527\,
            in2 => \_gnd_net_\,
            in3 => \N__38508\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__47321\,
            ce => \N__38739\,
            sr => \N__46911\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39917\,
            in1 => \N__38869\,
            in2 => \_gnd_net_\,
            in3 => \N__38850\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__47318\,
            ce => \N__38731\,
            sr => \N__46917\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39921\,
            in1 => \N__38845\,
            in2 => \_gnd_net_\,
            in3 => \N__38826\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__47318\,
            ce => \N__38731\,
            sr => \N__46917\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39918\,
            in1 => \N__38821\,
            in2 => \_gnd_net_\,
            in3 => \N__38802\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__47318\,
            ce => \N__38731\,
            sr => \N__46917\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39922\,
            in1 => \N__38797\,
            in2 => \_gnd_net_\,
            in3 => \N__38778\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__47318\,
            ce => \N__38731\,
            sr => \N__46917\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39919\,
            in1 => \N__38774\,
            in2 => \_gnd_net_\,
            in3 => \N__38760\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__47318\,
            ce => \N__38731\,
            sr => \N__46917\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__38753\,
            in1 => \N__39920\,
            in2 => \_gnd_net_\,
            in3 => \N__38757\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47318\,
            ce => \N__38731\,
            sr => \N__46917\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000000"
        )
    port map (
            in0 => \N__38925\,
            in1 => \N__38907\,
            in2 => \N__39099\,
            in3 => \N__39222\,
            lcout => \delay_measurement_inst.un1_elapsed_time_hc\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41335\,
            in1 => \N__41362\,
            in2 => \N__41285\,
            in3 => \N__41378\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64AN1_6_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__41182\,
            in1 => \N__41145\,
            in2 => \N__41258\,
            in3 => \N__41212\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__41705\,
            in1 => \N__41336\,
            in2 => \N__41609\,
            in3 => \N__41363\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINH2S1_14_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__41464\,
            in1 => \_gnd_net_\,
            in2 => \N__38937\,
            in3 => \N__41491\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINEU73_14_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001011101"
        )
    port map (
            in0 => \N__41492\,
            in1 => \N__39078\,
            in2 => \N__38934\,
            in3 => \N__41465\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_11_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41181\,
            in1 => \N__41579\,
            in2 => \N__41549\,
            in3 => \N__41213\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_11_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38898\,
            in1 => \N__39066\,
            in2 => \N__38916\,
            in3 => \N__38913\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclt31_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41250\,
            in1 => \N__41518\,
            in2 => \N__41150\,
            in3 => \N__41429\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41211\,
            in1 => \N__41180\,
            in2 => \N__41257\,
            in3 => \N__41463\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010011111100"
        )
    port map (
            in0 => \N__39060\,
            in1 => \N__41462\,
            in2 => \N__41149\,
            in3 => \N__38892\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100000000"
        )
    port map (
            in0 => \N__38883\,
            in1 => \N__39077\,
            in2 => \N__38874\,
            in3 => \N__39084\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41725\,
            in1 => \N__41404\,
            in2 => \N__41704\,
            in3 => \N__41428\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__41461\,
            in1 => \_gnd_net_\,
            in2 => \N__39087\,
            in3 => \N__41490\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41542\,
            in1 => \N__41572\,
            in2 => \N__41522\,
            in3 => \N__41602\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_17_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41405\,
            in1 => \N__41281\,
            in2 => \N__41312\,
            in3 => \N__41726\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41210\,
            in1 => \N__41305\,
            in2 => \N__41186\,
            in3 => \N__41460\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI339G_25_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41957\,
            in2 => \_gnd_net_\,
            in3 => \N__41630\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_27_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__41934\,
            in1 => \N__41943\,
            in2 => \N__39054\,
            in3 => \N__38943\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\,
            ltout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7L2RA_20_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__41675\,
            in1 => \N__39051\,
            in2 => \N__39045\,
            in3 => \N__46097\,
            lcout => \delay_measurement_inst.delay_hc_reg3lt31_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41925\,
            in1 => \N__41646\,
            in2 => \N__41916\,
            in3 => \N__41655\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02O13_20_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__46098\,
            in1 => \N__41676\,
            in2 => \N__41798\,
            in3 => \N__39228\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39213\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39192\,
            in2 => \N__39204\,
            in3 => \N__44152\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44135\,
            in1 => \N__39174\,
            in2 => \N__39186\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39156\,
            in2 => \N__39168\,
            in3 => \N__44099\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39141\,
            in2 => \N__39150\,
            in3 => \N__44063\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44042\,
            in1 => \N__39123\,
            in2 => \N__39135\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39105\,
            in2 => \N__39117\,
            in3 => \N__44018\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44573\,
            in1 => \N__39363\,
            in2 => \N__39372\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39348\,
            in2 => \N__39357\,
            in3 => \N__44546\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_16_12_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39330\,
            in2 => \N__39342\,
            in3 => \N__44525\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44504\,
            in1 => \N__39312\,
            in2 => \N__39324\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39288\,
            in2 => \N__39306\,
            in3 => \N__44480\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39267\,
            in2 => \N__39282\,
            in3 => \N__44453\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39261\,
            in2 => \N__39255\,
            in3 => \N__44423\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39234\,
            in2 => \N__39246\,
            in3 => \N__44390\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39471\,
            in2 => \N__39480\,
            in3 => \N__45005\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39453\,
            in2 => \N__39465\,
            in3 => \N__44981\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_16_13_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39432\,
            in2 => \N__39447\,
            in3 => \N__44960\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39411\,
            in2 => \N__39426\,
            in3 => \N__44936\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39390\,
            in2 => \N__39405\,
            in3 => \N__44915\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39384\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44647\,
            in2 => \N__39381\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__44648\,
            in1 => \N__44607\,
            in2 => \_gnd_net_\,
            in3 => \N__44156\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_7_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__45406\,
            in1 => \N__45574\,
            in2 => \N__45748\,
            in3 => \N__39558\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47375\,
            ce => 'H',
            sr => \N__46843\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_8_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__45575\,
            in1 => \N__45716\,
            in2 => \N__45441\,
            in3 => \N__39552\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47375\,
            ce => 'H',
            sr => \N__46843\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_9_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__45407\,
            in1 => \N__45576\,
            in2 => \N__45749\,
            in3 => \N__39546\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47375\,
            ce => 'H',
            sr => \N__46843\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39529\,
            in2 => \_gnd_net_\,
            in3 => \N__41072\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__45573\,
            in1 => \N__45715\,
            in2 => \_gnd_net_\,
            in3 => \N__45405\,
            lcout => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39530\,
            in2 => \_gnd_net_\,
            in3 => \N__41073\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_12_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__45446\,
            in1 => \N__45583\,
            in2 => \N__45750\,
            in3 => \N__39498\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47367\,
            ce => 'H',
            sr => \N__46846\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_18_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45726\,
            in1 => \N__45449\,
            in2 => \N__45598\,
            in3 => \N__39492\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47367\,
            ce => 'H',
            sr => \N__46846\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_10_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45724\,
            in1 => \N__45447\,
            in2 => \N__45596\,
            in3 => \N__39486\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47367\,
            ce => 'H',
            sr => \N__46846\
        );

    \delay_measurement_inst.delay_tr_reg_15_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__39699\,
            in1 => \N__39675\,
            in2 => \N__43253\,
            in3 => \N__39618\,
            lcout => measured_delay_tr_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47367\,
            ce => 'H',
            sr => \N__46846\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_11_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45725\,
            in1 => \N__45448\,
            in2 => \N__45597\,
            in3 => \N__39591\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47367\,
            ce => 'H',
            sr => \N__46846\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__47742\,
            in1 => \N__47605\,
            in2 => \N__47899\,
            in3 => \N__45108\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47367\,
            ce => 'H',
            sr => \N__46846\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001000000000"
        )
    port map (
            in0 => \N__40113\,
            in1 => \N__46155\,
            in2 => \N__40020\,
            in3 => \N__40053\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47359\,
            ce => \N__43067\,
            sr => \N__46854\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000101"
        )
    port map (
            in0 => \N__42823\,
            in1 => \N__42857\,
            in2 => \N__42783\,
            in3 => \N__43331\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47359\,
            ce => \N__43067\,
            sr => \N__46854\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__42781\,
            in1 => \N__46308\,
            in2 => \N__43343\,
            in3 => \N__42821\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47359\,
            ce => \N__43067\,
            sr => \N__46854\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__42777\,
            in1 => \N__42507\,
            in2 => \_gnd_net_\,
            in3 => \N__43332\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47359\,
            ce => \N__43067\,
            sr => \N__46854\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42776\,
            in2 => \N__43344\,
            in3 => \N__39585\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47359\,
            ce => \N__43067\,
            sr => \N__46854\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__42822\,
            in1 => \N__43330\,
            in2 => \N__46344\,
            in3 => \N__42782\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47359\,
            ce => \N__43067\,
            sr => \N__46854\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__43329\,
            in1 => \N__42894\,
            in2 => \_gnd_net_\,
            in3 => \N__43235\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47359\,
            ce => \N__43067\,
            sr => \N__46854\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011110011"
        )
    port map (
            in0 => \N__43234\,
            in1 => \N__43148\,
            in2 => \N__46260\,
            in3 => \N__46194\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47359\,
            ce => \N__43067\,
            sr => \N__46854\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40014\,
            in2 => \_gnd_net_\,
            in3 => \N__40112\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__46147\,
            in1 => \N__40077\,
            in2 => \N__40056\,
            in3 => \N__40048\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47353\,
            ce => \N__43062\,
            sr => \N__46864\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__40049\,
            in1 => \N__40015\,
            in2 => \_gnd_net_\,
            in3 => \N__46146\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47353\,
            ce => \N__43062\,
            sr => \N__46864\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39977\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39777\,
            in2 => \N__39810\,
            in3 => \N__39793\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_16_18_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39744\,
            in2 => \N__39771\,
            in3 => \N__39761\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39734\,
            in1 => \N__39705\,
            in2 => \N__39717\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40295\,
            in1 => \N__40278\,
            in2 => \N__42519\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40263\,
            in2 => \N__40272\,
            in3 => \N__45314\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40253\,
            in1 => \N__40239\,
            in2 => \N__42711\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40233\,
            in1 => \N__40218\,
            in2 => \N__42477\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40182\,
            in2 => \N__40212\,
            in3 => \N__40200\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40161\,
            in2 => \N__43398\,
            in3 => \N__40176\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40140\,
            in2 => \N__42693\,
            in3 => \N__40155\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40119\,
            in2 => \N__42657\,
            in3 => \N__40134\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40470\,
            in2 => \N__42624\,
            in3 => \N__40485\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40446\,
            in2 => \N__42579\,
            in3 => \N__40463\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40413\,
            in2 => \N__40440\,
            in3 => \N__40427\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40377\,
            in2 => \N__40407\,
            in3 => \N__40391\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40371\,
            in1 => \N__42864\,
            in2 => \N__40353\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40326\,
            in2 => \N__41040\,
            in3 => \N__40344\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_16_20_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40302\,
            in2 => \N__41031\,
            in3 => \N__40320\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41100\,
            in2 => \N__41022\,
            in3 => \N__41118\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41094\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_17_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46472\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47330\,
            ce => \N__43386\,
            sr => \N__46891\
        );

    \phase_controller_slave.stoper_tr.target_time_18_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46510\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47330\,
            ce => \N__43386\,
            sr => \N__46891\
        );

    \phase_controller_slave.stoper_tr.target_time_19_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46422\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47330\,
            ce => \N__43386\,
            sr => \N__46891\
        );

    \SB_DFF_inst_DELAY_HC1_LC_17_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41013\,
            lcout => delay_hc_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_17_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__40988\,
            in1 => \N__40959\,
            in2 => \_gnd_net_\,
            in3 => \N__43005\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_336_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_2_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__40877\,
            in1 => \N__40741\,
            in2 => \N__41367\,
            in3 => \N__40920\,
            lcout => measured_delay_hc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47444\,
            ce => 'H',
            sr => \N__46802\
        );

    \delay_measurement_inst.delay_hc_reg_15_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__40740\,
            in1 => \N__41469\,
            in2 => \N__40540\,
            in3 => \N__40644\,
            lcout => measured_delay_hc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47444\,
            ce => 'H',
            sr => \N__46802\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42969\,
            lcout => \delay_measurement_inst.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47437\,
            ce => \N__41747\,
            sr => \N__46805\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42948\,
            lcout => \delay_measurement_inst.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47437\,
            ce => \N__41747\,
            sr => \N__46805\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42968\,
            in2 => \N__42927\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_17_8_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__47429\,
            ce => \N__41748\,
            sr => \N__46808\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42947\,
            in2 => \N__43614\,
            in3 => \N__41292\,
            lcout => \delay_measurement_inst.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__47429\,
            ce => \N__41748\,
            sr => \N__46808\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42926\,
            in2 => \N__43590\,
            in3 => \N__41262\,
            lcout => \delay_measurement_inst.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__47429\,
            ce => \N__41748\,
            sr => \N__46808\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43613\,
            in2 => \N__43566\,
            in3 => \N__41223\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__47429\,
            ce => \N__41748\,
            sr => \N__46808\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43589\,
            in2 => \N__43542\,
            in3 => \N__41190\,
            lcout => \delay_measurement_inst.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__47429\,
            ce => \N__41748\,
            sr => \N__46808\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43565\,
            in2 => \N__43518\,
            in3 => \N__41157\,
            lcout => \delay_measurement_inst.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__47429\,
            ce => \N__41748\,
            sr => \N__46808\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43541\,
            in2 => \N__43494\,
            in3 => \N__41616\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__47429\,
            ce => \N__41748\,
            sr => \N__46808\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43517\,
            in2 => \N__43470\,
            in3 => \N__41586\,
            lcout => \delay_measurement_inst.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__47429\,
            ce => \N__41748\,
            sr => \N__46808\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43493\,
            in2 => \N__43446\,
            in3 => \N__41556\,
            lcout => \delay_measurement_inst.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__47422\,
            ce => \N__41749\,
            sr => \N__46811\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43469\,
            in2 => \N__43422\,
            in3 => \N__41526\,
            lcout => \delay_measurement_inst.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__47422\,
            ce => \N__41749\,
            sr => \N__46811\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43445\,
            in2 => \N__43806\,
            in3 => \N__41499\,
            lcout => \delay_measurement_inst.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__47422\,
            ce => \N__41749\,
            sr => \N__46811\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43421\,
            in2 => \N__43782\,
            in3 => \N__41472\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__47422\,
            ce => \N__41749\,
            sr => \N__46811\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43805\,
            in2 => \N__43758\,
            in3 => \N__41436\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__47422\,
            ce => \N__41749\,
            sr => \N__46811\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43781\,
            in2 => \N__43734\,
            in3 => \N__41412\,
            lcout => \delay_measurement_inst.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__47422\,
            ce => \N__41749\,
            sr => \N__46811\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43757\,
            in2 => \N__43710\,
            in3 => \N__41391\,
            lcout => \delay_measurement_inst.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__47422\,
            ce => \N__41749\,
            sr => \N__46811\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43733\,
            in2 => \N__43686\,
            in3 => \N__41712\,
            lcout => \delay_measurement_inst.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__47422\,
            ce => \N__41749\,
            sr => \N__46811\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43709\,
            in2 => \N__43662\,
            in3 => \N__41679\,
            lcout => \delay_measurement_inst.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__47415\,
            ce => \N__41750\,
            sr => \N__46815\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43685\,
            in2 => \N__43638\,
            in3 => \N__41664\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__47415\,
            ce => \N__41750\,
            sr => \N__46815\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43661\,
            in2 => \N__43998\,
            in3 => \N__41661\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__47415\,
            ce => \N__41750\,
            sr => \N__46815\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43637\,
            in2 => \N__43974\,
            in3 => \N__41658\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__47415\,
            ce => \N__41750\,
            sr => \N__46815\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43997\,
            in2 => \N__43950\,
            in3 => \N__41649\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__47415\,
            ce => \N__41750\,
            sr => \N__46815\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43973\,
            in2 => \N__43926\,
            in3 => \N__41640\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__47415\,
            ce => \N__41750\,
            sr => \N__46815\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43949\,
            in2 => \N__43902\,
            in3 => \N__41619\,
            lcout => \delay_measurement_inst.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__47415\,
            ce => \N__41750\,
            sr => \N__46815\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43925\,
            in2 => \N__43878\,
            in3 => \N__41946\,
            lcout => \delay_measurement_inst.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__47415\,
            ce => \N__41750\,
            sr => \N__46815\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43901\,
            in2 => \N__43854\,
            in3 => \N__41937\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__47407\,
            ce => \N__41751\,
            sr => \N__46820\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43877\,
            in2 => \N__43830\,
            in3 => \N__41928\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__47407\,
            ce => \N__41751\,
            sr => \N__46820\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43853\,
            in2 => \N__44367\,
            in3 => \N__41919\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__47407\,
            ce => \N__41751\,
            sr => \N__46820\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43829\,
            in2 => \N__44226\,
            in3 => \N__41907\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__47407\,
            ce => \N__41751\,
            sr => \N__46820\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41904\,
            lcout => \delay_measurement_inst.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47407\,
            ce => \N__41751\,
            sr => \N__46820\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_4_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__44752\,
            in1 => \N__44887\,
            in2 => \N__42222\,
            in3 => \N__44052\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47398\,
            ce => 'H',
            sr => \N__46825\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_5_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__44885\,
            in1 => \N__42207\,
            in2 => \N__44031\,
            in3 => \N__44758\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47398\,
            ce => 'H',
            sr => \N__46825\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_6_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__44753\,
            in1 => \N__44888\,
            in2 => \N__42223\,
            in3 => \N__44007\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47398\,
            ce => 'H',
            sr => \N__46825\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_7_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__44886\,
            in1 => \N__42208\,
            in2 => \N__44562\,
            in3 => \N__44759\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47398\,
            ce => 'H',
            sr => \N__46825\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_8_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__44754\,
            in1 => \N__44889\,
            in2 => \N__42224\,
            in3 => \N__44535\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47398\,
            ce => 'H',
            sr => \N__46825\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__44883\,
            in1 => \N__42205\,
            in2 => \N__44442\,
            in3 => \N__44756\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47398\,
            ce => 'H',
            sr => \N__46825\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_9_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__44755\,
            in1 => \N__44890\,
            in2 => \N__42225\,
            in3 => \N__44514\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47398\,
            ce => 'H',
            sr => \N__46825\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__44884\,
            in1 => \N__42206\,
            in2 => \N__44994\,
            in3 => \N__44757\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47398\,
            ce => 'H',
            sr => \N__46825\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_10_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__44875\,
            in1 => \N__44493\,
            in2 => \N__42218\,
            in3 => \N__44771\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47388\,
            ce => 'H',
            sr => \N__46830\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_14_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__44764\,
            in1 => \N__42176\,
            in2 => \N__44379\,
            in3 => \N__44879\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47388\,
            ce => 'H',
            sr => \N__46830\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__44876\,
            in1 => \N__44768\,
            in2 => \N__42219\,
            in3 => \N__44970\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47388\,
            ce => 'H',
            sr => \N__46830\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__44765\,
            in1 => \N__42177\,
            in2 => \N__44949\,
            in3 => \N__44880\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47388\,
            ce => 'H',
            sr => \N__46830\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__44877\,
            in1 => \N__44769\,
            in2 => \N__42220\,
            in3 => \N__44925\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47388\,
            ce => 'H',
            sr => \N__46830\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_19_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__44766\,
            in1 => \N__42178\,
            in2 => \N__44901\,
            in3 => \N__44881\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47388\,
            ce => 'H',
            sr => \N__46830\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_2_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__44878\,
            in1 => \N__44770\,
            in2 => \N__42221\,
            in3 => \N__44118\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47388\,
            ce => 'H',
            sr => \N__46830\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_3_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__44767\,
            in1 => \N__42179\,
            in2 => \N__44082\,
            in3 => \N__44882\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47388\,
            ce => 'H',
            sr => \N__46830\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__47572\,
            in1 => \N__47892\,
            in2 => \N__47743\,
            in3 => \N__45174\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47380\,
            ce => 'H',
            sr => \N__46835\
        );

    \phase_controller_inst1.start_timer_tr_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__42084\,
            in1 => \N__42071\,
            in2 => \N__47931\,
            in3 => \N__42033\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47380\,
            ce => 'H',
            sr => \N__46835\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__47571\,
            in1 => \N__47729\,
            in2 => \_gnd_net_\,
            in3 => \N__47891\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110111000000"
        )
    port map (
            in0 => \N__45959\,
            in1 => \N__41997\,
            in2 => \N__42012\,
            in3 => \N__45994\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47380\,
            ce => 'H',
            sr => \N__46835\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45987\,
            in2 => \_gnd_net_\,
            in3 => \N__45958\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__47730\,
            in1 => \N__45144\,
            in2 => \N__47930\,
            in3 => \N__47573\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47380\,
            ce => 'H',
            sr => \N__46835\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45923\,
            in1 => \N__41967\,
            in2 => \N__41979\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42345\,
            in2 => \N__42357\,
            in3 => \N__45119\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42324\,
            in2 => \N__42339\,
            in3 => \N__45278\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42309\,
            in2 => \N__42318\,
            in3 => \N__45248\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45221\,
            in1 => \N__42291\,
            in2 => \N__42303\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42276\,
            in2 => \N__42285\,
            in3 => \N__46070\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46043\,
            in1 => \N__42258\,
            in2 => \N__42270\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42252\,
            in2 => \N__42240\,
            in3 => \N__45077\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42456\,
            in2 => \N__42465\,
            in3 => \N__45044\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46013\,
            in1 => \N__42450\,
            in2 => \N__43083\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42432\,
            in2 => \N__42444\,
            in3 => \N__45890\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42414\,
            in2 => \N__42426\,
            in3 => \N__45863\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45833\,
            in1 => \N__42393\,
            in2 => \N__42408\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42375\,
            in2 => \N__42387\,
            in3 => \N__47957\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__47480\,
            in1 => \N__42369\,
            in2 => \N__43188\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45189\,
            in1 => \N__42363\,
            in2 => \N__43173\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42567\,
            in2 => \N__42546\,
            in3 => \N__45161\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42561\,
            in2 => \N__42537\,
            in3 => \N__45794\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42555\,
            in2 => \N__42528\,
            in3 => \N__45776\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42549\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46473\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47360\,
            ce => \N__43063\,
            sr => \N__46855\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46515\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47360\,
            ce => \N__43063\,
            sr => \N__46855\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46433\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47360\,
            ce => \N__43063\,
            sr => \N__46855\
        );

    \phase_controller_slave.stoper_tr.target_time_4_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__42773\,
            in1 => \N__43301\,
            in2 => \N__46307\,
            in3 => \N__42824\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47354\,
            ce => \N__43384\,
            sr => \N__46865\
        );

    \phase_controller_slave.stoper_tr.target_time_7_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__43300\,
            in1 => \N__42506\,
            in2 => \_gnd_net_\,
            in3 => \N__42774\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47354\,
            ce => \N__43384\,
            sr => \N__46865\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43239\,
            in2 => \_gnd_net_\,
            in3 => \N__42903\,
            lcout => \phase_controller_inst1.stoper_tr.N_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_16_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46383\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47354\,
            ce => \N__43384\,
            sr => \N__46865\
        );

    \phase_controller_slave.stoper_tr.target_time_6_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110000001101"
        )
    port map (
            in0 => \N__43299\,
            in1 => \N__42858\,
            in2 => \N__42828\,
            in3 => \N__42775\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47344\,
            ce => \N__43385\,
            sr => \N__46875\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__46471\,
            in1 => \N__46381\,
            in2 => \N__46432\,
            in3 => \N__46506\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42699\,
            in3 => \N__46272\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_10_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42696\,
            in3 => \N__43109\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47344\,
            ce => \N__43385\,
            sr => \N__46875\
        );

    \phase_controller_slave.stoper_tr.target_time_11_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43137\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42681\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47344\,
            ce => \N__43385\,
            sr => \N__46875\
        );

    \phase_controller_slave.stoper_tr.target_time_12_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43138\,
            in2 => \_gnd_net_\,
            in3 => \N__42648\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47344\,
            ce => \N__43385\,
            sr => \N__46875\
        );

    \phase_controller_slave.stoper_tr.target_time_13_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43139\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42607\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47344\,
            ce => \N__43385\,
            sr => \N__46875\
        );

    \phase_controller_slave.stoper_tr.target_time_9_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010111011"
        )
    port map (
            in0 => \N__46256\,
            in1 => \N__43140\,
            in2 => \N__43260\,
            in3 => \N__46193\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47344\,
            ce => \N__43385\,
            sr => \N__46875\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43302\,
            in2 => \_gnd_net_\,
            in3 => \N__43257\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47336\,
            ce => \N__43068\,
            sr => \N__46884\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46382\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47336\,
            ce => \N__43068\,
            sr => \N__46884\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43141\,
            in2 => \_gnd_net_\,
            in3 => \N__43110\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47336\,
            ce => \N__43068\,
            sr => \N__46884\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_18_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43001\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44320\,
            in1 => \N__42967\,
            in2 => \_gnd_net_\,
            in3 => \N__42951\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_7_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__47445\,
            ce => \N__44205\,
            sr => \N__46803\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44342\,
            in1 => \N__42946\,
            in2 => \_gnd_net_\,
            in3 => \N__42930\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__47445\,
            ce => \N__44205\,
            sr => \N__46803\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44321\,
            in1 => \N__42925\,
            in2 => \_gnd_net_\,
            in3 => \N__42906\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__47445\,
            ce => \N__44205\,
            sr => \N__46803\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44343\,
            in1 => \N__43612\,
            in2 => \_gnd_net_\,
            in3 => \N__43593\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__47445\,
            ce => \N__44205\,
            sr => \N__46803\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44322\,
            in1 => \N__43588\,
            in2 => \_gnd_net_\,
            in3 => \N__43569\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__47445\,
            ce => \N__44205\,
            sr => \N__46803\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44344\,
            in1 => \N__43564\,
            in2 => \_gnd_net_\,
            in3 => \N__43545\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__47445\,
            ce => \N__44205\,
            sr => \N__46803\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44323\,
            in1 => \N__43540\,
            in2 => \_gnd_net_\,
            in3 => \N__43521\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__47445\,
            ce => \N__44205\,
            sr => \N__46803\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44345\,
            in1 => \N__43516\,
            in2 => \_gnd_net_\,
            in3 => \N__43497\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__47445\,
            ce => \N__44205\,
            sr => \N__46803\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44333\,
            in1 => \N__43492\,
            in2 => \_gnd_net_\,
            in3 => \N__43473\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_18_8_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__47438\,
            ce => \N__44207\,
            sr => \N__46806\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44349\,
            in1 => \N__43468\,
            in2 => \_gnd_net_\,
            in3 => \N__43449\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__47438\,
            ce => \N__44207\,
            sr => \N__46806\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44330\,
            in1 => \N__43444\,
            in2 => \_gnd_net_\,
            in3 => \N__43425\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__47438\,
            ce => \N__44207\,
            sr => \N__46806\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44346\,
            in1 => \N__43420\,
            in2 => \_gnd_net_\,
            in3 => \N__43401\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__47438\,
            ce => \N__44207\,
            sr => \N__46806\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44331\,
            in1 => \N__43804\,
            in2 => \_gnd_net_\,
            in3 => \N__43785\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__47438\,
            ce => \N__44207\,
            sr => \N__46806\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44347\,
            in1 => \N__43780\,
            in2 => \_gnd_net_\,
            in3 => \N__43761\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__47438\,
            ce => \N__44207\,
            sr => \N__46806\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44332\,
            in1 => \N__43756\,
            in2 => \_gnd_net_\,
            in3 => \N__43737\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__47438\,
            ce => \N__44207\,
            sr => \N__46806\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44348\,
            in1 => \N__43732\,
            in2 => \_gnd_net_\,
            in3 => \N__43713\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__47438\,
            ce => \N__44207\,
            sr => \N__46806\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44334\,
            in1 => \N__43708\,
            in2 => \_gnd_net_\,
            in3 => \N__43689\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_18_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__47430\,
            ce => \N__44206\,
            sr => \N__46809\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44338\,
            in1 => \N__43684\,
            in2 => \_gnd_net_\,
            in3 => \N__43665\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__47430\,
            ce => \N__44206\,
            sr => \N__46809\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44335\,
            in1 => \N__43660\,
            in2 => \_gnd_net_\,
            in3 => \N__43641\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__47430\,
            ce => \N__44206\,
            sr => \N__46809\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44339\,
            in1 => \N__43636\,
            in2 => \_gnd_net_\,
            in3 => \N__43617\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__47430\,
            ce => \N__44206\,
            sr => \N__46809\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44336\,
            in1 => \N__43996\,
            in2 => \_gnd_net_\,
            in3 => \N__43977\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__47430\,
            ce => \N__44206\,
            sr => \N__46809\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44340\,
            in1 => \N__43972\,
            in2 => \_gnd_net_\,
            in3 => \N__43953\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__47430\,
            ce => \N__44206\,
            sr => \N__46809\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44337\,
            in1 => \N__43948\,
            in2 => \_gnd_net_\,
            in3 => \N__43929\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__47430\,
            ce => \N__44206\,
            sr => \N__46809\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44341\,
            in1 => \N__43924\,
            in2 => \_gnd_net_\,
            in3 => \N__43905\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__47430\,
            ce => \N__44206\,
            sr => \N__46809\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44324\,
            in1 => \N__43900\,
            in2 => \_gnd_net_\,
            in3 => \N__43881\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_18_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__47423\,
            ce => \N__44211\,
            sr => \N__46812\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44328\,
            in1 => \N__43876\,
            in2 => \_gnd_net_\,
            in3 => \N__43857\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__47423\,
            ce => \N__44211\,
            sr => \N__46812\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44325\,
            in1 => \N__43852\,
            in2 => \_gnd_net_\,
            in3 => \N__43833\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__47423\,
            ce => \N__44211\,
            sr => \N__46812\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44329\,
            in1 => \N__43828\,
            in2 => \_gnd_net_\,
            in3 => \N__43809\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__47423\,
            ce => \N__44211\,
            sr => \N__46812\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44326\,
            in1 => \N__44366\,
            in2 => \_gnd_net_\,
            in3 => \N__44352\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__47423\,
            ce => \N__44211\,
            sr => \N__46812\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__44225\,
            in1 => \N__44327\,
            in2 => \_gnd_net_\,
            in3 => \N__44229\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47423\,
            ce => \N__44211\,
            sr => \N__46812\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44175\,
            in2 => \N__44163\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_11_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44136\,
            in2 => \_gnd_net_\,
            in3 => \N__44106\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44583\,
            in2 => \N__44103\,
            in3 => \N__44067\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44064\,
            in2 => \_gnd_net_\,
            in3 => \N__44046\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44043\,
            in2 => \_gnd_net_\,
            in3 => \N__44022\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44019\,
            in2 => \_gnd_net_\,
            in3 => \N__44001\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44574\,
            in2 => \_gnd_net_\,
            in3 => \N__44550\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44547\,
            in2 => \_gnd_net_\,
            in3 => \N__44529\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44526\,
            in2 => \_gnd_net_\,
            in3 => \N__44508\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44505\,
            in2 => \_gnd_net_\,
            in3 => \N__44487\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44484\,
            in2 => \_gnd_net_\,
            in3 => \N__44457\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44454\,
            in2 => \_gnd_net_\,
            in3 => \N__44430\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44427\,
            in2 => \_gnd_net_\,
            in3 => \N__44394\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44391\,
            in2 => \_gnd_net_\,
            in3 => \N__44370\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45006\,
            in2 => \_gnd_net_\,
            in3 => \N__44985\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44982\,
            in2 => \_gnd_net_\,
            in3 => \N__44964\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44961\,
            in2 => \_gnd_net_\,
            in3 => \N__44940\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44937\,
            in2 => \_gnd_net_\,
            in3 => \N__44919\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44916\,
            in2 => \_gnd_net_\,
            in3 => \N__44904\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47734\,
            in2 => \_gnd_net_\,
            in3 => \N__47536\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44874\,
            in2 => \_gnd_net_\,
            in3 => \N__44763\,
            lcout => \phase_controller_slave.stoper_hc.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44643\,
            in2 => \_gnd_net_\,
            in3 => \N__44611\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45132\,
            in2 => \N__45927\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45126\,
            in2 => \_gnd_net_\,
            in3 => \N__45096\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45813\,
            in2 => \N__45282\,
            in3 => \N__45093\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45249\,
            in2 => \_gnd_net_\,
            in3 => \N__45090\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45222\,
            in2 => \_gnd_net_\,
            in3 => \N__45087\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46074\,
            in2 => \_gnd_net_\,
            in3 => \N__45084\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46044\,
            in2 => \_gnd_net_\,
            in3 => \N__45081\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45078\,
            in2 => \_gnd_net_\,
            in3 => \N__45048\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45045\,
            in2 => \_gnd_net_\,
            in3 => \N__45009\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46014\,
            in2 => \_gnd_net_\,
            in3 => \N__45207\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45891\,
            in2 => \_gnd_net_\,
            in3 => \N__45204\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45864\,
            in2 => \_gnd_net_\,
            in3 => \N__45201\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45834\,
            in2 => \_gnd_net_\,
            in3 => \N__45198\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47958\,
            in2 => \_gnd_net_\,
            in3 => \N__45195\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47481\,
            in2 => \_gnd_net_\,
            in3 => \N__45192\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45188\,
            in2 => \_gnd_net_\,
            in3 => \N__45168\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45165\,
            in2 => \_gnd_net_\,
            in3 => \N__45135\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45795\,
            in2 => \_gnd_net_\,
            in3 => \N__45819\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45777\,
            in2 => \_gnd_net_\,
            in3 => \N__45816\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45995\,
            in2 => \_gnd_net_\,
            in3 => \N__45956\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__47621\,
            in1 => \N__47789\,
            in2 => \N__45804\,
            in3 => \N__47921\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47368\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__47781\,
            in1 => \N__47624\,
            in2 => \N__47936\,
            in3 => \N__45783\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47368\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_5_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010000010"
        )
    port map (
            in0 => \N__45765\,
            in1 => \N__45731\,
            in2 => \N__45600\,
            in3 => \N__45450\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47368\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010001010"
        )
    port map (
            in0 => \N__45291\,
            in1 => \N__47627\,
            in2 => \N__47790\,
            in3 => \N__47924\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47368\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__47622\,
            in1 => \N__47922\,
            in2 => \N__45261\,
            in3 => \N__47784\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47368\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__47782\,
            in1 => \N__47625\,
            in2 => \N__47937\,
            in3 => \N__45231\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47368\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__47623\,
            in1 => \N__47923\,
            in2 => \N__46086\,
            in3 => \N__47785\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47368\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__47783\,
            in1 => \N__47626\,
            in2 => \N__47938\,
            in3 => \N__46056\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47368\,
            ce => 'H',
            sr => \N__46847\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__47774\,
            in1 => \N__47909\,
            in2 => \N__47628\,
            in3 => \N__46026\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47361\,
            ce => 'H',
            sr => \N__46856\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__45999\,
            in1 => \N__45922\,
            in2 => \_gnd_net_\,
            in3 => \N__45957\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__47777\,
            in1 => \N__47908\,
            in2 => \N__45930\,
            in3 => \N__47620\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47361\,
            ce => 'H',
            sr => \N__46856\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010100010"
        )
    port map (
            in0 => \N__45900\,
            in1 => \N__47778\,
            in2 => \N__47631\,
            in3 => \N__47925\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47361\,
            ce => 'H',
            sr => \N__46856\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__47775\,
            in1 => \N__47910\,
            in2 => \N__47629\,
            in3 => \N__45873\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47361\,
            ce => 'H',
            sr => \N__46856\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__47906\,
            in1 => \N__47779\,
            in2 => \N__45846\,
            in3 => \N__47615\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47361\,
            ce => 'H',
            sr => \N__46856\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__47776\,
            in1 => \N__47911\,
            in2 => \N__47630\,
            in3 => \N__47967\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47361\,
            ce => 'H',
            sr => \N__46856\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__47907\,
            in1 => \N__47780\,
            in2 => \N__47646\,
            in3 => \N__47616\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47361\,
            ce => 'H',
            sr => \N__46856\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__46514\,
            in1 => \N__46470\,
            in2 => \N__46434\,
            in3 => \N__46380\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__46340\,
            in1 => \N__46306\,
            in2 => \N__46275\,
            in3 => \N__46271\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__46248\,
            in1 => \N__46215\,
            in2 => \N__46197\,
            in3 => \N__46192\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46116\,
            in2 => \_gnd_net_\,
            in3 => \N__46107\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
