// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Oct 8 2025 23:57:57

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    start_stop,
    s2_phy,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    input start_stop;
    output s2_phy;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__22544;
    wire N__22543;
    wire N__22542;
    wire N__22533;
    wire N__22532;
    wire N__22531;
    wire N__22524;
    wire N__22523;
    wire N__22522;
    wire N__22515;
    wire N__22514;
    wire N__22513;
    wire N__22506;
    wire N__22505;
    wire N__22504;
    wire N__22497;
    wire N__22496;
    wire N__22495;
    wire N__22488;
    wire N__22487;
    wire N__22486;
    wire N__22479;
    wire N__22478;
    wire N__22477;
    wire N__22470;
    wire N__22469;
    wire N__22468;
    wire N__22461;
    wire N__22460;
    wire N__22459;
    wire N__22452;
    wire N__22451;
    wire N__22450;
    wire N__22443;
    wire N__22442;
    wire N__22441;
    wire N__22434;
    wire N__22433;
    wire N__22432;
    wire N__22415;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22378;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22361;
    wire N__22360;
    wire N__22359;
    wire N__22356;
    wire N__22353;
    wire N__22350;
    wire N__22343;
    wire N__22342;
    wire N__22341;
    wire N__22340;
    wire N__22339;
    wire N__22336;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22304;
    wire N__22303;
    wire N__22302;
    wire N__22301;
    wire N__22300;
    wire N__22299;
    wire N__22298;
    wire N__22297;
    wire N__22296;
    wire N__22295;
    wire N__22294;
    wire N__22293;
    wire N__22292;
    wire N__22291;
    wire N__22290;
    wire N__22289;
    wire N__22288;
    wire N__22287;
    wire N__22286;
    wire N__22285;
    wire N__22284;
    wire N__22283;
    wire N__22282;
    wire N__22281;
    wire N__22280;
    wire N__22279;
    wire N__22278;
    wire N__22277;
    wire N__22276;
    wire N__22275;
    wire N__22274;
    wire N__22273;
    wire N__22272;
    wire N__22271;
    wire N__22270;
    wire N__22269;
    wire N__22266;
    wire N__22265;
    wire N__22264;
    wire N__22263;
    wire N__22262;
    wire N__22261;
    wire N__22260;
    wire N__22259;
    wire N__22258;
    wire N__22257;
    wire N__22256;
    wire N__22255;
    wire N__22254;
    wire N__22253;
    wire N__22252;
    wire N__22251;
    wire N__22250;
    wire N__22249;
    wire N__22248;
    wire N__22247;
    wire N__22244;
    wire N__22243;
    wire N__22242;
    wire N__22241;
    wire N__22240;
    wire N__22239;
    wire N__22238;
    wire N__22237;
    wire N__22236;
    wire N__22235;
    wire N__22234;
    wire N__22233;
    wire N__22232;
    wire N__22231;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22075;
    wire N__22072;
    wire N__22071;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22051;
    wire N__22048;
    wire N__22043;
    wire N__22042;
    wire N__22041;
    wire N__22040;
    wire N__22039;
    wire N__22038;
    wire N__22037;
    wire N__22036;
    wire N__22035;
    wire N__22034;
    wire N__22033;
    wire N__22032;
    wire N__22031;
    wire N__22030;
    wire N__22029;
    wire N__22028;
    wire N__22027;
    wire N__22026;
    wire N__22025;
    wire N__22024;
    wire N__22023;
    wire N__22022;
    wire N__22021;
    wire N__22020;
    wire N__22019;
    wire N__22018;
    wire N__22017;
    wire N__22016;
    wire N__22015;
    wire N__22014;
    wire N__22013;
    wire N__22012;
    wire N__22011;
    wire N__22010;
    wire N__22009;
    wire N__22008;
    wire N__22007;
    wire N__22006;
    wire N__22005;
    wire N__22004;
    wire N__22003;
    wire N__22002;
    wire N__22001;
    wire N__22000;
    wire N__21999;
    wire N__21998;
    wire N__21997;
    wire N__21996;
    wire N__21995;
    wire N__21994;
    wire N__21993;
    wire N__21992;
    wire N__21991;
    wire N__21990;
    wire N__21989;
    wire N__21988;
    wire N__21987;
    wire N__21986;
    wire N__21985;
    wire N__21984;
    wire N__21983;
    wire N__21982;
    wire N__21981;
    wire N__21980;
    wire N__21979;
    wire N__21978;
    wire N__21977;
    wire N__21976;
    wire N__21975;
    wire N__21974;
    wire N__21973;
    wire N__21972;
    wire N__21971;
    wire N__21970;
    wire N__21969;
    wire N__21968;
    wire N__21967;
    wire N__21966;
    wire N__21965;
    wire N__21964;
    wire N__21963;
    wire N__21962;
    wire N__21961;
    wire N__21960;
    wire N__21959;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21781;
    wire N__21778;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21761;
    wire N__21760;
    wire N__21759;
    wire N__21756;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21710;
    wire N__21709;
    wire N__21708;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21660;
    wire N__21657;
    wire N__21652;
    wire N__21649;
    wire N__21644;
    wire N__21643;
    wire N__21642;
    wire N__21639;
    wire N__21638;
    wire N__21637;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21607;
    wire N__21606;
    wire N__21603;
    wire N__21600;
    wire N__21597;
    wire N__21596;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21556;
    wire N__21553;
    wire N__21552;
    wire N__21549;
    wire N__21548;
    wire N__21545;
    wire N__21540;
    wire N__21537;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21514;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21497;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21485;
    wire N__21484;
    wire N__21481;
    wire N__21480;
    wire N__21479;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21467;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21425;
    wire N__21422;
    wire N__21421;
    wire N__21420;
    wire N__21419;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21405;
    wire N__21402;
    wire N__21395;
    wire N__21394;
    wire N__21393;
    wire N__21392;
    wire N__21389;
    wire N__21384;
    wire N__21381;
    wire N__21374;
    wire N__21373;
    wire N__21372;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21350;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21342;
    wire N__21339;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21324;
    wire N__21319;
    wire N__21316;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21306;
    wire N__21301;
    wire N__21298;
    wire N__21293;
    wire N__21290;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21278;
    wire N__21275;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21248;
    wire N__21247;
    wire N__21244;
    wire N__21241;
    wire N__21240;
    wire N__21235;
    wire N__21232;
    wire N__21227;
    wire N__21226;
    wire N__21223;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21206;
    wire N__21205;
    wire N__21204;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21182;
    wire N__21181;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21130;
    wire N__21127;
    wire N__21126;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21076;
    wire N__21075;
    wire N__21074;
    wire N__21073;
    wire N__21072;
    wire N__21067;
    wire N__21066;
    wire N__21065;
    wire N__21064;
    wire N__21063;
    wire N__21062;
    wire N__21061;
    wire N__21060;
    wire N__21059;
    wire N__21058;
    wire N__21057;
    wire N__21056;
    wire N__21055;
    wire N__21046;
    wire N__21045;
    wire N__21044;
    wire N__21043;
    wire N__21042;
    wire N__21041;
    wire N__21040;
    wire N__21039;
    wire N__21038;
    wire N__21037;
    wire N__21036;
    wire N__21035;
    wire N__21034;
    wire N__21031;
    wire N__21022;
    wire N__21013;
    wire N__21004;
    wire N__21001;
    wire N__20992;
    wire N__20983;
    wire N__20974;
    wire N__20969;
    wire N__20962;
    wire N__20951;
    wire N__20948;
    wire N__20947;
    wire N__20946;
    wire N__20945;
    wire N__20944;
    wire N__20943;
    wire N__20942;
    wire N__20941;
    wire N__20940;
    wire N__20939;
    wire N__20938;
    wire N__20937;
    wire N__20936;
    wire N__20935;
    wire N__20932;
    wire N__20921;
    wire N__20914;
    wire N__20907;
    wire N__20902;
    wire N__20899;
    wire N__20896;
    wire N__20889;
    wire N__20886;
    wire N__20881;
    wire N__20878;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20854;
    wire N__20849;
    wire N__20846;
    wire N__20845;
    wire N__20844;
    wire N__20843;
    wire N__20842;
    wire N__20841;
    wire N__20840;
    wire N__20839;
    wire N__20838;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20827;
    wire N__20826;
    wire N__20825;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20815;
    wire N__20814;
    wire N__20813;
    wire N__20812;
    wire N__20811;
    wire N__20810;
    wire N__20809;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20781;
    wire N__20780;
    wire N__20779;
    wire N__20778;
    wire N__20775;
    wire N__20766;
    wire N__20763;
    wire N__20746;
    wire N__20743;
    wire N__20738;
    wire N__20735;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20718;
    wire N__20715;
    wire N__20712;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20690;
    wire N__20689;
    wire N__20684;
    wire N__20681;
    wire N__20680;
    wire N__20679;
    wire N__20674;
    wire N__20671;
    wire N__20666;
    wire N__20663;
    wire N__20660;
    wire N__20657;
    wire N__20656;
    wire N__20655;
    wire N__20654;
    wire N__20653;
    wire N__20652;
    wire N__20651;
    wire N__20650;
    wire N__20649;
    wire N__20648;
    wire N__20647;
    wire N__20646;
    wire N__20645;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20634;
    wire N__20633;
    wire N__20632;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20617;
    wire N__20616;
    wire N__20615;
    wire N__20612;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20595;
    wire N__20594;
    wire N__20581;
    wire N__20572;
    wire N__20565;
    wire N__20560;
    wire N__20551;
    wire N__20546;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20534;
    wire N__20527;
    wire N__20524;
    wire N__20523;
    wire N__20520;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20498;
    wire N__20497;
    wire N__20496;
    wire N__20491;
    wire N__20488;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20472;
    wire N__20465;
    wire N__20464;
    wire N__20463;
    wire N__20458;
    wire N__20455;
    wire N__20450;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20438;
    wire N__20437;
    wire N__20436;
    wire N__20435;
    wire N__20432;
    wire N__20427;
    wire N__20424;
    wire N__20417;
    wire N__20416;
    wire N__20411;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20403;
    wire N__20400;
    wire N__20397;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20374;
    wire N__20369;
    wire N__20366;
    wire N__20365;
    wire N__20362;
    wire N__20359;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20344;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20300;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20288;
    wire N__20287;
    wire N__20286;
    wire N__20285;
    wire N__20282;
    wire N__20277;
    wire N__20274;
    wire N__20267;
    wire N__20266;
    wire N__20263;
    wire N__20262;
    wire N__20257;
    wire N__20254;
    wire N__20249;
    wire N__20248;
    wire N__20245;
    wire N__20242;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20209;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20191;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20137;
    wire N__20136;
    wire N__20135;
    wire N__20132;
    wire N__20131;
    wire N__20130;
    wire N__20129;
    wire N__20128;
    wire N__20121;
    wire N__20120;
    wire N__20119;
    wire N__20118;
    wire N__20117;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20109;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20089;
    wire N__20086;
    wire N__20083;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20071;
    wire N__20070;
    wire N__20067;
    wire N__20062;
    wire N__20059;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20033;
    wire N__20032;
    wire N__20031;
    wire N__20028;
    wire N__20027;
    wire N__20026;
    wire N__20021;
    wire N__20020;
    wire N__20019;
    wire N__20018;
    wire N__20015;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19997;
    wire N__19996;
    wire N__19993;
    wire N__19986;
    wire N__19983;
    wire N__19978;
    wire N__19975;
    wire N__19970;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19945;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19930;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19907;
    wire N__19906;
    wire N__19905;
    wire N__19904;
    wire N__19903;
    wire N__19902;
    wire N__19901;
    wire N__19900;
    wire N__19899;
    wire N__19898;
    wire N__19895;
    wire N__19894;
    wire N__19893;
    wire N__19892;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19878;
    wire N__19877;
    wire N__19874;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19860;
    wire N__19859;
    wire N__19858;
    wire N__19857;
    wire N__19854;
    wire N__19837;
    wire N__19830;
    wire N__19827;
    wire N__19810;
    wire N__19807;
    wire N__19802;
    wire N__19799;
    wire N__19794;
    wire N__19791;
    wire N__19790;
    wire N__19789;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19758;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19735;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19718;
    wire N__19715;
    wire N__19714;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19706;
    wire N__19705;
    wire N__19702;
    wire N__19697;
    wire N__19692;
    wire N__19685;
    wire N__19684;
    wire N__19683;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19669;
    wire N__19664;
    wire N__19661;
    wire N__19660;
    wire N__19659;
    wire N__19656;
    wire N__19653;
    wire N__19650;
    wire N__19645;
    wire N__19640;
    wire N__19637;
    wire N__19636;
    wire N__19635;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19616;
    wire N__19613;
    wire N__19612;
    wire N__19611;
    wire N__19608;
    wire N__19605;
    wire N__19602;
    wire N__19599;
    wire N__19592;
    wire N__19589;
    wire N__19588;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19573;
    wire N__19568;
    wire N__19565;
    wire N__19564;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19549;
    wire N__19544;
    wire N__19541;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19495;
    wire N__19494;
    wire N__19491;
    wire N__19488;
    wire N__19485;
    wire N__19480;
    wire N__19475;
    wire N__19472;
    wire N__19471;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19456;
    wire N__19451;
    wire N__19448;
    wire N__19447;
    wire N__19446;
    wire N__19443;
    wire N__19440;
    wire N__19437;
    wire N__19434;
    wire N__19427;
    wire N__19424;
    wire N__19423;
    wire N__19422;
    wire N__19419;
    wire N__19416;
    wire N__19413;
    wire N__19410;
    wire N__19403;
    wire N__19400;
    wire N__19399;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19384;
    wire N__19379;
    wire N__19376;
    wire N__19375;
    wire N__19374;
    wire N__19371;
    wire N__19368;
    wire N__19365;
    wire N__19360;
    wire N__19355;
    wire N__19352;
    wire N__19351;
    wire N__19350;
    wire N__19347;
    wire N__19342;
    wire N__19337;
    wire N__19334;
    wire N__19333;
    wire N__19332;
    wire N__19329;
    wire N__19324;
    wire N__19319;
    wire N__19316;
    wire N__19315;
    wire N__19314;
    wire N__19311;
    wire N__19306;
    wire N__19301;
    wire N__19298;
    wire N__19297;
    wire N__19296;
    wire N__19293;
    wire N__19290;
    wire N__19287;
    wire N__19282;
    wire N__19277;
    wire N__19274;
    wire N__19273;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19258;
    wire N__19253;
    wire N__19250;
    wire N__19249;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19229;
    wire N__19226;
    wire N__19225;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19205;
    wire N__19202;
    wire N__19201;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19186;
    wire N__19181;
    wire N__19178;
    wire N__19177;
    wire N__19176;
    wire N__19173;
    wire N__19170;
    wire N__19167;
    wire N__19162;
    wire N__19157;
    wire N__19154;
    wire N__19153;
    wire N__19152;
    wire N__19149;
    wire N__19144;
    wire N__19139;
    wire N__19136;
    wire N__19135;
    wire N__19134;
    wire N__19131;
    wire N__19126;
    wire N__19121;
    wire N__19118;
    wire N__19117;
    wire N__19116;
    wire N__19115;
    wire N__19114;
    wire N__19113;
    wire N__19112;
    wire N__19111;
    wire N__19110;
    wire N__19109;
    wire N__19108;
    wire N__19107;
    wire N__19106;
    wire N__19105;
    wire N__19104;
    wire N__19103;
    wire N__19102;
    wire N__19101;
    wire N__19100;
    wire N__19099;
    wire N__19098;
    wire N__19097;
    wire N__19096;
    wire N__19095;
    wire N__19094;
    wire N__19093;
    wire N__19092;
    wire N__19089;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19081;
    wire N__19078;
    wire N__19077;
    wire N__19074;
    wire N__19073;
    wire N__19072;
    wire N__19055;
    wire N__19038;
    wire N__19021;
    wire N__19004;
    wire N__18995;
    wire N__18994;
    wire N__18993;
    wire N__18992;
    wire N__18991;
    wire N__18990;
    wire N__18989;
    wire N__18988;
    wire N__18987;
    wire N__18986;
    wire N__18985;
    wire N__18984;
    wire N__18983;
    wire N__18982;
    wire N__18981;
    wire N__18980;
    wire N__18979;
    wire N__18978;
    wire N__18965;
    wire N__18954;
    wire N__18949;
    wire N__18938;
    wire N__18929;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18896;
    wire N__18893;
    wire N__18892;
    wire N__18889;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18869;
    wire N__18868;
    wire N__18867;
    wire N__18866;
    wire N__18865;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18847;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18830;
    wire N__18827;
    wire N__18826;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18816;
    wire N__18809;
    wire N__18806;
    wire N__18805;
    wire N__18804;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18790;
    wire N__18785;
    wire N__18782;
    wire N__18781;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18766;
    wire N__18761;
    wire N__18758;
    wire N__18757;
    wire N__18756;
    wire N__18753;
    wire N__18748;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18736;
    wire N__18735;
    wire N__18732;
    wire N__18729;
    wire N__18726;
    wire N__18721;
    wire N__18718;
    wire N__18715;
    wire N__18710;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18692;
    wire N__18691;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18674;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18659;
    wire N__18658;
    wire N__18655;
    wire N__18652;
    wire N__18647;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18635;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18623;
    wire N__18622;
    wire N__18619;
    wire N__18616;
    wire N__18611;
    wire N__18610;
    wire N__18609;
    wire N__18608;
    wire N__18607;
    wire N__18606;
    wire N__18605;
    wire N__18604;
    wire N__18603;
    wire N__18602;
    wire N__18601;
    wire N__18600;
    wire N__18599;
    wire N__18598;
    wire N__18593;
    wire N__18586;
    wire N__18573;
    wire N__18566;
    wire N__18557;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18545;
    wire N__18544;
    wire N__18541;
    wire N__18538;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18520;
    wire N__18517;
    wire N__18514;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18499;
    wire N__18496;
    wire N__18493;
    wire N__18492;
    wire N__18491;
    wire N__18488;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18467;
    wire N__18464;
    wire N__18459;
    wire N__18456;
    wire N__18451;
    wire N__18446;
    wire N__18443;
    wire N__18442;
    wire N__18439;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18429;
    wire N__18422;
    wire N__18419;
    wire N__18418;
    wire N__18415;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18405;
    wire N__18398;
    wire N__18395;
    wire N__18394;
    wire N__18393;
    wire N__18392;
    wire N__18389;
    wire N__18388;
    wire N__18387;
    wire N__18384;
    wire N__18379;
    wire N__18376;
    wire N__18371;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18349;
    wire N__18348;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18337;
    wire N__18336;
    wire N__18335;
    wire N__18334;
    wire N__18333;
    wire N__18332;
    wire N__18331;
    wire N__18330;
    wire N__18329;
    wire N__18328;
    wire N__18327;
    wire N__18326;
    wire N__18325;
    wire N__18324;
    wire N__18323;
    wire N__18322;
    wire N__18321;
    wire N__18318;
    wire N__18317;
    wire N__18316;
    wire N__18309;
    wire N__18302;
    wire N__18285;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18267;
    wire N__18262;
    wire N__18255;
    wire N__18248;
    wire N__18245;
    wire N__18236;
    wire N__18235;
    wire N__18234;
    wire N__18233;
    wire N__18232;
    wire N__18231;
    wire N__18230;
    wire N__18229;
    wire N__18228;
    wire N__18227;
    wire N__18226;
    wire N__18225;
    wire N__18224;
    wire N__18223;
    wire N__18222;
    wire N__18221;
    wire N__18220;
    wire N__18219;
    wire N__18218;
    wire N__18217;
    wire N__18216;
    wire N__18215;
    wire N__18212;
    wire N__18211;
    wire N__18198;
    wire N__18181;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18163;
    wire N__18158;
    wire N__18155;
    wire N__18146;
    wire N__18143;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18109;
    wire N__18106;
    wire N__18103;
    wire N__18102;
    wire N__18101;
    wire N__18098;
    wire N__18091;
    wire N__18088;
    wire N__18085;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18061;
    wire N__18060;
    wire N__18057;
    wire N__18052;
    wire N__18051;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18039;
    wire N__18032;
    wire N__18031;
    wire N__18028;
    wire N__18025;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18010;
    wire N__18007;
    wire N__18004;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17989;
    wire N__17986;
    wire N__17983;
    wire N__17978;
    wire N__17975;
    wire N__17972;
    wire N__17969;
    wire N__17968;
    wire N__17965;
    wire N__17962;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17947;
    wire N__17944;
    wire N__17941;
    wire N__17936;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17926;
    wire N__17923;
    wire N__17920;
    wire N__17917;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17902;
    wire N__17899;
    wire N__17896;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17878;
    wire N__17875;
    wire N__17872;
    wire N__17867;
    wire N__17866;
    wire N__17863;
    wire N__17860;
    wire N__17855;
    wire N__17852;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17827;
    wire N__17824;
    wire N__17821;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17807;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17765;
    wire N__17764;
    wire N__17761;
    wire N__17758;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17737;
    wire N__17734;
    wire N__17731;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17689;
    wire N__17686;
    wire N__17683;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17644;
    wire N__17641;
    wire N__17638;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17602;
    wire N__17599;
    wire N__17596;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17581;
    wire N__17578;
    wire N__17575;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17560;
    wire N__17559;
    wire N__17558;
    wire N__17557;
    wire N__17556;
    wire N__17553;
    wire N__17550;
    wire N__17547;
    wire N__17544;
    wire N__17543;
    wire N__17542;
    wire N__17541;
    wire N__17540;
    wire N__17539;
    wire N__17536;
    wire N__17533;
    wire N__17532;
    wire N__17531;
    wire N__17530;
    wire N__17529;
    wire N__17528;
    wire N__17527;
    wire N__17526;
    wire N__17525;
    wire N__17516;
    wire N__17509;
    wire N__17508;
    wire N__17507;
    wire N__17506;
    wire N__17501;
    wire N__17496;
    wire N__17479;
    wire N__17474;
    wire N__17471;
    wire N__17470;
    wire N__17469;
    wire N__17466;
    wire N__17463;
    wire N__17460;
    wire N__17453;
    wire N__17446;
    wire N__17435;
    wire N__17432;
    wire N__17431;
    wire N__17430;
    wire N__17429;
    wire N__17428;
    wire N__17427;
    wire N__17426;
    wire N__17425;
    wire N__17422;
    wire N__17407;
    wire N__17406;
    wire N__17405;
    wire N__17404;
    wire N__17403;
    wire N__17402;
    wire N__17401;
    wire N__17400;
    wire N__17399;
    wire N__17398;
    wire N__17397;
    wire N__17396;
    wire N__17395;
    wire N__17394;
    wire N__17391;
    wire N__17388;
    wire N__17373;
    wire N__17372;
    wire N__17371;
    wire N__17370;
    wire N__17367;
    wire N__17364;
    wire N__17355;
    wire N__17352;
    wire N__17347;
    wire N__17340;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17311;
    wire N__17308;
    wire N__17305;
    wire N__17300;
    wire N__17297;
    wire N__17294;
    wire N__17291;
    wire N__17290;
    wire N__17287;
    wire N__17284;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17249;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17237;
    wire N__17234;
    wire N__17231;
    wire N__17228;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17203;
    wire N__17200;
    wire N__17197;
    wire N__17192;
    wire N__17189;
    wire N__17186;
    wire N__17183;
    wire N__17180;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17135;
    wire N__17132;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17120;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17096;
    wire N__17095;
    wire N__17092;
    wire N__17087;
    wire N__17084;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17072;
    wire N__17071;
    wire N__17068;
    wire N__17067;
    wire N__17064;
    wire N__17061;
    wire N__17058;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17014;
    wire N__17011;
    wire N__17008;
    wire N__17003;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16981;
    wire N__16978;
    wire N__16975;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16939;
    wire N__16936;
    wire N__16933;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16915;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16834;
    wire N__16833;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16813;
    wire N__16810;
    wire N__16807;
    wire N__16802;
    wire N__16799;
    wire N__16798;
    wire N__16797;
    wire N__16796;
    wire N__16795;
    wire N__16794;
    wire N__16793;
    wire N__16792;
    wire N__16789;
    wire N__16786;
    wire N__16783;
    wire N__16774;
    wire N__16769;
    wire N__16762;
    wire N__16759;
    wire N__16754;
    wire N__16751;
    wire N__16748;
    wire N__16747;
    wire N__16746;
    wire N__16743;
    wire N__16740;
    wire N__16737;
    wire N__16732;
    wire N__16729;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16717;
    wire N__16714;
    wire N__16711;
    wire N__16710;
    wire N__16705;
    wire N__16702;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16683;
    wire N__16678;
    wire N__16675;
    wire N__16670;
    wire N__16667;
    wire N__16666;
    wire N__16663;
    wire N__16662;
    wire N__16659;
    wire N__16656;
    wire N__16653;
    wire N__16650;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16634;
    wire N__16633;
    wire N__16630;
    wire N__16627;
    wire N__16622;
    wire N__16619;
    wire N__16618;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16597;
    wire N__16596;
    wire N__16593;
    wire N__16590;
    wire N__16587;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16573;
    wire N__16572;
    wire N__16569;
    wire N__16566;
    wire N__16563;
    wire N__16556;
    wire N__16553;
    wire N__16550;
    wire N__16549;
    wire N__16548;
    wire N__16545;
    wire N__16540;
    wire N__16535;
    wire N__16532;
    wire N__16531;
    wire N__16528;
    wire N__16525;
    wire N__16524;
    wire N__16521;
    wire N__16516;
    wire N__16511;
    wire N__16508;
    wire N__16507;
    wire N__16504;
    wire N__16503;
    wire N__16500;
    wire N__16497;
    wire N__16494;
    wire N__16493;
    wire N__16490;
    wire N__16485;
    wire N__16482;
    wire N__16475;
    wire N__16472;
    wire N__16469;
    wire N__16468;
    wire N__16467;
    wire N__16464;
    wire N__16459;
    wire N__16454;
    wire N__16451;
    wire N__16450;
    wire N__16449;
    wire N__16446;
    wire N__16441;
    wire N__16438;
    wire N__16435;
    wire N__16430;
    wire N__16427;
    wire N__16426;
    wire N__16425;
    wire N__16422;
    wire N__16419;
    wire N__16416;
    wire N__16413;
    wire N__16408;
    wire N__16403;
    wire N__16400;
    wire N__16399;
    wire N__16396;
    wire N__16393;
    wire N__16392;
    wire N__16389;
    wire N__16386;
    wire N__16383;
    wire N__16378;
    wire N__16373;
    wire N__16370;
    wire N__16367;
    wire N__16366;
    wire N__16361;
    wire N__16358;
    wire N__16357;
    wire N__16354;
    wire N__16351;
    wire N__16346;
    wire N__16345;
    wire N__16344;
    wire N__16339;
    wire N__16336;
    wire N__16331;
    wire N__16328;
    wire N__16325;
    wire N__16322;
    wire N__16319;
    wire N__16316;
    wire N__16315;
    wire N__16312;
    wire N__16309;
    wire N__16304;
    wire N__16301;
    wire N__16300;
    wire N__16297;
    wire N__16294;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16284;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16263;
    wire N__16258;
    wire N__16255;
    wire N__16250;
    wire N__16247;
    wire N__16244;
    wire N__16241;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16226;
    wire N__16223;
    wire N__16220;
    wire N__16217;
    wire N__16216;
    wire N__16211;
    wire N__16208;
    wire N__16205;
    wire N__16202;
    wire N__16199;
    wire N__16196;
    wire N__16195;
    wire N__16194;
    wire N__16191;
    wire N__16190;
    wire N__16187;
    wire N__16186;
    wire N__16185;
    wire N__16178;
    wire N__16175;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16163;
    wire N__16160;
    wire N__16155;
    wire N__16148;
    wire N__16147;
    wire N__16146;
    wire N__16143;
    wire N__16140;
    wire N__16139;
    wire N__16138;
    wire N__16135;
    wire N__16130;
    wire N__16127;
    wire N__16124;
    wire N__16121;
    wire N__16118;
    wire N__16113;
    wire N__16106;
    wire N__16103;
    wire N__16102;
    wire N__16099;
    wire N__16096;
    wire N__16095;
    wire N__16094;
    wire N__16093;
    wire N__16090;
    wire N__16087;
    wire N__16082;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16070;
    wire N__16061;
    wire N__16060;
    wire N__16059;
    wire N__16056;
    wire N__16055;
    wire N__16052;
    wire N__16049;
    wire N__16046;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16018;
    wire N__16013;
    wire N__16010;
    wire N__16009;
    wire N__16008;
    wire N__16007;
    wire N__16006;
    wire N__16003;
    wire N__16000;
    wire N__15997;
    wire N__15994;
    wire N__15991;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15974;
    wire N__15965;
    wire N__15962;
    wire N__15961;
    wire N__15960;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15952;
    wire N__15949;
    wire N__15946;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15920;
    wire N__15917;
    wire N__15916;
    wire N__15915;
    wire N__15908;
    wire N__15907;
    wire N__15906;
    wire N__15905;
    wire N__15904;
    wire N__15903;
    wire N__15900;
    wire N__15897;
    wire N__15896;
    wire N__15895;
    wire N__15894;
    wire N__15893;
    wire N__15892;
    wire N__15889;
    wire N__15886;
    wire N__15885;
    wire N__15884;
    wire N__15883;
    wire N__15882;
    wire N__15877;
    wire N__15876;
    wire N__15875;
    wire N__15874;
    wire N__15873;
    wire N__15872;
    wire N__15871;
    wire N__15866;
    wire N__15861;
    wire N__15856;
    wire N__15847;
    wire N__15844;
    wire N__15839;
    wire N__15838;
    wire N__15835;
    wire N__15824;
    wire N__15821;
    wire N__15814;
    wire N__15807;
    wire N__15804;
    wire N__15797;
    wire N__15792;
    wire N__15785;
    wire N__15784;
    wire N__15783;
    wire N__15780;
    wire N__15779;
    wire N__15778;
    wire N__15775;
    wire N__15772;
    wire N__15769;
    wire N__15766;
    wire N__15763;
    wire N__15760;
    wire N__15757;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15737;
    wire N__15736;
    wire N__15735;
    wire N__15734;
    wire N__15733;
    wire N__15732;
    wire N__15731;
    wire N__15730;
    wire N__15729;
    wire N__15726;
    wire N__15723;
    wire N__15720;
    wire N__15717;
    wire N__15716;
    wire N__15715;
    wire N__15714;
    wire N__15711;
    wire N__15710;
    wire N__15707;
    wire N__15704;
    wire N__15703;
    wire N__15702;
    wire N__15701;
    wire N__15700;
    wire N__15699;
    wire N__15698;
    wire N__15691;
    wire N__15678;
    wire N__15673;
    wire N__15666;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15653;
    wire N__15652;
    wire N__15651;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15637;
    wire N__15634;
    wire N__15633;
    wire N__15618;
    wire N__15615;
    wire N__15608;
    wire N__15605;
    wire N__15602;
    wire N__15599;
    wire N__15596;
    wire N__15587;
    wire N__15586;
    wire N__15581;
    wire N__15580;
    wire N__15579;
    wire N__15578;
    wire N__15577;
    wire N__15576;
    wire N__15573;
    wire N__15566;
    wire N__15563;
    wire N__15562;
    wire N__15561;
    wire N__15560;
    wire N__15559;
    wire N__15558;
    wire N__15555;
    wire N__15554;
    wire N__15553;
    wire N__15548;
    wire N__15545;
    wire N__15534;
    wire N__15533;
    wire N__15532;
    wire N__15531;
    wire N__15530;
    wire N__15527;
    wire N__15522;
    wire N__15515;
    wire N__15506;
    wire N__15497;
    wire N__15494;
    wire N__15491;
    wire N__15488;
    wire N__15485;
    wire N__15482;
    wire N__15479;
    wire N__15476;
    wire N__15473;
    wire N__15470;
    wire N__15467;
    wire N__15466;
    wire N__15465;
    wire N__15464;
    wire N__15463;
    wire N__15462;
    wire N__15457;
    wire N__15456;
    wire N__15455;
    wire N__15454;
    wire N__15453;
    wire N__15452;
    wire N__15451;
    wire N__15450;
    wire N__15449;
    wire N__15440;
    wire N__15439;
    wire N__15438;
    wire N__15437;
    wire N__15436;
    wire N__15435;
    wire N__15434;
    wire N__15431;
    wire N__15420;
    wire N__15413;
    wire N__15412;
    wire N__15411;
    wire N__15408;
    wire N__15395;
    wire N__15388;
    wire N__15383;
    wire N__15374;
    wire N__15373;
    wire N__15370;
    wire N__15367;
    wire N__15362;
    wire N__15361;
    wire N__15360;
    wire N__15359;
    wire N__15358;
    wire N__15357;
    wire N__15356;
    wire N__15355;
    wire N__15354;
    wire N__15353;
    wire N__15352;
    wire N__15351;
    wire N__15350;
    wire N__15349;
    wire N__15346;
    wire N__15337;
    wire N__15334;
    wire N__15333;
    wire N__15332;
    wire N__15331;
    wire N__15330;
    wire N__15329;
    wire N__15318;
    wire N__15311;
    wire N__15310;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15290;
    wire N__15285;
    wire N__15280;
    wire N__15269;
    wire N__15266;
    wire N__15263;
    wire N__15262;
    wire N__15261;
    wire N__15260;
    wire N__15259;
    wire N__15258;
    wire N__15257;
    wire N__15256;
    wire N__15255;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15238;
    wire N__15237;
    wire N__15236;
    wire N__15235;
    wire N__15234;
    wire N__15233;
    wire N__15232;
    wire N__15231;
    wire N__15230;
    wire N__15229;
    wire N__15228;
    wire N__15227;
    wire N__15224;
    wire N__15215;
    wire N__15212;
    wire N__15203;
    wire N__15200;
    wire N__15197;
    wire N__15190;
    wire N__15175;
    wire N__15172;
    wire N__15171;
    wire N__15170;
    wire N__15165;
    wire N__15158;
    wire N__15153;
    wire N__15150;
    wire N__15147;
    wire N__15144;
    wire N__15141;
    wire N__15138;
    wire N__15131;
    wire N__15122;
    wire N__15119;
    wire N__15118;
    wire N__15115;
    wire N__15112;
    wire N__15111;
    wire N__15106;
    wire N__15103;
    wire N__15102;
    wire N__15101;
    wire N__15098;
    wire N__15095;
    wire N__15090;
    wire N__15083;
    wire N__15080;
    wire N__15079;
    wire N__15078;
    wire N__15077;
    wire N__15076;
    wire N__15075;
    wire N__15074;
    wire N__15073;
    wire N__15072;
    wire N__15071;
    wire N__15070;
    wire N__15069;
    wire N__15068;
    wire N__15067;
    wire N__15066;
    wire N__15065;
    wire N__15064;
    wire N__15063;
    wire N__15062;
    wire N__15061;
    wire N__15058;
    wire N__15053;
    wire N__15036;
    wire N__15033;
    wire N__15016;
    wire N__15009;
    wire N__15008;
    wire N__15003;
    wire N__15002;
    wire N__15001;
    wire N__14998;
    wire N__14997;
    wire N__14994;
    wire N__14991;
    wire N__14988;
    wire N__14985;
    wire N__14982;
    wire N__14979;
    wire N__14976;
    wire N__14971;
    wire N__14960;
    wire N__14957;
    wire N__14954;
    wire N__14953;
    wire N__14950;
    wire N__14947;
    wire N__14946;
    wire N__14945;
    wire N__14942;
    wire N__14937;
    wire N__14934;
    wire N__14927;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14902;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14876;
    wire N__14875;
    wire N__14874;
    wire N__14873;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14852;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14840;
    wire N__14831;
    wire N__14830;
    wire N__14829;
    wire N__14828;
    wire N__14825;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14815;
    wire N__14814;
    wire N__14811;
    wire N__14808;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14789;
    wire N__14786;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14731;
    wire N__14730;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14722;
    wire N__14719;
    wire N__14716;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14684;
    wire N__14683;
    wire N__14682;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14666;
    wire N__14665;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14652;
    wire N__14651;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14625;
    wire N__14618;
    wire N__14617;
    wire N__14616;
    wire N__14615;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14605;
    wire N__14602;
    wire N__14599;
    wire N__14596;
    wire N__14593;
    wire N__14588;
    wire N__14585;
    wire N__14580;
    wire N__14577;
    wire N__14570;
    wire N__14569;
    wire N__14566;
    wire N__14565;
    wire N__14562;
    wire N__14559;
    wire N__14558;
    wire N__14555;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14530;
    wire N__14525;
    wire N__14520;
    wire N__14515;
    wire N__14510;
    wire N__14509;
    wire N__14508;
    wire N__14507;
    wire N__14504;
    wire N__14501;
    wire N__14498;
    wire N__14497;
    wire N__14494;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14475;
    wire N__14472;
    wire N__14469;
    wire N__14466;
    wire N__14459;
    wire N__14458;
    wire N__14457;
    wire N__14454;
    wire N__14451;
    wire N__14450;
    wire N__14449;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14428;
    wire N__14425;
    wire N__14422;
    wire N__14419;
    wire N__14416;
    wire N__14413;
    wire N__14410;
    wire N__14399;
    wire N__14398;
    wire N__14397;
    wire N__14394;
    wire N__14393;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14385;
    wire N__14382;
    wire N__14379;
    wire N__14376;
    wire N__14373;
    wire N__14370;
    wire N__14367;
    wire N__14360;
    wire N__14355;
    wire N__14352;
    wire N__14349;
    wire N__14346;
    wire N__14339;
    wire N__14338;
    wire N__14337;
    wire N__14334;
    wire N__14333;
    wire N__14332;
    wire N__14329;
    wire N__14326;
    wire N__14323;
    wire N__14320;
    wire N__14317;
    wire N__14308;
    wire N__14305;
    wire N__14302;
    wire N__14297;
    wire N__14294;
    wire N__14291;
    wire N__14288;
    wire N__14285;
    wire N__14282;
    wire N__14279;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14264;
    wire N__14263;
    wire N__14262;
    wire N__14259;
    wire N__14256;
    wire N__14253;
    wire N__14252;
    wire N__14251;
    wire N__14246;
    wire N__14243;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14229;
    wire N__14222;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14214;
    wire N__14211;
    wire N__14208;
    wire N__14207;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14197;
    wire N__14192;
    wire N__14189;
    wire N__14186;
    wire N__14183;
    wire N__14180;
    wire N__14171;
    wire N__14170;
    wire N__14169;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14153;
    wire N__14150;
    wire N__14149;
    wire N__14148;
    wire N__14143;
    wire N__14140;
    wire N__14137;
    wire N__14132;
    wire N__14129;
    wire N__14126;
    wire N__14123;
    wire N__14122;
    wire N__14121;
    wire N__14120;
    wire N__14117;
    wire N__14114;
    wire N__14111;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14090;
    wire N__14087;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14075;
    wire N__14072;
    wire N__14069;
    wire N__14066;
    wire N__14063;
    wire N__14060;
    wire N__14057;
    wire N__14054;
    wire N__14051;
    wire N__14048;
    wire N__14045;
    wire N__14042;
    wire N__14039;
    wire N__14036;
    wire N__14033;
    wire N__14030;
    wire N__14027;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13997;
    wire N__13994;
    wire N__13991;
    wire N__13988;
    wire N__13985;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13967;
    wire N__13964;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13937;
    wire N__13934;
    wire N__13931;
    wire N__13928;
    wire N__13925;
    wire N__13922;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13844;
    wire N__13841;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13826;
    wire N__13823;
    wire N__13822;
    wire N__13819;
    wire N__13816;
    wire N__13813;
    wire N__13812;
    wire N__13809;
    wire N__13806;
    wire N__13803;
    wire N__13800;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13784;
    wire N__13783;
    wire N__13782;
    wire N__13779;
    wire N__13776;
    wire N__13773;
    wire N__13770;
    wire N__13769;
    wire N__13766;
    wire N__13763;
    wire N__13760;
    wire N__13757;
    wire N__13754;
    wire N__13749;
    wire N__13746;
    wire N__13739;
    wire N__13736;
    wire N__13733;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13723;
    wire N__13720;
    wire N__13719;
    wire N__13718;
    wire N__13715;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13690;
    wire N__13687;
    wire N__13684;
    wire N__13681;
    wire N__13678;
    wire N__13677;
    wire N__13676;
    wire N__13671;
    wire N__13668;
    wire N__13665;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13648;
    wire N__13645;
    wire N__13644;
    wire N__13641;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13631;
    wire N__13628;
    wire N__13623;
    wire N__13616;
    wire N__13613;
    wire N__13610;
    wire N__13607;
    wire N__13606;
    wire N__13605;
    wire N__13604;
    wire N__13595;
    wire N__13592;
    wire N__13591;
    wire N__13590;
    wire N__13589;
    wire N__13588;
    wire N__13585;
    wire N__13576;
    wire N__13573;
    wire N__13570;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13523;
    wire N__13520;
    wire N__13517;
    wire N__13514;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13415;
    wire N__13412;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13391;
    wire N__13388;
    wire N__13385;
    wire N__13382;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13367;
    wire N__13364;
    wire N__13361;
    wire N__13358;
    wire N__13355;
    wire N__13354;
    wire N__13353;
    wire N__13350;
    wire N__13347;
    wire N__13344;
    wire N__13337;
    wire N__13336;
    wire N__13331;
    wire N__13328;
    wire N__13327;
    wire N__13326;
    wire N__13325;
    wire N__13322;
    wire N__13317;
    wire N__13314;
    wire N__13307;
    wire N__13306;
    wire N__13303;
    wire N__13302;
    wire N__13301;
    wire N__13294;
    wire N__13293;
    wire N__13290;
    wire N__13289;
    wire N__13286;
    wire N__13279;
    wire N__13276;
    wire N__13273;
    wire N__13268;
    wire N__13267;
    wire N__13266;
    wire N__13265;
    wire N__13264;
    wire N__13263;
    wire N__13256;
    wire N__13249;
    wire N__13246;
    wire N__13243;
    wire N__13240;
    wire N__13235;
    wire N__13234;
    wire N__13233;
    wire N__13232;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13224;
    wire N__13221;
    wire N__13218;
    wire N__13213;
    wire N__13208;
    wire N__13205;
    wire N__13200;
    wire N__13195;
    wire N__13192;
    wire N__13187;
    wire N__13184;
    wire N__13183;
    wire N__13180;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13170;
    wire N__13167;
    wire N__13162;
    wire N__13157;
    wire N__13156;
    wire N__13155;
    wire N__13154;
    wire N__13153;
    wire N__13146;
    wire N__13141;
    wire N__13140;
    wire N__13139;
    wire N__13138;
    wire N__13137;
    wire N__13136;
    wire N__13133;
    wire N__13130;
    wire N__13119;
    wire N__13118;
    wire N__13115;
    wire N__13110;
    wire N__13107;
    wire N__13100;
    wire N__13097;
    wire N__13094;
    wire N__13091;
    wire N__13088;
    wire N__13085;
    wire N__13082;
    wire N__13079;
    wire N__13076;
    wire N__13073;
    wire N__13070;
    wire N__13067;
    wire N__13064;
    wire N__13061;
    wire N__13058;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13040;
    wire N__13037;
    wire N__13034;
    wire N__13031;
    wire N__13028;
    wire N__13025;
    wire N__13022;
    wire N__13019;
    wire N__13016;
    wire N__13015;
    wire N__13012;
    wire N__13009;
    wire N__13008;
    wire N__13003;
    wire N__13000;
    wire N__12995;
    wire N__12994;
    wire N__12991;
    wire N__12988;
    wire N__12987;
    wire N__12984;
    wire N__12981;
    wire N__12978;
    wire N__12975;
    wire N__12972;
    wire N__12969;
    wire N__12962;
    wire N__12961;
    wire N__12958;
    wire N__12957;
    wire N__12956;
    wire N__12953;
    wire N__12952;
    wire N__12949;
    wire N__12944;
    wire N__12941;
    wire N__12938;
    wire N__12933;
    wire N__12926;
    wire N__12925;
    wire N__12924;
    wire N__12923;
    wire N__12922;
    wire N__12911;
    wire N__12910;
    wire N__12907;
    wire N__12906;
    wire N__12905;
    wire N__12904;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12886;
    wire N__12881;
    wire N__12880;
    wire N__12877;
    wire N__12874;
    wire N__12873;
    wire N__12870;
    wire N__12867;
    wire N__12864;
    wire N__12857;
    wire N__12856;
    wire N__12853;
    wire N__12850;
    wire N__12847;
    wire N__12844;
    wire N__12843;
    wire N__12840;
    wire N__12837;
    wire N__12834;
    wire N__12827;
    wire N__12824;
    wire N__12823;
    wire N__12822;
    wire N__12819;
    wire N__12818;
    wire N__12817;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12803;
    wire N__12800;
    wire N__12795;
    wire N__12792;
    wire N__12789;
    wire N__12782;
    wire N__12779;
    wire N__12778;
    wire N__12777;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12764;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12743;
    wire N__12740;
    wire N__12739;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12724;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12712;
    wire N__12709;
    wire N__12706;
    wire N__12701;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12691;
    wire N__12688;
    wire N__12685;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12668;
    wire N__12665;
    wire N__12662;
    wire N__12659;
    wire N__12656;
    wire N__12655;
    wire N__12652;
    wire N__12649;
    wire N__12644;
    wire N__12641;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12626;
    wire N__12623;
    wire N__12620;
    wire N__12617;
    wire N__12614;
    wire N__12611;
    wire N__12610;
    wire N__12607;
    wire N__12604;
    wire N__12603;
    wire N__12600;
    wire N__12597;
    wire N__12594;
    wire N__12587;
    wire N__12586;
    wire N__12583;
    wire N__12580;
    wire N__12577;
    wire N__12574;
    wire N__12571;
    wire N__12568;
    wire N__12567;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12555;
    wire N__12548;
    wire N__12545;
    wire N__12544;
    wire N__12541;
    wire N__12538;
    wire N__12537;
    wire N__12536;
    wire N__12535;
    wire N__12532;
    wire N__12529;
    wire N__12522;
    wire N__12515;
    wire N__12514;
    wire N__12511;
    wire N__12508;
    wire N__12503;
    wire N__12500;
    wire N__12499;
    wire N__12498;
    wire N__12497;
    wire N__12496;
    wire N__12495;
    wire N__12492;
    wire N__12489;
    wire N__12486;
    wire N__12485;
    wire N__12484;
    wire N__12483;
    wire N__12482;
    wire N__12481;
    wire N__12480;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12469;
    wire N__12468;
    wire N__12467;
    wire N__12466;
    wire N__12465;
    wire N__12464;
    wire N__12457;
    wire N__12448;
    wire N__12441;
    wire N__12434;
    wire N__12427;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12417;
    wire N__12416;
    wire N__12415;
    wire N__12414;
    wire N__12407;
    wire N__12400;
    wire N__12397;
    wire N__12396;
    wire N__12393;
    wire N__12388;
    wire N__12383;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12359;
    wire N__12358;
    wire N__12357;
    wire N__12356;
    wire N__12355;
    wire N__12354;
    wire N__12353;
    wire N__12352;
    wire N__12351;
    wire N__12350;
    wire N__12349;
    wire N__12348;
    wire N__12347;
    wire N__12346;
    wire N__12345;
    wire N__12344;
    wire N__12343;
    wire N__12342;
    wire N__12341;
    wire N__12326;
    wire N__12319;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12296;
    wire N__12295;
    wire N__12294;
    wire N__12293;
    wire N__12288;
    wire N__12283;
    wire N__12280;
    wire N__12279;
    wire N__12274;
    wire N__12267;
    wire N__12262;
    wire N__12259;
    wire N__12256;
    wire N__12245;
    wire N__12242;
    wire N__12241;
    wire N__12240;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12230;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12194;
    wire N__12191;
    wire N__12188;
    wire N__12185;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12173;
    wire N__12170;
    wire N__12167;
    wire N__12164;
    wire N__12161;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12151;
    wire N__12146;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12133;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12123;
    wire N__12118;
    wire N__12113;
    wire N__12110;
    wire N__12109;
    wire N__12108;
    wire N__12105;
    wire N__12102;
    wire N__12099;
    wire N__12094;
    wire N__12089;
    wire N__12086;
    wire N__12085;
    wire N__12084;
    wire N__12081;
    wire N__12078;
    wire N__12075;
    wire N__12072;
    wire N__12065;
    wire N__12062;
    wire N__12061;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12051;
    wire N__12048;
    wire N__12041;
    wire N__12038;
    wire N__12037;
    wire N__12036;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12022;
    wire N__12017;
    wire N__12014;
    wire N__12013;
    wire N__12012;
    wire N__12009;
    wire N__12006;
    wire N__12003;
    wire N__11998;
    wire N__11993;
    wire N__11990;
    wire N__11989;
    wire N__11986;
    wire N__11983;
    wire N__11978;
    wire N__11975;
    wire N__11974;
    wire N__11973;
    wire N__11972;
    wire N__11971;
    wire N__11970;
    wire N__11969;
    wire N__11968;
    wire N__11967;
    wire N__11966;
    wire N__11965;
    wire N__11964;
    wire N__11963;
    wire N__11962;
    wire N__11961;
    wire N__11960;
    wire N__11959;
    wire N__11958;
    wire N__11957;
    wire N__11956;
    wire N__11955;
    wire N__11954;
    wire N__11953;
    wire N__11952;
    wire N__11951;
    wire N__11950;
    wire N__11949;
    wire N__11948;
    wire N__11947;
    wire N__11946;
    wire N__11937;
    wire N__11928;
    wire N__11923;
    wire N__11914;
    wire N__11905;
    wire N__11896;
    wire N__11887;
    wire N__11878;
    wire N__11875;
    wire N__11860;
    wire N__11855;
    wire N__11852;
    wire N__11851;
    wire N__11848;
    wire N__11845;
    wire N__11840;
    wire N__11839;
    wire N__11838;
    wire N__11837;
    wire N__11828;
    wire N__11825;
    wire N__11822;
    wire N__11821;
    wire N__11820;
    wire N__11817;
    wire N__11812;
    wire N__11807;
    wire N__11804;
    wire N__11803;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11788;
    wire N__11783;
    wire N__11780;
    wire N__11779;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11764;
    wire N__11759;
    wire N__11756;
    wire N__11755;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11735;
    wire N__11732;
    wire N__11731;
    wire N__11730;
    wire N__11727;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11711;
    wire N__11708;
    wire N__11707;
    wire N__11706;
    wire N__11703;
    wire N__11700;
    wire N__11697;
    wire N__11692;
    wire N__11687;
    wire N__11684;
    wire N__11683;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11673;
    wire N__11668;
    wire N__11663;
    wire N__11660;
    wire N__11659;
    wire N__11658;
    wire N__11655;
    wire N__11650;
    wire N__11645;
    wire N__11642;
    wire N__11641;
    wire N__11640;
    wire N__11637;
    wire N__11632;
    wire N__11627;
    wire N__11626;
    wire N__11625;
    wire N__11622;
    wire N__11617;
    wire N__11612;
    wire N__11609;
    wire N__11608;
    wire N__11607;
    wire N__11604;
    wire N__11601;
    wire N__11598;
    wire N__11593;
    wire N__11588;
    wire N__11585;
    wire N__11584;
    wire N__11583;
    wire N__11580;
    wire N__11577;
    wire N__11574;
    wire N__11569;
    wire N__11564;
    wire N__11561;
    wire N__11560;
    wire N__11559;
    wire N__11556;
    wire N__11553;
    wire N__11550;
    wire N__11543;
    wire N__11540;
    wire N__11539;
    wire N__11538;
    wire N__11535;
    wire N__11532;
    wire N__11529;
    wire N__11526;
    wire N__11519;
    wire N__11516;
    wire N__11515;
    wire N__11514;
    wire N__11511;
    wire N__11508;
    wire N__11505;
    wire N__11500;
    wire N__11495;
    wire N__11492;
    wire N__11491;
    wire N__11490;
    wire N__11487;
    wire N__11484;
    wire N__11481;
    wire N__11476;
    wire N__11471;
    wire N__11468;
    wire N__11467;
    wire N__11466;
    wire N__11463;
    wire N__11458;
    wire N__11453;
    wire N__11450;
    wire N__11449;
    wire N__11448;
    wire N__11445;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11429;
    wire N__11428;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11416;
    wire N__11413;
    wire N__11410;
    wire N__11405;
    wire N__11404;
    wire N__11401;
    wire N__11400;
    wire N__11397;
    wire N__11392;
    wire N__11389;
    wire N__11386;
    wire N__11381;
    wire N__11380;
    wire N__11379;
    wire N__11378;
    wire N__11377;
    wire N__11370;
    wire N__11365;
    wire N__11364;
    wire N__11363;
    wire N__11362;
    wire N__11361;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11347;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11331;
    wire N__11324;
    wire N__11323;
    wire N__11322;
    wire N__11321;
    wire N__11320;
    wire N__11315;
    wire N__11308;
    wire N__11303;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11282;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11274;
    wire N__11271;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11256;
    wire N__11249;
    wire N__11246;
    wire N__11243;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11235;
    wire N__11232;
    wire N__11229;
    wire N__11226;
    wire N__11219;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11209;
    wire N__11208;
    wire N__11205;
    wire N__11202;
    wire N__11199;
    wire N__11192;
    wire N__11189;
    wire N__11188;
    wire N__11187;
    wire N__11184;
    wire N__11181;
    wire N__11178;
    wire N__11173;
    wire N__11168;
    wire N__11165;
    wire N__11164;
    wire N__11163;
    wire N__11160;
    wire N__11157;
    wire N__11154;
    wire N__11149;
    wire N__11144;
    wire N__11141;
    wire N__11140;
    wire N__11139;
    wire N__11136;
    wire N__11131;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11098;
    wire N__11095;
    wire N__11094;
    wire N__11091;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11079;
    wire N__11072;
    wire N__11071;
    wire N__11070;
    wire N__11069;
    wire N__11068;
    wire N__11067;
    wire N__11066;
    wire N__11061;
    wire N__11060;
    wire N__11049;
    wire N__11046;
    wire N__11043;
    wire N__11036;
    wire N__11035;
    wire N__11034;
    wire N__11033;
    wire N__11032;
    wire N__11031;
    wire N__11030;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11018;
    wire N__11007;
    wire N__11000;
    wire N__10999;
    wire N__10998;
    wire N__10995;
    wire N__10992;
    wire N__10991;
    wire N__10990;
    wire N__10987;
    wire N__10986;
    wire N__10983;
    wire N__10972;
    wire N__10969;
    wire N__10966;
    wire N__10961;
    wire N__10960;
    wire N__10957;
    wire N__10954;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10907;
    wire N__10904;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10726;
    wire N__10725;
    wire N__10724;
    wire N__10723;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10613;
    wire N__10610;
    wire N__10609;
    wire N__10606;
    wire N__10603;
    wire N__10600;
    wire N__10597;
    wire N__10592;
    wire N__10589;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10571;
    wire N__10568;
    wire N__10565;
    wire N__10564;
    wire N__10563;
    wire N__10562;
    wire N__10561;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10544;
    wire N__10537;
    wire N__10532;
    wire N__10529;
    wire N__10528;
    wire N__10525;
    wire N__10524;
    wire N__10521;
    wire N__10520;
    wire N__10519;
    wire N__10518;
    wire N__10513;
    wire N__10510;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10492;
    wire N__10489;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10477;
    wire N__10476;
    wire N__10473;
    wire N__10468;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10456;
    wire N__10455;
    wire N__10452;
    wire N__10449;
    wire N__10448;
    wire N__10443;
    wire N__10440;
    wire N__10437;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10423;
    wire N__10420;
    wire N__10417;
    wire N__10412;
    wire N__10411;
    wire N__10408;
    wire N__10405;
    wire N__10404;
    wire N__10401;
    wire N__10398;
    wire N__10395;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10360;
    wire N__10357;
    wire N__10354;
    wire N__10353;
    wire N__10350;
    wire N__10347;
    wire N__10344;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10330;
    wire N__10329;
    wire N__10326;
    wire N__10323;
    wire N__10320;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10303;
    wire N__10302;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10286;
    wire N__10283;
    wire N__10282;
    wire N__10279;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10255;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10238;
    wire N__10235;
    wire N__10232;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10222;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10210;
    wire N__10207;
    wire N__10204;
    wire N__10201;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10189;
    wire N__10186;
    wire N__10183;
    wire N__10180;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10168;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10156;
    wire N__10153;
    wire N__10152;
    wire N__10149;
    wire N__10146;
    wire N__10143;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10114;
    wire N__10111;
    wire N__10108;
    wire N__10105;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10093;
    wire N__10090;
    wire N__10087;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10066;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10054;
    wire N__10051;
    wire N__10048;
    wire N__10045;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10033;
    wire N__10030;
    wire N__10027;
    wire N__10024;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9916;
    wire N__9913;
    wire N__9910;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9895;
    wire N__9892;
    wire N__9889;
    wire N__9886;
    wire N__9883;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9865;
    wire N__9862;
    wire N__9859;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9841;
    wire N__9838;
    wire N__9835;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9793;
    wire N__9790;
    wire N__9787;
    wire N__9782;
    wire N__9779;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9727;
    wire N__9724;
    wire N__9721;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9703;
    wire N__9700;
    wire N__9697;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9608;
    wire N__9605;
    wire N__9604;
    wire N__9601;
    wire N__9598;
    wire N__9593;
    wire N__9592;
    wire N__9591;
    wire N__9586;
    wire N__9583;
    wire N__9580;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9313;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9274;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9262;
    wire N__9259;
    wire N__9256;
    wire N__9253;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9025;
    wire N__9022;
    wire N__9019;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__9001;
    wire N__8998;
    wire N__8995;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8977;
    wire N__8974;
    wire N__8971;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8911;
    wire N__8908;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8898;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8872;
    wire N__8869;
    wire N__8866;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8758;
    wire N__8757;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire GNDG0;
    wire VCCG0;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0 ;
    wire bfn_1_18_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_1_19_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire bfn_1_20_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire N_27_i_i;
    wire un7_start_stop;
    wire CONSTANT_ONE_NET;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_1 ;
    wire bfn_2_15_0_;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_9 ;
    wire bfn_2_16_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_17 ;
    wire bfn_2_17_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_ ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ;
    wire bfn_2_22_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ;
    wire bfn_2_23_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire bfn_2_24_0_;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \delay_measurement_inst.N_212_cascade_ ;
    wire \delay_measurement_inst.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5_cascade_ ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19 ;
    wire bfn_3_19_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_8 ;
    wire bfn_3_20_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_16 ;
    wire bfn_3_21_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \delay_measurement_inst.N_168 ;
    wire \delay_measurement_inst.N_81_i ;
    wire \delay_measurement_inst.N_81_i_cascade_ ;
    wire \delay_measurement_inst.N_200 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_ ;
    wire \delay_measurement_inst.un1_tr_state_1_i_0_a2_0_7 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_203 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_2 ;
    wire \delay_measurement_inst.elapsed_time_tr_3 ;
    wire bfn_4_15_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.elapsed_time_tr_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.elapsed_time_tr_11 ;
    wire bfn_4_16_0_;
    wire \delay_measurement_inst.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.elapsed_time_tr_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.elapsed_time_tr_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire bfn_4_17_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_4_18_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_138_i_g ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_0 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_15_cascade_ ;
    wire il_max_comp2_c;
    wire il_max_comp2_D1;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_4Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_6Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.N_92_cascade_ ;
    wire \delay_measurement_inst.elapsed_time_tr_9 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ;
    wire \delay_measurement_inst.N_165 ;
    wire \delay_measurement_inst.N_212 ;
    wire \delay_measurement_inst.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.elapsed_time_tr_19 ;
    wire \delay_measurement_inst.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ;
    wire \delay_measurement_inst.N_197_1 ;
    wire \delay_measurement_inst.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.N_81_i_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire bfn_5_15_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_5_16_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_5_17_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_5_18_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_139_i_g ;
    wire \phase_controller_inst1.stoper_hc.un1_m3_eZ0Z_1 ;
    wire phase_controller_inst1_stoper_hc_un1_startlto19_2;
    wire phase_controller_inst1_stoper_hc_un1_startlto19_2_cascade_;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto31_a0Z0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto31_aZ0Z2_cascade_ ;
    wire d_N_5_mux;
    wire \phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_2_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_N_6_mux ;
    wire \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_m2_eZ0 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30_2_0Z0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire measured_delay_tr_11;
    wire measured_delay_tr_9;
    wire \phase_controller_inst1.stoper_tr.N_98 ;
    wire measured_delay_tr_12;
    wire measured_delay_tr_13;
    wire measured_delay_tr_14;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ;
    wire measured_delay_tr_10;
    wire measured_delay_tr_4;
    wire measured_delay_tr_7;
    wire measured_delay_tr_8;
    wire measured_delay_tr_5;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ;
    wire measured_delay_tr_1;
    wire measured_delay_tr_2;
    wire measured_delay_tr_3;
    wire \phase_controller_inst1.stoper_tr.N_109 ;
    wire \phase_controller_inst1.stoper_tr.N_110 ;
    wire \phase_controller_inst1.stoper_tr.N_92 ;
    wire measured_delay_tr_6;
    wire \phase_controller_inst1.stoper_tr.N_95 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_7_14_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_7_15_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_17 ;
    wire bfn_7_16_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_ ;
    wire \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ;
    wire measured_delay_tr_19;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire measured_delay_tr_17;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire measured_delay_tr_18;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire measured_delay_tr_16;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlt31 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ;
    wire bfn_7_19_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire bfn_7_20_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_16 ;
    wire bfn_7_21_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.time_passed11_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire measured_delay_hc_4;
    wire measured_delay_hc_1;
    wire measured_delay_hc_22;
    wire measured_delay_hc_21;
    wire measured_delay_hc_0;
    wire measured_delay_hc_5;
    wire measured_delay_hc_20;
    wire measured_delay_hc_3;
    wire measured_delay_hc_17;
    wire measured_delay_hc_6;
    wire measured_delay_hc_13;
    wire measured_delay_hc_19;
    wire measured_delay_hc_15;
    wire measured_delay_hc_18;
    wire measured_delay_hc_16;
    wire measured_delay_hc_14;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_0_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_0_0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ;
    wire il_min_comp2_c;
    wire \phase_controller_slave.stoper_tr.time_passed11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_inst1.stoper_tr.time_passed11_cascade_ ;
    wire \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_slave.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.un1_start ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto31_d ;
    wire \phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire measured_delay_hc_9;
    wire measured_delay_hc_7;
    wire measured_delay_hc_2;
    wire measured_delay_hc_8;
    wire measured_delay_hc_12;
    wire measured_delay_hc_10;
    wire measured_delay_hc_31;
    wire measured_delay_hc_11;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5FBM1Z0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_2 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2Z0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2Z0Z_6_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_3 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_2 ;
    wire \delay_measurement_inst.elapsed_time_hc_3 ;
    wire bfn_8_26_0_;
    wire \delay_measurement_inst.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_reg3lto6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_reg3lto9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.elapsed_time_hc_11 ;
    wire bfn_8_27_0_;
    wire \delay_measurement_inst.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_reg3lto14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_reg3lto15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.elapsed_time_hc_19 ;
    wire bfn_8_28_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire bfn_8_29_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ;
    wire bfn_9_13_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ;
    wire bfn_9_14_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ;
    wire bfn_9_15_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ;
    wire bfn_9_17_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ;
    wire bfn_9_18_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ;
    wire bfn_9_19_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.time_passed11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_slave.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_slave.N_21 ;
    wire s3_phy_c;
    wire \phase_controller_slave.stoper_hc.time_passed11 ;
    wire \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4 ;
    wire measured_delay_hc_30;
    wire measured_delay_hc_24;
    wire measured_delay_hc_25;
    wire measured_delay_hc_28;
    wire measured_delay_hc_29;
    wire \delay_measurement_inst.delay_hc_reg3 ;
    wire measured_delay_hc_23;
    wire measured_delay_hc_27;
    wire \delay_measurement_inst.un1_elapsed_time_hc ;
    wire \delay_measurement_inst.delay_hc_reg3lto31_0_0 ;
    wire measured_delay_hc_26;
    wire \delay_measurement_inst.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.N_136_i_g ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_9_26_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_9_27_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_9_28_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_9_29_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_138_i ;
    wire il_max_comp1_c;
    wire il_max_comp1_D1;
    wire il_min_comp1_c;
    wire il_min_comp1_D1;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ;
    wire measured_delay_tr_15;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ;
    wire \phase_controller_slave.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ;
    wire \phase_controller_inst1.stoper_tr.time_passed11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_slave.start_timer_tr_0_sqmuxa ;
    wire il_min_comp2_D1;
    wire \phase_controller_slave.N_20 ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.T01_0_sqmuxa ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.N_83 ;
    wire il_max_comp1_D2;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_slave.tr_time_passed ;
    wire \phase_controller_slave.stateZ0Z_0 ;
    wire shift_flag_start;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst1.N_88 ;
    wire il_max_comp2_D2;
    wire \phase_controller_slave.stateZ0Z_4 ;
    wire \phase_controller_slave.un1_startZ0 ;
    wire \phase_controller_slave.stateZ0Z_3 ;
    wire il_min_comp2_D2;
    wire \phase_controller_slave.stateZ0Z_2 ;
    wire \phase_controller_slave.hc_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire \phase_controller_slave.stateZ0Z_1 ;
    wire s4_phy_c;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.un1_tr_state_1_i_0_0 ;
    wire start_stop_c;
    wire \phase_controller_inst1.stateZ0Z_4 ;
    wire \phase_controller_inst1.N_86 ;
    wire \delay_measurement_inst.delay_hc_timer.N_137_i_g ;
    wire \phase_controller_inst1.stateZ0Z_3 ;
    wire s1_phy_c;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_139_i ;
    wire delay_tr_input_c;
    wire delay_tr_d1;
    wire delay_tr_d2;
    wire \delay_measurement_inst.prev_tr_sigZ0 ;
    wire \delay_measurement_inst.tr_stateZ0Z_0 ;
    wire red_c_i;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire delay_hc_input_c;
    wire delay_hc_d1;
    wire \delay_measurement_inst.prev_hc_sigZ0 ;
    wire \delay_measurement_inst.hc_stateZ0Z_0 ;
    wire red_c_g;
    wire delay_hc_d2;
    wire clk_100mhz;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.N_136_i ;
    wire _gnd_net_;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__12626),
            .RESETB(N__21350),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__22542),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__22544),
            .DIN(N__22543),
            .DOUT(N__22542),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__22544),
            .PADOUT(N__22543),
            .PADIN(N__22542),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__22533),
            .DIN(N__22532),
            .DOUT(N__22531),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__22533),
            .PADOUT(N__22532),
            .PADIN(N__22531),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__22524),
            .DIN(N__22523),
            .DOUT(N__22522),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__22524),
            .PADOUT(N__22523),
            .PADIN(N__22522),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21530),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__22515),
            .DIN(N__22514),
            .DOUT(N__22513),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__22515),
            .PADOUT(N__22514),
            .PADIN(N__22513),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21092),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__22506),
            .DIN(N__22505),
            .DOUT(N__22504),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__22506),
            .PADOUT(N__22505),
            .PADIN(N__22504),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__22497),
            .DIN(N__22496),
            .DOUT(N__22495),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__22497),
            .PADOUT(N__22496),
            .PADIN(N__22495),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__22488),
            .DIN(N__22487),
            .DOUT(N__22486),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__22488),
            .PADOUT(N__22487),
            .PADIN(N__22486),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__22479),
            .DIN(N__22478),
            .DOUT(N__22477),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__22479),
            .PADOUT(N__22478),
            .PADIN(N__22477),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__22470),
            .DIN(N__22469),
            .DOUT(N__22468),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__22470),
            .PADOUT(N__22469),
            .PADIN(N__22468),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__22461),
            .DIN(N__22460),
            .DOUT(N__22459),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__22461),
            .PADOUT(N__22460),
            .PADIN(N__22459),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21149),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__22452),
            .DIN(N__22451),
            .DOUT(N__22450),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__22452),
            .PADOUT(N__22451),
            .PADIN(N__22450),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18119),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_iopad (
            .OE(N__22443),
            .DIN(N__22442),
            .DOUT(N__22441),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_preio (
            .PADOEN(N__22443),
            .PADOUT(N__22442),
            .PADIN(N__22441),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_iopad (
            .OE(N__22434),
            .DIN(N__22433),
            .DOUT(N__22432),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_preio (
            .PADOEN(N__22434),
            .PADOUT(N__22433),
            .PADIN(N__22432),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__5331 (
            .O(N__22415),
            .I(N__22411));
    InMux I__5330 (
            .O(N__22414),
            .I(N__22408));
    LocalMux I__5329 (
            .O(N__22411),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    LocalMux I__5328 (
            .O(N__22408),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__5327 (
            .O(N__22403),
            .I(N__22400));
    LocalMux I__5326 (
            .O(N__22400),
            .I(N__22397));
    Span12Mux_h I__5325 (
            .O(N__22397),
            .I(N__22394));
    Span12Mux_v I__5324 (
            .O(N__22394),
            .I(N__22391));
    Odrv12 I__5323 (
            .O(N__22391),
            .I(delay_hc_input_c));
    InMux I__5322 (
            .O(N__22388),
            .I(N__22385));
    LocalMux I__5321 (
            .O(N__22385),
            .I(N__22382));
    Odrv12 I__5320 (
            .O(N__22382),
            .I(delay_hc_d1));
    InMux I__5319 (
            .O(N__22379),
            .I(N__22374));
    InMux I__5318 (
            .O(N__22378),
            .I(N__22371));
    InMux I__5317 (
            .O(N__22377),
            .I(N__22368));
    LocalMux I__5316 (
            .O(N__22374),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__5315 (
            .O(N__22371),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__5314 (
            .O(N__22368),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    InMux I__5313 (
            .O(N__22361),
            .I(N__22356));
    InMux I__5312 (
            .O(N__22360),
            .I(N__22353));
    InMux I__5311 (
            .O(N__22359),
            .I(N__22350));
    LocalMux I__5310 (
            .O(N__22356),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__5309 (
            .O(N__22353),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__5308 (
            .O(N__22350),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    CascadeMux I__5307 (
            .O(N__22343),
            .I(N__22336));
    InMux I__5306 (
            .O(N__22342),
            .I(N__22332));
    InMux I__5305 (
            .O(N__22341),
            .I(N__22329));
    InMux I__5304 (
            .O(N__22340),
            .I(N__22326));
    InMux I__5303 (
            .O(N__22339),
            .I(N__22323));
    InMux I__5302 (
            .O(N__22336),
            .I(N__22320));
    InMux I__5301 (
            .O(N__22335),
            .I(N__22317));
    LocalMux I__5300 (
            .O(N__22332),
            .I(N__22314));
    LocalMux I__5299 (
            .O(N__22329),
            .I(N__22311));
    LocalMux I__5298 (
            .O(N__22326),
            .I(N__22308));
    LocalMux I__5297 (
            .O(N__22323),
            .I(N__22305));
    LocalMux I__5296 (
            .O(N__22320),
            .I(N__22266));
    LocalMux I__5295 (
            .O(N__22317),
            .I(N__22244));
    Glb2LocalMux I__5294 (
            .O(N__22314),
            .I(N__22082));
    Glb2LocalMux I__5293 (
            .O(N__22311),
            .I(N__22082));
    Glb2LocalMux I__5292 (
            .O(N__22308),
            .I(N__22082));
    Glb2LocalMux I__5291 (
            .O(N__22305),
            .I(N__22082));
    SRMux I__5290 (
            .O(N__22304),
            .I(N__22082));
    SRMux I__5289 (
            .O(N__22303),
            .I(N__22082));
    SRMux I__5288 (
            .O(N__22302),
            .I(N__22082));
    SRMux I__5287 (
            .O(N__22301),
            .I(N__22082));
    SRMux I__5286 (
            .O(N__22300),
            .I(N__22082));
    SRMux I__5285 (
            .O(N__22299),
            .I(N__22082));
    SRMux I__5284 (
            .O(N__22298),
            .I(N__22082));
    SRMux I__5283 (
            .O(N__22297),
            .I(N__22082));
    SRMux I__5282 (
            .O(N__22296),
            .I(N__22082));
    SRMux I__5281 (
            .O(N__22295),
            .I(N__22082));
    SRMux I__5280 (
            .O(N__22294),
            .I(N__22082));
    SRMux I__5279 (
            .O(N__22293),
            .I(N__22082));
    SRMux I__5278 (
            .O(N__22292),
            .I(N__22082));
    SRMux I__5277 (
            .O(N__22291),
            .I(N__22082));
    SRMux I__5276 (
            .O(N__22290),
            .I(N__22082));
    SRMux I__5275 (
            .O(N__22289),
            .I(N__22082));
    SRMux I__5274 (
            .O(N__22288),
            .I(N__22082));
    SRMux I__5273 (
            .O(N__22287),
            .I(N__22082));
    SRMux I__5272 (
            .O(N__22286),
            .I(N__22082));
    SRMux I__5271 (
            .O(N__22285),
            .I(N__22082));
    SRMux I__5270 (
            .O(N__22284),
            .I(N__22082));
    SRMux I__5269 (
            .O(N__22283),
            .I(N__22082));
    SRMux I__5268 (
            .O(N__22282),
            .I(N__22082));
    SRMux I__5267 (
            .O(N__22281),
            .I(N__22082));
    SRMux I__5266 (
            .O(N__22280),
            .I(N__22082));
    SRMux I__5265 (
            .O(N__22279),
            .I(N__22082));
    SRMux I__5264 (
            .O(N__22278),
            .I(N__22082));
    SRMux I__5263 (
            .O(N__22277),
            .I(N__22082));
    SRMux I__5262 (
            .O(N__22276),
            .I(N__22082));
    SRMux I__5261 (
            .O(N__22275),
            .I(N__22082));
    SRMux I__5260 (
            .O(N__22274),
            .I(N__22082));
    SRMux I__5259 (
            .O(N__22273),
            .I(N__22082));
    SRMux I__5258 (
            .O(N__22272),
            .I(N__22082));
    SRMux I__5257 (
            .O(N__22271),
            .I(N__22082));
    SRMux I__5256 (
            .O(N__22270),
            .I(N__22082));
    SRMux I__5255 (
            .O(N__22269),
            .I(N__22082));
    Glb2LocalMux I__5254 (
            .O(N__22266),
            .I(N__22082));
    SRMux I__5253 (
            .O(N__22265),
            .I(N__22082));
    SRMux I__5252 (
            .O(N__22264),
            .I(N__22082));
    SRMux I__5251 (
            .O(N__22263),
            .I(N__22082));
    SRMux I__5250 (
            .O(N__22262),
            .I(N__22082));
    SRMux I__5249 (
            .O(N__22261),
            .I(N__22082));
    SRMux I__5248 (
            .O(N__22260),
            .I(N__22082));
    SRMux I__5247 (
            .O(N__22259),
            .I(N__22082));
    SRMux I__5246 (
            .O(N__22258),
            .I(N__22082));
    SRMux I__5245 (
            .O(N__22257),
            .I(N__22082));
    SRMux I__5244 (
            .O(N__22256),
            .I(N__22082));
    SRMux I__5243 (
            .O(N__22255),
            .I(N__22082));
    SRMux I__5242 (
            .O(N__22254),
            .I(N__22082));
    SRMux I__5241 (
            .O(N__22253),
            .I(N__22082));
    SRMux I__5240 (
            .O(N__22252),
            .I(N__22082));
    SRMux I__5239 (
            .O(N__22251),
            .I(N__22082));
    SRMux I__5238 (
            .O(N__22250),
            .I(N__22082));
    SRMux I__5237 (
            .O(N__22249),
            .I(N__22082));
    SRMux I__5236 (
            .O(N__22248),
            .I(N__22082));
    SRMux I__5235 (
            .O(N__22247),
            .I(N__22082));
    Glb2LocalMux I__5234 (
            .O(N__22244),
            .I(N__22082));
    SRMux I__5233 (
            .O(N__22243),
            .I(N__22082));
    SRMux I__5232 (
            .O(N__22242),
            .I(N__22082));
    SRMux I__5231 (
            .O(N__22241),
            .I(N__22082));
    SRMux I__5230 (
            .O(N__22240),
            .I(N__22082));
    SRMux I__5229 (
            .O(N__22239),
            .I(N__22082));
    SRMux I__5228 (
            .O(N__22238),
            .I(N__22082));
    SRMux I__5227 (
            .O(N__22237),
            .I(N__22082));
    SRMux I__5226 (
            .O(N__22236),
            .I(N__22082));
    SRMux I__5225 (
            .O(N__22235),
            .I(N__22082));
    SRMux I__5224 (
            .O(N__22234),
            .I(N__22082));
    SRMux I__5223 (
            .O(N__22233),
            .I(N__22082));
    SRMux I__5222 (
            .O(N__22232),
            .I(N__22082));
    SRMux I__5221 (
            .O(N__22231),
            .I(N__22082));
    GlobalMux I__5220 (
            .O(N__22082),
            .I(N__22079));
    gio2CtrlBuf I__5219 (
            .O(N__22079),
            .I(red_c_g));
    InMux I__5218 (
            .O(N__22076),
            .I(N__22072));
    InMux I__5217 (
            .O(N__22075),
            .I(N__22067));
    LocalMux I__5216 (
            .O(N__22072),
            .I(N__22064));
    InMux I__5215 (
            .O(N__22071),
            .I(N__22061));
    InMux I__5214 (
            .O(N__22070),
            .I(N__22058));
    LocalMux I__5213 (
            .O(N__22067),
            .I(N__22051));
    Span4Mux_v I__5212 (
            .O(N__22064),
            .I(N__22051));
    LocalMux I__5211 (
            .O(N__22061),
            .I(N__22051));
    LocalMux I__5210 (
            .O(N__22058),
            .I(N__22048));
    Odrv4 I__5209 (
            .O(N__22051),
            .I(delay_hc_d2));
    Odrv12 I__5208 (
            .O(N__22048),
            .I(delay_hc_d2));
    ClkMux I__5207 (
            .O(N__22043),
            .I(N__21788));
    ClkMux I__5206 (
            .O(N__22042),
            .I(N__21788));
    ClkMux I__5205 (
            .O(N__22041),
            .I(N__21788));
    ClkMux I__5204 (
            .O(N__22040),
            .I(N__21788));
    ClkMux I__5203 (
            .O(N__22039),
            .I(N__21788));
    ClkMux I__5202 (
            .O(N__22038),
            .I(N__21788));
    ClkMux I__5201 (
            .O(N__22037),
            .I(N__21788));
    ClkMux I__5200 (
            .O(N__22036),
            .I(N__21788));
    ClkMux I__5199 (
            .O(N__22035),
            .I(N__21788));
    ClkMux I__5198 (
            .O(N__22034),
            .I(N__21788));
    ClkMux I__5197 (
            .O(N__22033),
            .I(N__21788));
    ClkMux I__5196 (
            .O(N__22032),
            .I(N__21788));
    ClkMux I__5195 (
            .O(N__22031),
            .I(N__21788));
    ClkMux I__5194 (
            .O(N__22030),
            .I(N__21788));
    ClkMux I__5193 (
            .O(N__22029),
            .I(N__21788));
    ClkMux I__5192 (
            .O(N__22028),
            .I(N__21788));
    ClkMux I__5191 (
            .O(N__22027),
            .I(N__21788));
    ClkMux I__5190 (
            .O(N__22026),
            .I(N__21788));
    ClkMux I__5189 (
            .O(N__22025),
            .I(N__21788));
    ClkMux I__5188 (
            .O(N__22024),
            .I(N__21788));
    ClkMux I__5187 (
            .O(N__22023),
            .I(N__21788));
    ClkMux I__5186 (
            .O(N__22022),
            .I(N__21788));
    ClkMux I__5185 (
            .O(N__22021),
            .I(N__21788));
    ClkMux I__5184 (
            .O(N__22020),
            .I(N__21788));
    ClkMux I__5183 (
            .O(N__22019),
            .I(N__21788));
    ClkMux I__5182 (
            .O(N__22018),
            .I(N__21788));
    ClkMux I__5181 (
            .O(N__22017),
            .I(N__21788));
    ClkMux I__5180 (
            .O(N__22016),
            .I(N__21788));
    ClkMux I__5179 (
            .O(N__22015),
            .I(N__21788));
    ClkMux I__5178 (
            .O(N__22014),
            .I(N__21788));
    ClkMux I__5177 (
            .O(N__22013),
            .I(N__21788));
    ClkMux I__5176 (
            .O(N__22012),
            .I(N__21788));
    ClkMux I__5175 (
            .O(N__22011),
            .I(N__21788));
    ClkMux I__5174 (
            .O(N__22010),
            .I(N__21788));
    ClkMux I__5173 (
            .O(N__22009),
            .I(N__21788));
    ClkMux I__5172 (
            .O(N__22008),
            .I(N__21788));
    ClkMux I__5171 (
            .O(N__22007),
            .I(N__21788));
    ClkMux I__5170 (
            .O(N__22006),
            .I(N__21788));
    ClkMux I__5169 (
            .O(N__22005),
            .I(N__21788));
    ClkMux I__5168 (
            .O(N__22004),
            .I(N__21788));
    ClkMux I__5167 (
            .O(N__22003),
            .I(N__21788));
    ClkMux I__5166 (
            .O(N__22002),
            .I(N__21788));
    ClkMux I__5165 (
            .O(N__22001),
            .I(N__21788));
    ClkMux I__5164 (
            .O(N__22000),
            .I(N__21788));
    ClkMux I__5163 (
            .O(N__21999),
            .I(N__21788));
    ClkMux I__5162 (
            .O(N__21998),
            .I(N__21788));
    ClkMux I__5161 (
            .O(N__21997),
            .I(N__21788));
    ClkMux I__5160 (
            .O(N__21996),
            .I(N__21788));
    ClkMux I__5159 (
            .O(N__21995),
            .I(N__21788));
    ClkMux I__5158 (
            .O(N__21994),
            .I(N__21788));
    ClkMux I__5157 (
            .O(N__21993),
            .I(N__21788));
    ClkMux I__5156 (
            .O(N__21992),
            .I(N__21788));
    ClkMux I__5155 (
            .O(N__21991),
            .I(N__21788));
    ClkMux I__5154 (
            .O(N__21990),
            .I(N__21788));
    ClkMux I__5153 (
            .O(N__21989),
            .I(N__21788));
    ClkMux I__5152 (
            .O(N__21988),
            .I(N__21788));
    ClkMux I__5151 (
            .O(N__21987),
            .I(N__21788));
    ClkMux I__5150 (
            .O(N__21986),
            .I(N__21788));
    ClkMux I__5149 (
            .O(N__21985),
            .I(N__21788));
    ClkMux I__5148 (
            .O(N__21984),
            .I(N__21788));
    ClkMux I__5147 (
            .O(N__21983),
            .I(N__21788));
    ClkMux I__5146 (
            .O(N__21982),
            .I(N__21788));
    ClkMux I__5145 (
            .O(N__21981),
            .I(N__21788));
    ClkMux I__5144 (
            .O(N__21980),
            .I(N__21788));
    ClkMux I__5143 (
            .O(N__21979),
            .I(N__21788));
    ClkMux I__5142 (
            .O(N__21978),
            .I(N__21788));
    ClkMux I__5141 (
            .O(N__21977),
            .I(N__21788));
    ClkMux I__5140 (
            .O(N__21976),
            .I(N__21788));
    ClkMux I__5139 (
            .O(N__21975),
            .I(N__21788));
    ClkMux I__5138 (
            .O(N__21974),
            .I(N__21788));
    ClkMux I__5137 (
            .O(N__21973),
            .I(N__21788));
    ClkMux I__5136 (
            .O(N__21972),
            .I(N__21788));
    ClkMux I__5135 (
            .O(N__21971),
            .I(N__21788));
    ClkMux I__5134 (
            .O(N__21970),
            .I(N__21788));
    ClkMux I__5133 (
            .O(N__21969),
            .I(N__21788));
    ClkMux I__5132 (
            .O(N__21968),
            .I(N__21788));
    ClkMux I__5131 (
            .O(N__21967),
            .I(N__21788));
    ClkMux I__5130 (
            .O(N__21966),
            .I(N__21788));
    ClkMux I__5129 (
            .O(N__21965),
            .I(N__21788));
    ClkMux I__5128 (
            .O(N__21964),
            .I(N__21788));
    ClkMux I__5127 (
            .O(N__21963),
            .I(N__21788));
    ClkMux I__5126 (
            .O(N__21962),
            .I(N__21788));
    ClkMux I__5125 (
            .O(N__21961),
            .I(N__21788));
    ClkMux I__5124 (
            .O(N__21960),
            .I(N__21788));
    ClkMux I__5123 (
            .O(N__21959),
            .I(N__21788));
    GlobalMux I__5122 (
            .O(N__21788),
            .I(clk_100mhz));
    InMux I__5121 (
            .O(N__21785),
            .I(N__21782));
    LocalMux I__5120 (
            .O(N__21782),
            .I(N__21778));
    InMux I__5119 (
            .O(N__21781),
            .I(N__21774));
    Span4Mux_h I__5118 (
            .O(N__21778),
            .I(N__21771));
    InMux I__5117 (
            .O(N__21777),
            .I(N__21768));
    LocalMux I__5116 (
            .O(N__21774),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv4 I__5115 (
            .O(N__21771),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    LocalMux I__5114 (
            .O(N__21768),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__5113 (
            .O(N__21761),
            .I(N__21756));
    InMux I__5112 (
            .O(N__21760),
            .I(N__21752));
    InMux I__5111 (
            .O(N__21759),
            .I(N__21749));
    LocalMux I__5110 (
            .O(N__21756),
            .I(N__21746));
    InMux I__5109 (
            .O(N__21755),
            .I(N__21743));
    LocalMux I__5108 (
            .O(N__21752),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__5107 (
            .O(N__21749),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__5106 (
            .O(N__21746),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__5105 (
            .O(N__21743),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    IoInMux I__5104 (
            .O(N__21734),
            .I(N__21731));
    LocalMux I__5103 (
            .O(N__21731),
            .I(N__21728));
    Odrv12 I__5102 (
            .O(N__21728),
            .I(\delay_measurement_inst.delay_hc_timer.N_136_i ));
    InMux I__5101 (
            .O(N__21725),
            .I(N__21722));
    LocalMux I__5100 (
            .O(N__21722),
            .I(N__21718));
    InMux I__5099 (
            .O(N__21721),
            .I(N__21715));
    Span4Mux_s1_v I__5098 (
            .O(N__21718),
            .I(N__21710));
    LocalMux I__5097 (
            .O(N__21715),
            .I(N__21710));
    Span4Mux_v I__5096 (
            .O(N__21710),
            .I(N__21704));
    InMux I__5095 (
            .O(N__21709),
            .I(N__21701));
    InMux I__5094 (
            .O(N__21708),
            .I(N__21698));
    InMux I__5093 (
            .O(N__21707),
            .I(N__21695));
    Span4Mux_h I__5092 (
            .O(N__21704),
            .I(N__21692));
    LocalMux I__5091 (
            .O(N__21701),
            .I(N__21687));
    LocalMux I__5090 (
            .O(N__21698),
            .I(N__21687));
    LocalMux I__5089 (
            .O(N__21695),
            .I(N__21684));
    Sp12to4 I__5088 (
            .O(N__21692),
            .I(N__21681));
    Span4Mux_v I__5087 (
            .O(N__21687),
            .I(N__21678));
    Span4Mux_h I__5086 (
            .O(N__21684),
            .I(N__21675));
    Span12Mux_v I__5085 (
            .O(N__21681),
            .I(N__21672));
    Sp12to4 I__5084 (
            .O(N__21678),
            .I(N__21669));
    Span4Mux_h I__5083 (
            .O(N__21675),
            .I(N__21666));
    Span12Mux_v I__5082 (
            .O(N__21672),
            .I(N__21663));
    Span12Mux_h I__5081 (
            .O(N__21669),
            .I(N__21660));
    Sp12to4 I__5080 (
            .O(N__21666),
            .I(N__21657));
    Span12Mux_h I__5079 (
            .O(N__21663),
            .I(N__21652));
    Span12Mux_v I__5078 (
            .O(N__21660),
            .I(N__21652));
    Span12Mux_v I__5077 (
            .O(N__21657),
            .I(N__21649));
    Odrv12 I__5076 (
            .O(N__21652),
            .I(start_stop_c));
    Odrv12 I__5075 (
            .O(N__21649),
            .I(start_stop_c));
    CascadeMux I__5074 (
            .O(N__21644),
            .I(N__21639));
    InMux I__5073 (
            .O(N__21643),
            .I(N__21630));
    InMux I__5072 (
            .O(N__21642),
            .I(N__21630));
    InMux I__5071 (
            .O(N__21639),
            .I(N__21630));
    InMux I__5070 (
            .O(N__21638),
            .I(N__21627));
    InMux I__5069 (
            .O(N__21637),
            .I(N__21624));
    LocalMux I__5068 (
            .O(N__21630),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__5067 (
            .O(N__21627),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__5066 (
            .O(N__21624),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    CascadeMux I__5065 (
            .O(N__21617),
            .I(N__21614));
    InMux I__5064 (
            .O(N__21614),
            .I(N__21611));
    LocalMux I__5063 (
            .O(N__21611),
            .I(\phase_controller_inst1.N_86 ));
    CEMux I__5062 (
            .O(N__21608),
            .I(N__21603));
    CEMux I__5061 (
            .O(N__21607),
            .I(N__21600));
    CEMux I__5060 (
            .O(N__21606),
            .I(N__21597));
    LocalMux I__5059 (
            .O(N__21603),
            .I(N__21593));
    LocalMux I__5058 (
            .O(N__21600),
            .I(N__21590));
    LocalMux I__5057 (
            .O(N__21597),
            .I(N__21587));
    CEMux I__5056 (
            .O(N__21596),
            .I(N__21584));
    Span4Mux_h I__5055 (
            .O(N__21593),
            .I(N__21581));
    Span4Mux_h I__5054 (
            .O(N__21590),
            .I(N__21578));
    Span4Mux_h I__5053 (
            .O(N__21587),
            .I(N__21575));
    LocalMux I__5052 (
            .O(N__21584),
            .I(N__21572));
    Odrv4 I__5051 (
            .O(N__21581),
            .I(\delay_measurement_inst.delay_hc_timer.N_137_i_g ));
    Odrv4 I__5050 (
            .O(N__21578),
            .I(\delay_measurement_inst.delay_hc_timer.N_137_i_g ));
    Odrv4 I__5049 (
            .O(N__21575),
            .I(\delay_measurement_inst.delay_hc_timer.N_137_i_g ));
    Odrv12 I__5048 (
            .O(N__21572),
            .I(\delay_measurement_inst.delay_hc_timer.N_137_i_g ));
    InMux I__5047 (
            .O(N__21563),
            .I(N__21560));
    LocalMux I__5046 (
            .O(N__21560),
            .I(N__21557));
    Span4Mux_v I__5045 (
            .O(N__21557),
            .I(N__21553));
    CascadeMux I__5044 (
            .O(N__21556),
            .I(N__21549));
    Span4Mux_v I__5043 (
            .O(N__21553),
            .I(N__21545));
    InMux I__5042 (
            .O(N__21552),
            .I(N__21540));
    InMux I__5041 (
            .O(N__21549),
            .I(N__21540));
    InMux I__5040 (
            .O(N__21548),
            .I(N__21537));
    Odrv4 I__5039 (
            .O(N__21545),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__5038 (
            .O(N__21540),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__5037 (
            .O(N__21537),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    IoInMux I__5036 (
            .O(N__21530),
            .I(N__21527));
    LocalMux I__5035 (
            .O(N__21527),
            .I(N__21524));
    Span4Mux_s3_v I__5034 (
            .O(N__21524),
            .I(N__21521));
    Span4Mux_h I__5033 (
            .O(N__21521),
            .I(N__21518));
    Odrv4 I__5032 (
            .O(N__21518),
            .I(s1_phy_c));
    InMux I__5031 (
            .O(N__21515),
            .I(N__21510));
    InMux I__5030 (
            .O(N__21514),
            .I(N__21507));
    InMux I__5029 (
            .O(N__21513),
            .I(N__21504));
    LocalMux I__5028 (
            .O(N__21510),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__5027 (
            .O(N__21507),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__5026 (
            .O(N__21504),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__5025 (
            .O(N__21497),
            .I(N__21493));
    InMux I__5024 (
            .O(N__21496),
            .I(N__21490));
    LocalMux I__5023 (
            .O(N__21493),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__5022 (
            .O(N__21490),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    InMux I__5021 (
            .O(N__21485),
            .I(N__21481));
    InMux I__5020 (
            .O(N__21484),
            .I(N__21476));
    LocalMux I__5019 (
            .O(N__21481),
            .I(N__21473));
    InMux I__5018 (
            .O(N__21480),
            .I(N__21470));
    InMux I__5017 (
            .O(N__21479),
            .I(N__21467));
    LocalMux I__5016 (
            .O(N__21476),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv12 I__5015 (
            .O(N__21473),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__5014 (
            .O(N__21470),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__5013 (
            .O(N__21467),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    IoInMux I__5012 (
            .O(N__21458),
            .I(N__21455));
    LocalMux I__5011 (
            .O(N__21455),
            .I(N__21452));
    Span12Mux_s2_v I__5010 (
            .O(N__21452),
            .I(N__21449));
    Odrv12 I__5009 (
            .O(N__21449),
            .I(\delay_measurement_inst.delay_tr_timer.N_139_i ));
    InMux I__5008 (
            .O(N__21446),
            .I(N__21443));
    LocalMux I__5007 (
            .O(N__21443),
            .I(N__21440));
    Span4Mux_h I__5006 (
            .O(N__21440),
            .I(N__21437));
    Span4Mux_v I__5005 (
            .O(N__21437),
            .I(N__21434));
    Span4Mux_v I__5004 (
            .O(N__21434),
            .I(N__21431));
    Odrv4 I__5003 (
            .O(N__21431),
            .I(delay_tr_input_c));
    InMux I__5002 (
            .O(N__21428),
            .I(N__21425));
    LocalMux I__5001 (
            .O(N__21425),
            .I(delay_tr_d1));
    CascadeMux I__5000 (
            .O(N__21422),
            .I(N__21415));
    InMux I__4999 (
            .O(N__21421),
            .I(N__21412));
    InMux I__4998 (
            .O(N__21420),
            .I(N__21405));
    InMux I__4997 (
            .O(N__21419),
            .I(N__21405));
    InMux I__4996 (
            .O(N__21418),
            .I(N__21405));
    InMux I__4995 (
            .O(N__21415),
            .I(N__21402));
    LocalMux I__4994 (
            .O(N__21412),
            .I(delay_tr_d2));
    LocalMux I__4993 (
            .O(N__21405),
            .I(delay_tr_d2));
    LocalMux I__4992 (
            .O(N__21402),
            .I(delay_tr_d2));
    InMux I__4991 (
            .O(N__21395),
            .I(N__21389));
    InMux I__4990 (
            .O(N__21394),
            .I(N__21384));
    InMux I__4989 (
            .O(N__21393),
            .I(N__21384));
    InMux I__4988 (
            .O(N__21392),
            .I(N__21381));
    LocalMux I__4987 (
            .O(N__21389),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__4986 (
            .O(N__21384),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__4985 (
            .O(N__21381),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    InMux I__4984 (
            .O(N__21374),
            .I(N__21368));
    InMux I__4983 (
            .O(N__21373),
            .I(N__21365));
    InMux I__4982 (
            .O(N__21372),
            .I(N__21362));
    InMux I__4981 (
            .O(N__21371),
            .I(N__21359));
    LocalMux I__4980 (
            .O(N__21368),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__4979 (
            .O(N__21365),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__4978 (
            .O(N__21362),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__4977 (
            .O(N__21359),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    IoInMux I__4976 (
            .O(N__21350),
            .I(N__21346));
    CEMux I__4975 (
            .O(N__21349),
            .I(N__21343));
    LocalMux I__4974 (
            .O(N__21346),
            .I(N__21339));
    LocalMux I__4973 (
            .O(N__21343),
            .I(N__21335));
    CEMux I__4972 (
            .O(N__21342),
            .I(N__21332));
    IoSpan4Mux I__4971 (
            .O(N__21339),
            .I(N__21328));
    CEMux I__4970 (
            .O(N__21338),
            .I(N__21325));
    Span4Mux_h I__4969 (
            .O(N__21335),
            .I(N__21319));
    LocalMux I__4968 (
            .O(N__21332),
            .I(N__21319));
    CEMux I__4967 (
            .O(N__21331),
            .I(N__21316));
    Span4Mux_s2_v I__4966 (
            .O(N__21328),
            .I(N__21312));
    LocalMux I__4965 (
            .O(N__21325),
            .I(N__21309));
    CEMux I__4964 (
            .O(N__21324),
            .I(N__21306));
    Span4Mux_v I__4963 (
            .O(N__21319),
            .I(N__21301));
    LocalMux I__4962 (
            .O(N__21316),
            .I(N__21301));
    CEMux I__4961 (
            .O(N__21315),
            .I(N__21298));
    Span4Mux_h I__4960 (
            .O(N__21312),
            .I(N__21293));
    Span4Mux_h I__4959 (
            .O(N__21309),
            .I(N__21293));
    LocalMux I__4958 (
            .O(N__21306),
            .I(N__21290));
    Span4Mux_h I__4957 (
            .O(N__21301),
            .I(N__21286));
    LocalMux I__4956 (
            .O(N__21298),
            .I(N__21283));
    Span4Mux_v I__4955 (
            .O(N__21293),
            .I(N__21278));
    Span4Mux_v I__4954 (
            .O(N__21290),
            .I(N__21278));
    CEMux I__4953 (
            .O(N__21289),
            .I(N__21275));
    Span4Mux_h I__4952 (
            .O(N__21286),
            .I(N__21270));
    Span4Mux_v I__4951 (
            .O(N__21283),
            .I(N__21270));
    Span4Mux_h I__4950 (
            .O(N__21278),
            .I(N__21267));
    LocalMux I__4949 (
            .O(N__21275),
            .I(N__21264));
    Span4Mux_v I__4948 (
            .O(N__21270),
            .I(N__21261));
    Span4Mux_h I__4947 (
            .O(N__21267),
            .I(N__21258));
    Span4Mux_v I__4946 (
            .O(N__21264),
            .I(N__21255));
    Odrv4 I__4945 (
            .O(N__21261),
            .I(red_c_i));
    Odrv4 I__4944 (
            .O(N__21258),
            .I(red_c_i));
    Odrv4 I__4943 (
            .O(N__21255),
            .I(red_c_i));
    InMux I__4942 (
            .O(N__21248),
            .I(N__21244));
    InMux I__4941 (
            .O(N__21247),
            .I(N__21241));
    LocalMux I__4940 (
            .O(N__21244),
            .I(N__21235));
    LocalMux I__4939 (
            .O(N__21241),
            .I(N__21235));
    InMux I__4938 (
            .O(N__21240),
            .I(N__21232));
    Odrv12 I__4937 (
            .O(N__21235),
            .I(il_min_comp2_D2));
    LocalMux I__4936 (
            .O(N__21232),
            .I(il_min_comp2_D2));
    CascadeMux I__4935 (
            .O(N__21227),
            .I(N__21223));
    InMux I__4934 (
            .O(N__21226),
            .I(N__21219));
    InMux I__4933 (
            .O(N__21223),
            .I(N__21216));
    InMux I__4932 (
            .O(N__21222),
            .I(N__21213));
    LocalMux I__4931 (
            .O(N__21219),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    LocalMux I__4930 (
            .O(N__21216),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    LocalMux I__4929 (
            .O(N__21213),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    InMux I__4928 (
            .O(N__21206),
            .I(N__21200));
    InMux I__4927 (
            .O(N__21205),
            .I(N__21197));
    InMux I__4926 (
            .O(N__21204),
            .I(N__21194));
    InMux I__4925 (
            .O(N__21203),
            .I(N__21191));
    LocalMux I__4924 (
            .O(N__21200),
            .I(\phase_controller_slave.hc_time_passed ));
    LocalMux I__4923 (
            .O(N__21197),
            .I(\phase_controller_slave.hc_time_passed ));
    LocalMux I__4922 (
            .O(N__21194),
            .I(\phase_controller_slave.hc_time_passed ));
    LocalMux I__4921 (
            .O(N__21191),
            .I(\phase_controller_slave.hc_time_passed ));
    InMux I__4920 (
            .O(N__21182),
            .I(N__21177));
    InMux I__4919 (
            .O(N__21181),
            .I(N__21174));
    CascadeMux I__4918 (
            .O(N__21180),
            .I(N__21171));
    LocalMux I__4917 (
            .O(N__21177),
            .I(N__21167));
    LocalMux I__4916 (
            .O(N__21174),
            .I(N__21164));
    InMux I__4915 (
            .O(N__21171),
            .I(N__21161));
    InMux I__4914 (
            .O(N__21170),
            .I(N__21158));
    Odrv12 I__4913 (
            .O(N__21167),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__4912 (
            .O(N__21164),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__4911 (
            .O(N__21161),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__4910 (
            .O(N__21158),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__4909 (
            .O(N__21149),
            .I(N__21146));
    LocalMux I__4908 (
            .O(N__21146),
            .I(N__21143));
    Span4Mux_s0_v I__4907 (
            .O(N__21143),
            .I(N__21140));
    Span4Mux_v I__4906 (
            .O(N__21140),
            .I(N__21137));
    Span4Mux_v I__4905 (
            .O(N__21137),
            .I(N__21134));
    Odrv4 I__4904 (
            .O(N__21134),
            .I(s2_phy_c));
    CascadeMux I__4903 (
            .O(N__21131),
            .I(N__21127));
    InMux I__4902 (
            .O(N__21130),
            .I(N__21122));
    InMux I__4901 (
            .O(N__21127),
            .I(N__21119));
    CascadeMux I__4900 (
            .O(N__21126),
            .I(N__21116));
    InMux I__4899 (
            .O(N__21125),
            .I(N__21113));
    LocalMux I__4898 (
            .O(N__21122),
            .I(N__21110));
    LocalMux I__4897 (
            .O(N__21119),
            .I(N__21107));
    InMux I__4896 (
            .O(N__21116),
            .I(N__21104));
    LocalMux I__4895 (
            .O(N__21113),
            .I(N__21101));
    Odrv12 I__4894 (
            .O(N__21110),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    Odrv4 I__4893 (
            .O(N__21107),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    LocalMux I__4892 (
            .O(N__21104),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    Odrv12 I__4891 (
            .O(N__21101),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    IoInMux I__4890 (
            .O(N__21092),
            .I(N__21089));
    LocalMux I__4889 (
            .O(N__21089),
            .I(N__21086));
    Span4Mux_s1_v I__4888 (
            .O(N__21086),
            .I(N__21083));
    Span4Mux_v I__4887 (
            .O(N__21083),
            .I(N__21080));
    Odrv4 I__4886 (
            .O(N__21080),
            .I(s4_phy_c));
    InMux I__4885 (
            .O(N__21077),
            .I(N__21067));
    InMux I__4884 (
            .O(N__21076),
            .I(N__21067));
    InMux I__4883 (
            .O(N__21075),
            .I(N__21046));
    InMux I__4882 (
            .O(N__21074),
            .I(N__21046));
    InMux I__4881 (
            .O(N__21073),
            .I(N__21046));
    InMux I__4880 (
            .O(N__21072),
            .I(N__21046));
    LocalMux I__4879 (
            .O(N__21067),
            .I(N__21031));
    InMux I__4878 (
            .O(N__21066),
            .I(N__21022));
    InMux I__4877 (
            .O(N__21065),
            .I(N__21022));
    InMux I__4876 (
            .O(N__21064),
            .I(N__21022));
    InMux I__4875 (
            .O(N__21063),
            .I(N__21022));
    InMux I__4874 (
            .O(N__21062),
            .I(N__21013));
    InMux I__4873 (
            .O(N__21061),
            .I(N__21013));
    InMux I__4872 (
            .O(N__21060),
            .I(N__21013));
    InMux I__4871 (
            .O(N__21059),
            .I(N__21013));
    InMux I__4870 (
            .O(N__21058),
            .I(N__21004));
    InMux I__4869 (
            .O(N__21057),
            .I(N__21004));
    InMux I__4868 (
            .O(N__21056),
            .I(N__21004));
    InMux I__4867 (
            .O(N__21055),
            .I(N__21004));
    LocalMux I__4866 (
            .O(N__21046),
            .I(N__21001));
    InMux I__4865 (
            .O(N__21045),
            .I(N__20992));
    InMux I__4864 (
            .O(N__21044),
            .I(N__20992));
    InMux I__4863 (
            .O(N__21043),
            .I(N__20992));
    InMux I__4862 (
            .O(N__21042),
            .I(N__20992));
    InMux I__4861 (
            .O(N__21041),
            .I(N__20983));
    InMux I__4860 (
            .O(N__21040),
            .I(N__20983));
    InMux I__4859 (
            .O(N__21039),
            .I(N__20983));
    InMux I__4858 (
            .O(N__21038),
            .I(N__20983));
    InMux I__4857 (
            .O(N__21037),
            .I(N__20974));
    InMux I__4856 (
            .O(N__21036),
            .I(N__20974));
    InMux I__4855 (
            .O(N__21035),
            .I(N__20974));
    InMux I__4854 (
            .O(N__21034),
            .I(N__20974));
    Span4Mux_h I__4853 (
            .O(N__21031),
            .I(N__20969));
    LocalMux I__4852 (
            .O(N__21022),
            .I(N__20969));
    LocalMux I__4851 (
            .O(N__21013),
            .I(N__20962));
    LocalMux I__4850 (
            .O(N__21004),
            .I(N__20962));
    Span4Mux_h I__4849 (
            .O(N__21001),
            .I(N__20962));
    LocalMux I__4848 (
            .O(N__20992),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__4847 (
            .O(N__20983),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__4846 (
            .O(N__20974),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__4845 (
            .O(N__20969),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__4844 (
            .O(N__20962),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__4843 (
            .O(N__20951),
            .I(N__20948));
    LocalMux I__4842 (
            .O(N__20948),
            .I(N__20932));
    InMux I__4841 (
            .O(N__20947),
            .I(N__20921));
    InMux I__4840 (
            .O(N__20946),
            .I(N__20921));
    InMux I__4839 (
            .O(N__20945),
            .I(N__20921));
    InMux I__4838 (
            .O(N__20944),
            .I(N__20921));
    InMux I__4837 (
            .O(N__20943),
            .I(N__20921));
    InMux I__4836 (
            .O(N__20942),
            .I(N__20914));
    InMux I__4835 (
            .O(N__20941),
            .I(N__20914));
    InMux I__4834 (
            .O(N__20940),
            .I(N__20914));
    InMux I__4833 (
            .O(N__20939),
            .I(N__20907));
    InMux I__4832 (
            .O(N__20938),
            .I(N__20907));
    InMux I__4831 (
            .O(N__20937),
            .I(N__20907));
    InMux I__4830 (
            .O(N__20936),
            .I(N__20902));
    InMux I__4829 (
            .O(N__20935),
            .I(N__20902));
    Span4Mux_h I__4828 (
            .O(N__20932),
            .I(N__20899));
    LocalMux I__4827 (
            .O(N__20921),
            .I(N__20896));
    LocalMux I__4826 (
            .O(N__20914),
            .I(N__20889));
    LocalMux I__4825 (
            .O(N__20907),
            .I(N__20889));
    LocalMux I__4824 (
            .O(N__20902),
            .I(N__20889));
    Span4Mux_v I__4823 (
            .O(N__20899),
            .I(N__20886));
    Span4Mux_h I__4822 (
            .O(N__20896),
            .I(N__20881));
    Span4Mux_v I__4821 (
            .O(N__20889),
            .I(N__20881));
    Span4Mux_h I__4820 (
            .O(N__20886),
            .I(N__20878));
    Odrv4 I__4819 (
            .O(N__20881),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__4818 (
            .O(N__20878),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    CascadeMux I__4817 (
            .O(N__20873),
            .I(N__20870));
    InMux I__4816 (
            .O(N__20870),
            .I(N__20867));
    LocalMux I__4815 (
            .O(N__20867),
            .I(N__20864));
    Span4Mux_h I__4814 (
            .O(N__20864),
            .I(N__20861));
    Span4Mux_h I__4813 (
            .O(N__20861),
            .I(N__20858));
    Odrv4 I__4812 (
            .O(N__20858),
            .I(\delay_measurement_inst.un1_tr_state_1_i_0_0 ));
    InMux I__4811 (
            .O(N__20855),
            .I(N__20849));
    InMux I__4810 (
            .O(N__20854),
            .I(N__20849));
    LocalMux I__4809 (
            .O(N__20849),
            .I(\phase_controller_inst1.T01_0_sqmuxa ));
    CascadeMux I__4808 (
            .O(N__20846),
            .I(N__20834));
    CascadeMux I__4807 (
            .O(N__20845),
            .I(N__20831));
    CascadeMux I__4806 (
            .O(N__20844),
            .I(N__20828));
    CascadeMux I__4805 (
            .O(N__20843),
            .I(N__20821));
    CascadeMux I__4804 (
            .O(N__20842),
            .I(N__20818));
    CascadeMux I__4803 (
            .O(N__20841),
            .I(N__20815));
    CascadeMux I__4802 (
            .O(N__20840),
            .I(N__20805));
    CascadeMux I__4801 (
            .O(N__20839),
            .I(N__20802));
    CascadeMux I__4800 (
            .O(N__20838),
            .I(N__20799));
    CascadeMux I__4799 (
            .O(N__20837),
            .I(N__20796));
    InMux I__4798 (
            .O(N__20834),
            .I(N__20781));
    InMux I__4797 (
            .O(N__20831),
            .I(N__20781));
    InMux I__4796 (
            .O(N__20828),
            .I(N__20781));
    InMux I__4795 (
            .O(N__20827),
            .I(N__20781));
    InMux I__4794 (
            .O(N__20826),
            .I(N__20781));
    InMux I__4793 (
            .O(N__20825),
            .I(N__20781));
    InMux I__4792 (
            .O(N__20824),
            .I(N__20781));
    InMux I__4791 (
            .O(N__20821),
            .I(N__20775));
    InMux I__4790 (
            .O(N__20818),
            .I(N__20766));
    InMux I__4789 (
            .O(N__20815),
            .I(N__20766));
    InMux I__4788 (
            .O(N__20814),
            .I(N__20766));
    InMux I__4787 (
            .O(N__20813),
            .I(N__20766));
    CascadeMux I__4786 (
            .O(N__20812),
            .I(N__20763));
    InMux I__4785 (
            .O(N__20811),
            .I(N__20746));
    InMux I__4784 (
            .O(N__20810),
            .I(N__20746));
    InMux I__4783 (
            .O(N__20809),
            .I(N__20746));
    InMux I__4782 (
            .O(N__20808),
            .I(N__20746));
    InMux I__4781 (
            .O(N__20805),
            .I(N__20746));
    InMux I__4780 (
            .O(N__20802),
            .I(N__20746));
    InMux I__4779 (
            .O(N__20799),
            .I(N__20746));
    InMux I__4778 (
            .O(N__20796),
            .I(N__20746));
    LocalMux I__4777 (
            .O(N__20781),
            .I(N__20743));
    InMux I__4776 (
            .O(N__20780),
            .I(N__20738));
    InMux I__4775 (
            .O(N__20779),
            .I(N__20738));
    CascadeMux I__4774 (
            .O(N__20778),
            .I(N__20735));
    LocalMux I__4773 (
            .O(N__20775),
            .I(N__20730));
    LocalMux I__4772 (
            .O(N__20766),
            .I(N__20730));
    InMux I__4771 (
            .O(N__20763),
            .I(N__20727));
    LocalMux I__4770 (
            .O(N__20746),
            .I(N__20724));
    Span4Mux_h I__4769 (
            .O(N__20743),
            .I(N__20721));
    LocalMux I__4768 (
            .O(N__20738),
            .I(N__20718));
    InMux I__4767 (
            .O(N__20735),
            .I(N__20715));
    Span4Mux_v I__4766 (
            .O(N__20730),
            .I(N__20712));
    LocalMux I__4765 (
            .O(N__20727),
            .I(N__20707));
    Span4Mux_h I__4764 (
            .O(N__20724),
            .I(N__20707));
    Span4Mux_v I__4763 (
            .O(N__20721),
            .I(N__20704));
    Span4Mux_h I__4762 (
            .O(N__20718),
            .I(N__20701));
    LocalMux I__4761 (
            .O(N__20715),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__4760 (
            .O(N__20712),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__4759 (
            .O(N__20707),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__4758 (
            .O(N__20704),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__4757 (
            .O(N__20701),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__4756 (
            .O(N__20690),
            .I(N__20684));
    InMux I__4755 (
            .O(N__20689),
            .I(N__20684));
    LocalMux I__4754 (
            .O(N__20684),
            .I(\phase_controller_inst1.N_83 ));
    InMux I__4753 (
            .O(N__20681),
            .I(N__20674));
    InMux I__4752 (
            .O(N__20680),
            .I(N__20674));
    InMux I__4751 (
            .O(N__20679),
            .I(N__20671));
    LocalMux I__4750 (
            .O(N__20674),
            .I(N__20666));
    LocalMux I__4749 (
            .O(N__20671),
            .I(N__20666));
    Odrv12 I__4748 (
            .O(N__20666),
            .I(il_max_comp1_D2));
    InMux I__4747 (
            .O(N__20663),
            .I(N__20660));
    LocalMux I__4746 (
            .O(N__20660),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    CascadeMux I__4745 (
            .O(N__20657),
            .I(N__20641));
    CascadeMux I__4744 (
            .O(N__20656),
            .I(N__20638));
    CascadeMux I__4743 (
            .O(N__20655),
            .I(N__20635));
    CascadeMux I__4742 (
            .O(N__20654),
            .I(N__20629));
    CascadeMux I__4741 (
            .O(N__20653),
            .I(N__20626));
    CascadeMux I__4740 (
            .O(N__20652),
            .I(N__20623));
    CascadeMux I__4739 (
            .O(N__20651),
            .I(N__20620));
    CascadeMux I__4738 (
            .O(N__20650),
            .I(N__20617));
    CascadeMux I__4737 (
            .O(N__20649),
            .I(N__20612));
    CascadeMux I__4736 (
            .O(N__20648),
            .I(N__20608));
    CascadeMux I__4735 (
            .O(N__20647),
            .I(N__20605));
    CascadeMux I__4734 (
            .O(N__20646),
            .I(N__20602));
    CascadeMux I__4733 (
            .O(N__20645),
            .I(N__20599));
    CascadeMux I__4732 (
            .O(N__20644),
            .I(N__20596));
    InMux I__4731 (
            .O(N__20641),
            .I(N__20581));
    InMux I__4730 (
            .O(N__20638),
            .I(N__20581));
    InMux I__4729 (
            .O(N__20635),
            .I(N__20581));
    InMux I__4728 (
            .O(N__20634),
            .I(N__20581));
    InMux I__4727 (
            .O(N__20633),
            .I(N__20581));
    InMux I__4726 (
            .O(N__20632),
            .I(N__20581));
    InMux I__4725 (
            .O(N__20629),
            .I(N__20572));
    InMux I__4724 (
            .O(N__20626),
            .I(N__20572));
    InMux I__4723 (
            .O(N__20623),
            .I(N__20572));
    InMux I__4722 (
            .O(N__20620),
            .I(N__20572));
    InMux I__4721 (
            .O(N__20617),
            .I(N__20565));
    InMux I__4720 (
            .O(N__20616),
            .I(N__20565));
    InMux I__4719 (
            .O(N__20615),
            .I(N__20565));
    InMux I__4718 (
            .O(N__20612),
            .I(N__20560));
    InMux I__4717 (
            .O(N__20611),
            .I(N__20560));
    InMux I__4716 (
            .O(N__20608),
            .I(N__20551));
    InMux I__4715 (
            .O(N__20605),
            .I(N__20551));
    InMux I__4714 (
            .O(N__20602),
            .I(N__20551));
    InMux I__4713 (
            .O(N__20599),
            .I(N__20551));
    InMux I__4712 (
            .O(N__20596),
            .I(N__20546));
    InMux I__4711 (
            .O(N__20595),
            .I(N__20546));
    CascadeMux I__4710 (
            .O(N__20594),
            .I(N__20542));
    LocalMux I__4709 (
            .O(N__20581),
            .I(N__20539));
    LocalMux I__4708 (
            .O(N__20572),
            .I(N__20534));
    LocalMux I__4707 (
            .O(N__20565),
            .I(N__20534));
    LocalMux I__4706 (
            .O(N__20560),
            .I(N__20527));
    LocalMux I__4705 (
            .O(N__20551),
            .I(N__20527));
    LocalMux I__4704 (
            .O(N__20546),
            .I(N__20527));
    InMux I__4703 (
            .O(N__20545),
            .I(N__20524));
    InMux I__4702 (
            .O(N__20542),
            .I(N__20520));
    Span4Mux_h I__4701 (
            .O(N__20539),
            .I(N__20513));
    Span4Mux_v I__4700 (
            .O(N__20534),
            .I(N__20513));
    Span4Mux_v I__4699 (
            .O(N__20527),
            .I(N__20513));
    LocalMux I__4698 (
            .O(N__20524),
            .I(N__20510));
    InMux I__4697 (
            .O(N__20523),
            .I(N__20507));
    LocalMux I__4696 (
            .O(N__20520),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__4695 (
            .O(N__20513),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__4694 (
            .O(N__20510),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__4693 (
            .O(N__20507),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__4692 (
            .O(N__20498),
            .I(N__20491));
    InMux I__4691 (
            .O(N__20497),
            .I(N__20491));
    InMux I__4690 (
            .O(N__20496),
            .I(N__20488));
    LocalMux I__4689 (
            .O(N__20491),
            .I(N__20484));
    LocalMux I__4688 (
            .O(N__20488),
            .I(N__20481));
    InMux I__4687 (
            .O(N__20487),
            .I(N__20478));
    Span4Mux_h I__4686 (
            .O(N__20484),
            .I(N__20475));
    Span4Mux_h I__4685 (
            .O(N__20481),
            .I(N__20472));
    LocalMux I__4684 (
            .O(N__20478),
            .I(\phase_controller_slave.tr_time_passed ));
    Odrv4 I__4683 (
            .O(N__20475),
            .I(\phase_controller_slave.tr_time_passed ));
    Odrv4 I__4682 (
            .O(N__20472),
            .I(\phase_controller_slave.tr_time_passed ));
    InMux I__4681 (
            .O(N__20465),
            .I(N__20458));
    InMux I__4680 (
            .O(N__20464),
            .I(N__20458));
    InMux I__4679 (
            .O(N__20463),
            .I(N__20455));
    LocalMux I__4678 (
            .O(N__20458),
            .I(\phase_controller_slave.stateZ0Z_0 ));
    LocalMux I__4677 (
            .O(N__20455),
            .I(\phase_controller_slave.stateZ0Z_0 ));
    InMux I__4676 (
            .O(N__20450),
            .I(N__20446));
    InMux I__4675 (
            .O(N__20449),
            .I(N__20443));
    LocalMux I__4674 (
            .O(N__20446),
            .I(shift_flag_start));
    LocalMux I__4673 (
            .O(N__20443),
            .I(shift_flag_start));
    InMux I__4672 (
            .O(N__20438),
            .I(N__20432));
    InMux I__4671 (
            .O(N__20437),
            .I(N__20427));
    InMux I__4670 (
            .O(N__20436),
            .I(N__20427));
    InMux I__4669 (
            .O(N__20435),
            .I(N__20424));
    LocalMux I__4668 (
            .O(N__20432),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__4667 (
            .O(N__20427),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__4666 (
            .O(N__20424),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    InMux I__4665 (
            .O(N__20417),
            .I(N__20411));
    InMux I__4664 (
            .O(N__20416),
            .I(N__20411));
    LocalMux I__4663 (
            .O(N__20411),
            .I(N__20407));
    InMux I__4662 (
            .O(N__20410),
            .I(N__20404));
    Span4Mux_h I__4661 (
            .O(N__20407),
            .I(N__20400));
    LocalMux I__4660 (
            .O(N__20404),
            .I(N__20397));
    InMux I__4659 (
            .O(N__20403),
            .I(N__20394));
    Sp12to4 I__4658 (
            .O(N__20400),
            .I(N__20391));
    Span4Mux_h I__4657 (
            .O(N__20397),
            .I(N__20388));
    LocalMux I__4656 (
            .O(N__20394),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv12 I__4655 (
            .O(N__20391),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__4654 (
            .O(N__20388),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__4653 (
            .O(N__20381),
            .I(N__20378));
    LocalMux I__4652 (
            .O(N__20378),
            .I(\phase_controller_inst1.N_88 ));
    InMux I__4651 (
            .O(N__20375),
            .I(N__20369));
    InMux I__4650 (
            .O(N__20374),
            .I(N__20369));
    LocalMux I__4649 (
            .O(N__20369),
            .I(N__20366));
    Span4Mux_h I__4648 (
            .O(N__20366),
            .I(N__20362));
    InMux I__4647 (
            .O(N__20365),
            .I(N__20359));
    Sp12to4 I__4646 (
            .O(N__20362),
            .I(N__20354));
    LocalMux I__4645 (
            .O(N__20359),
            .I(N__20354));
    Span12Mux_v I__4644 (
            .O(N__20354),
            .I(N__20351));
    Odrv12 I__4643 (
            .O(N__20351),
            .I(il_max_comp2_D2));
    CascadeMux I__4642 (
            .O(N__20348),
            .I(N__20345));
    InMux I__4641 (
            .O(N__20345),
            .I(N__20340));
    CascadeMux I__4640 (
            .O(N__20344),
            .I(N__20337));
    CascadeMux I__4639 (
            .O(N__20343),
            .I(N__20334));
    LocalMux I__4638 (
            .O(N__20340),
            .I(N__20330));
    InMux I__4637 (
            .O(N__20337),
            .I(N__20327));
    InMux I__4636 (
            .O(N__20334),
            .I(N__20324));
    CascadeMux I__4635 (
            .O(N__20333),
            .I(N__20321));
    Span4Mux_h I__4634 (
            .O(N__20330),
            .I(N__20318));
    LocalMux I__4633 (
            .O(N__20327),
            .I(N__20315));
    LocalMux I__4632 (
            .O(N__20324),
            .I(N__20312));
    InMux I__4631 (
            .O(N__20321),
            .I(N__20309));
    Odrv4 I__4630 (
            .O(N__20318),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    Odrv4 I__4629 (
            .O(N__20315),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    Odrv4 I__4628 (
            .O(N__20312),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    LocalMux I__4627 (
            .O(N__20309),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    InMux I__4626 (
            .O(N__20300),
            .I(N__20296));
    InMux I__4625 (
            .O(N__20299),
            .I(N__20293));
    LocalMux I__4624 (
            .O(N__20296),
            .I(\phase_controller_slave.un1_startZ0 ));
    LocalMux I__4623 (
            .O(N__20293),
            .I(\phase_controller_slave.un1_startZ0 ));
    InMux I__4622 (
            .O(N__20288),
            .I(N__20282));
    InMux I__4621 (
            .O(N__20287),
            .I(N__20277));
    InMux I__4620 (
            .O(N__20286),
            .I(N__20277));
    InMux I__4619 (
            .O(N__20285),
            .I(N__20274));
    LocalMux I__4618 (
            .O(N__20282),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    LocalMux I__4617 (
            .O(N__20277),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    LocalMux I__4616 (
            .O(N__20274),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    CascadeMux I__4615 (
            .O(N__20267),
            .I(N__20263));
    InMux I__4614 (
            .O(N__20266),
            .I(N__20257));
    InMux I__4613 (
            .O(N__20263),
            .I(N__20257));
    InMux I__4612 (
            .O(N__20262),
            .I(N__20254));
    LocalMux I__4611 (
            .O(N__20257),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__4610 (
            .O(N__20254),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__4609 (
            .O(N__20249),
            .I(N__20245));
    InMux I__4608 (
            .O(N__20248),
            .I(N__20242));
    LocalMux I__4607 (
            .O(N__20245),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__4606 (
            .O(N__20242),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__4605 (
            .O(N__20237),
            .I(N__20234));
    LocalMux I__4604 (
            .O(N__20234),
            .I(\phase_controller_slave.start_timer_tr_0_sqmuxa ));
    InMux I__4603 (
            .O(N__20231),
            .I(N__20228));
    LocalMux I__4602 (
            .O(N__20228),
            .I(N__20225));
    Span4Mux_v I__4601 (
            .O(N__20225),
            .I(N__20222));
    Span4Mux_v I__4600 (
            .O(N__20222),
            .I(N__20219));
    Odrv4 I__4599 (
            .O(N__20219),
            .I(il_min_comp2_D1));
    InMux I__4598 (
            .O(N__20216),
            .I(N__20213));
    LocalMux I__4597 (
            .O(N__20213),
            .I(\phase_controller_slave.N_20 ));
    InMux I__4596 (
            .O(N__20210),
            .I(N__20205));
    InMux I__4595 (
            .O(N__20209),
            .I(N__20202));
    InMux I__4594 (
            .O(N__20208),
            .I(N__20199));
    LocalMux I__4593 (
            .O(N__20205),
            .I(N__20196));
    LocalMux I__4592 (
            .O(N__20202),
            .I(N__20191));
    LocalMux I__4591 (
            .O(N__20199),
            .I(N__20191));
    Odrv12 I__4590 (
            .O(N__20196),
            .I(il_min_comp1_D2));
    Odrv4 I__4589 (
            .O(N__20191),
            .I(il_min_comp1_D2));
    InMux I__4588 (
            .O(N__20186),
            .I(N__20183));
    LocalMux I__4587 (
            .O(N__20183),
            .I(N__20180));
    Span4Mux_h I__4586 (
            .O(N__20180),
            .I(N__20177));
    Span4Mux_v I__4585 (
            .O(N__20177),
            .I(N__20174));
    Span4Mux_v I__4584 (
            .O(N__20174),
            .I(N__20171));
    Odrv4 I__4583 (
            .O(N__20171),
            .I(il_max_comp1_c));
    InMux I__4582 (
            .O(N__20168),
            .I(N__20165));
    LocalMux I__4581 (
            .O(N__20165),
            .I(il_max_comp1_D1));
    InMux I__4580 (
            .O(N__20162),
            .I(N__20159));
    LocalMux I__4579 (
            .O(N__20159),
            .I(N__20156));
    Span4Mux_v I__4578 (
            .O(N__20156),
            .I(N__20153));
    Sp12to4 I__4577 (
            .O(N__20153),
            .I(N__20150));
    Span12Mux_h I__4576 (
            .O(N__20150),
            .I(N__20147));
    Odrv12 I__4575 (
            .O(N__20147),
            .I(il_min_comp1_c));
    InMux I__4574 (
            .O(N__20144),
            .I(N__20141));
    LocalMux I__4573 (
            .O(N__20141),
            .I(il_min_comp1_D1));
    InMux I__4572 (
            .O(N__20138),
            .I(N__20132));
    InMux I__4571 (
            .O(N__20137),
            .I(N__20121));
    InMux I__4570 (
            .O(N__20136),
            .I(N__20121));
    InMux I__4569 (
            .O(N__20135),
            .I(N__20121));
    LocalMux I__4568 (
            .O(N__20132),
            .I(N__20113));
    CascadeMux I__4567 (
            .O(N__20131),
            .I(N__20110));
    InMux I__4566 (
            .O(N__20130),
            .I(N__20104));
    InMux I__4565 (
            .O(N__20129),
            .I(N__20104));
    InMux I__4564 (
            .O(N__20128),
            .I(N__20101));
    LocalMux I__4563 (
            .O(N__20121),
            .I(N__20098));
    InMux I__4562 (
            .O(N__20120),
            .I(N__20089));
    InMux I__4561 (
            .O(N__20119),
            .I(N__20089));
    InMux I__4560 (
            .O(N__20118),
            .I(N__20089));
    InMux I__4559 (
            .O(N__20117),
            .I(N__20089));
    InMux I__4558 (
            .O(N__20116),
            .I(N__20086));
    Span4Mux_h I__4557 (
            .O(N__20113),
            .I(N__20083));
    InMux I__4556 (
            .O(N__20110),
            .I(N__20078));
    InMux I__4555 (
            .O(N__20109),
            .I(N__20078));
    LocalMux I__4554 (
            .O(N__20104),
            .I(N__20075));
    LocalMux I__4553 (
            .O(N__20101),
            .I(N__20072));
    Span4Mux_v I__4552 (
            .O(N__20098),
            .I(N__20067));
    LocalMux I__4551 (
            .O(N__20089),
            .I(N__20062));
    LocalMux I__4550 (
            .O(N__20086),
            .I(N__20062));
    Span4Mux_h I__4549 (
            .O(N__20083),
            .I(N__20059));
    LocalMux I__4548 (
            .O(N__20078),
            .I(N__20052));
    Span4Mux_h I__4547 (
            .O(N__20075),
            .I(N__20052));
    Span4Mux_h I__4546 (
            .O(N__20072),
            .I(N__20052));
    InMux I__4545 (
            .O(N__20071),
            .I(N__20049));
    InMux I__4544 (
            .O(N__20070),
            .I(N__20046));
    Odrv4 I__4543 (
            .O(N__20067),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    Odrv4 I__4542 (
            .O(N__20062),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    Odrv4 I__4541 (
            .O(N__20059),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    Odrv4 I__4540 (
            .O(N__20052),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    LocalMux I__4539 (
            .O(N__20049),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    LocalMux I__4538 (
            .O(N__20046),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    InMux I__4537 (
            .O(N__20033),
            .I(N__20028));
    InMux I__4536 (
            .O(N__20032),
            .I(N__20021));
    InMux I__4535 (
            .O(N__20031),
            .I(N__20021));
    LocalMux I__4534 (
            .O(N__20028),
            .I(N__20015));
    CascadeMux I__4533 (
            .O(N__20027),
            .I(N__20011));
    CascadeMux I__4532 (
            .O(N__20026),
            .I(N__20008));
    LocalMux I__4531 (
            .O(N__20021),
            .I(N__20005));
    InMux I__4530 (
            .O(N__20020),
            .I(N__20002));
    InMux I__4529 (
            .O(N__20019),
            .I(N__19997));
    InMux I__4528 (
            .O(N__20018),
            .I(N__19997));
    Span4Mux_v I__4527 (
            .O(N__20015),
            .I(N__19993));
    InMux I__4526 (
            .O(N__20014),
            .I(N__19986));
    InMux I__4525 (
            .O(N__20011),
            .I(N__19986));
    InMux I__4524 (
            .O(N__20008),
            .I(N__19986));
    Span4Mux_h I__4523 (
            .O(N__20005),
            .I(N__19983));
    LocalMux I__4522 (
            .O(N__20002),
            .I(N__19978));
    LocalMux I__4521 (
            .O(N__19997),
            .I(N__19978));
    InMux I__4520 (
            .O(N__19996),
            .I(N__19975));
    Sp12to4 I__4519 (
            .O(N__19993),
            .I(N__19970));
    LocalMux I__4518 (
            .O(N__19986),
            .I(N__19970));
    Odrv4 I__4517 (
            .O(N__19983),
            .I(measured_delay_tr_15));
    Odrv4 I__4516 (
            .O(N__19978),
            .I(measured_delay_tr_15));
    LocalMux I__4515 (
            .O(N__19975),
            .I(measured_delay_tr_15));
    Odrv12 I__4514 (
            .O(N__19970),
            .I(measured_delay_tr_15));
    InMux I__4513 (
            .O(N__19961),
            .I(N__19958));
    LocalMux I__4512 (
            .O(N__19958),
            .I(N__19955));
    Span4Mux_h I__4511 (
            .O(N__19955),
            .I(N__19952));
    Odrv4 I__4510 (
            .O(N__19952),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    CEMux I__4509 (
            .O(N__19949),
            .I(N__19946));
    LocalMux I__4508 (
            .O(N__19946),
            .I(N__19941));
    CEMux I__4507 (
            .O(N__19945),
            .I(N__19938));
    CEMux I__4506 (
            .O(N__19944),
            .I(N__19935));
    Span4Mux_v I__4505 (
            .O(N__19941),
            .I(N__19930));
    LocalMux I__4504 (
            .O(N__19938),
            .I(N__19930));
    LocalMux I__4503 (
            .O(N__19935),
            .I(N__19926));
    Span4Mux_h I__4502 (
            .O(N__19930),
            .I(N__19923));
    CEMux I__4501 (
            .O(N__19929),
            .I(N__19920));
    Span4Mux_h I__4500 (
            .O(N__19926),
            .I(N__19917));
    Span4Mux_h I__4499 (
            .O(N__19923),
            .I(N__19914));
    LocalMux I__4498 (
            .O(N__19920),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__4497 (
            .O(N__19917),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__4496 (
            .O(N__19914),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    CascadeMux I__4495 (
            .O(N__19907),
            .I(N__19895));
    CascadeMux I__4494 (
            .O(N__19906),
            .I(N__19888));
    CascadeMux I__4493 (
            .O(N__19905),
            .I(N__19885));
    CascadeMux I__4492 (
            .O(N__19904),
            .I(N__19882));
    CascadeMux I__4491 (
            .O(N__19903),
            .I(N__19879));
    CascadeMux I__4490 (
            .O(N__19902),
            .I(N__19874));
    CascadeMux I__4489 (
            .O(N__19901),
            .I(N__19870));
    CascadeMux I__4488 (
            .O(N__19900),
            .I(N__19867));
    CascadeMux I__4487 (
            .O(N__19899),
            .I(N__19864));
    CascadeMux I__4486 (
            .O(N__19898),
            .I(N__19861));
    InMux I__4485 (
            .O(N__19895),
            .I(N__19854));
    InMux I__4484 (
            .O(N__19894),
            .I(N__19837));
    InMux I__4483 (
            .O(N__19893),
            .I(N__19837));
    InMux I__4482 (
            .O(N__19892),
            .I(N__19837));
    InMux I__4481 (
            .O(N__19891),
            .I(N__19837));
    InMux I__4480 (
            .O(N__19888),
            .I(N__19837));
    InMux I__4479 (
            .O(N__19885),
            .I(N__19837));
    InMux I__4478 (
            .O(N__19882),
            .I(N__19837));
    InMux I__4477 (
            .O(N__19879),
            .I(N__19837));
    InMux I__4476 (
            .O(N__19878),
            .I(N__19830));
    InMux I__4475 (
            .O(N__19877),
            .I(N__19830));
    InMux I__4474 (
            .O(N__19874),
            .I(N__19830));
    CascadeMux I__4473 (
            .O(N__19873),
            .I(N__19827));
    InMux I__4472 (
            .O(N__19870),
            .I(N__19810));
    InMux I__4471 (
            .O(N__19867),
            .I(N__19810));
    InMux I__4470 (
            .O(N__19864),
            .I(N__19810));
    InMux I__4469 (
            .O(N__19861),
            .I(N__19810));
    InMux I__4468 (
            .O(N__19860),
            .I(N__19810));
    InMux I__4467 (
            .O(N__19859),
            .I(N__19810));
    InMux I__4466 (
            .O(N__19858),
            .I(N__19810));
    InMux I__4465 (
            .O(N__19857),
            .I(N__19810));
    LocalMux I__4464 (
            .O(N__19854),
            .I(N__19807));
    LocalMux I__4463 (
            .O(N__19837),
            .I(N__19802));
    LocalMux I__4462 (
            .O(N__19830),
            .I(N__19802));
    InMux I__4461 (
            .O(N__19827),
            .I(N__19799));
    LocalMux I__4460 (
            .O(N__19810),
            .I(N__19794));
    Span4Mux_v I__4459 (
            .O(N__19807),
            .I(N__19794));
    Span4Mux_v I__4458 (
            .O(N__19802),
            .I(N__19791));
    LocalMux I__4457 (
            .O(N__19799),
            .I(N__19785));
    Sp12to4 I__4456 (
            .O(N__19794),
            .I(N__19782));
    Span4Mux_h I__4455 (
            .O(N__19791),
            .I(N__19779));
    InMux I__4454 (
            .O(N__19790),
            .I(N__19776));
    InMux I__4453 (
            .O(N__19789),
            .I(N__19773));
    InMux I__4452 (
            .O(N__19788),
            .I(N__19770));
    Span4Mux_h I__4451 (
            .O(N__19785),
            .I(N__19767));
    Span12Mux_s5_h I__4450 (
            .O(N__19782),
            .I(N__19758));
    Sp12to4 I__4449 (
            .O(N__19779),
            .I(N__19758));
    LocalMux I__4448 (
            .O(N__19776),
            .I(N__19758));
    LocalMux I__4447 (
            .O(N__19773),
            .I(N__19758));
    LocalMux I__4446 (
            .O(N__19770),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__4445 (
            .O(N__19767),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv12 I__4444 (
            .O(N__19758),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    InMux I__4443 (
            .O(N__19751),
            .I(N__19748));
    LocalMux I__4442 (
            .O(N__19748),
            .I(N__19745));
    Odrv4 I__4441 (
            .O(N__19745),
            .I(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ));
    CascadeMux I__4440 (
            .O(N__19742),
            .I(N__19739));
    InMux I__4439 (
            .O(N__19739),
            .I(N__19736));
    LocalMux I__4438 (
            .O(N__19736),
            .I(N__19731));
    InMux I__4437 (
            .O(N__19735),
            .I(N__19728));
    InMux I__4436 (
            .O(N__19734),
            .I(N__19725));
    Odrv12 I__4435 (
            .O(N__19731),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    LocalMux I__4434 (
            .O(N__19728),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    LocalMux I__4433 (
            .O(N__19725),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    InMux I__4432 (
            .O(N__19718),
            .I(N__19715));
    LocalMux I__4431 (
            .O(N__19715),
            .I(N__19710));
    InMux I__4430 (
            .O(N__19714),
            .I(N__19707));
    InMux I__4429 (
            .O(N__19713),
            .I(N__19702));
    Span4Mux_h I__4428 (
            .O(N__19710),
            .I(N__19697));
    LocalMux I__4427 (
            .O(N__19707),
            .I(N__19697));
    InMux I__4426 (
            .O(N__19706),
            .I(N__19692));
    InMux I__4425 (
            .O(N__19705),
            .I(N__19692));
    LocalMux I__4424 (
            .O(N__19702),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__4423 (
            .O(N__19697),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__4422 (
            .O(N__19692),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__4421 (
            .O(N__19685),
            .I(N__19680));
    CascadeMux I__4420 (
            .O(N__19684),
            .I(N__19677));
    InMux I__4419 (
            .O(N__19683),
            .I(N__19674));
    InMux I__4418 (
            .O(N__19680),
            .I(N__19669));
    InMux I__4417 (
            .O(N__19677),
            .I(N__19669));
    LocalMux I__4416 (
            .O(N__19674),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__4415 (
            .O(N__19669),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__4414 (
            .O(N__19664),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    CascadeMux I__4413 (
            .O(N__19661),
            .I(N__19656));
    CascadeMux I__4412 (
            .O(N__19660),
            .I(N__19653));
    InMux I__4411 (
            .O(N__19659),
            .I(N__19650));
    InMux I__4410 (
            .O(N__19656),
            .I(N__19645));
    InMux I__4409 (
            .O(N__19653),
            .I(N__19645));
    LocalMux I__4408 (
            .O(N__19650),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__4407 (
            .O(N__19645),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__4406 (
            .O(N__19640),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__4405 (
            .O(N__19637),
            .I(N__19632));
    InMux I__4404 (
            .O(N__19636),
            .I(N__19629));
    InMux I__4403 (
            .O(N__19635),
            .I(N__19626));
    LocalMux I__4402 (
            .O(N__19632),
            .I(N__19623));
    LocalMux I__4401 (
            .O(N__19629),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__4400 (
            .O(N__19626),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__4399 (
            .O(N__19623),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__4398 (
            .O(N__19616),
            .I(bfn_9_29_0_));
    InMux I__4397 (
            .O(N__19613),
            .I(N__19608));
    InMux I__4396 (
            .O(N__19612),
            .I(N__19605));
    InMux I__4395 (
            .O(N__19611),
            .I(N__19602));
    LocalMux I__4394 (
            .O(N__19608),
            .I(N__19599));
    LocalMux I__4393 (
            .O(N__19605),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__4392 (
            .O(N__19602),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__4391 (
            .O(N__19599),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__4390 (
            .O(N__19592),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    CascadeMux I__4389 (
            .O(N__19589),
            .I(N__19584));
    CascadeMux I__4388 (
            .O(N__19588),
            .I(N__19581));
    InMux I__4387 (
            .O(N__19587),
            .I(N__19578));
    InMux I__4386 (
            .O(N__19584),
            .I(N__19573));
    InMux I__4385 (
            .O(N__19581),
            .I(N__19573));
    LocalMux I__4384 (
            .O(N__19578),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__4383 (
            .O(N__19573),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__4382 (
            .O(N__19568),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    CascadeMux I__4381 (
            .O(N__19565),
            .I(N__19560));
    CascadeMux I__4380 (
            .O(N__19564),
            .I(N__19557));
    InMux I__4379 (
            .O(N__19563),
            .I(N__19554));
    InMux I__4378 (
            .O(N__19560),
            .I(N__19549));
    InMux I__4377 (
            .O(N__19557),
            .I(N__19549));
    LocalMux I__4376 (
            .O(N__19554),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__4375 (
            .O(N__19549),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__4374 (
            .O(N__19544),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__4373 (
            .O(N__19541),
            .I(N__19537));
    InMux I__4372 (
            .O(N__19540),
            .I(N__19534));
    LocalMux I__4371 (
            .O(N__19537),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    LocalMux I__4370 (
            .O(N__19534),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__4369 (
            .O(N__19529),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__4368 (
            .O(N__19526),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__4367 (
            .O(N__19523),
            .I(N__19519));
    InMux I__4366 (
            .O(N__19522),
            .I(N__19516));
    LocalMux I__4365 (
            .O(N__19519),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    LocalMux I__4364 (
            .O(N__19516),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    IoInMux I__4363 (
            .O(N__19511),
            .I(N__19508));
    LocalMux I__4362 (
            .O(N__19508),
            .I(N__19505));
    Span12Mux_s6_v I__4361 (
            .O(N__19505),
            .I(N__19502));
    Span12Mux_v I__4360 (
            .O(N__19502),
            .I(N__19499));
    Odrv12 I__4359 (
            .O(N__19499),
            .I(\delay_measurement_inst.delay_tr_timer.N_138_i ));
    CascadeMux I__4358 (
            .O(N__19496),
            .I(N__19491));
    CascadeMux I__4357 (
            .O(N__19495),
            .I(N__19488));
    InMux I__4356 (
            .O(N__19494),
            .I(N__19485));
    InMux I__4355 (
            .O(N__19491),
            .I(N__19480));
    InMux I__4354 (
            .O(N__19488),
            .I(N__19480));
    LocalMux I__4353 (
            .O(N__19485),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__4352 (
            .O(N__19480),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__4351 (
            .O(N__19475),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    CascadeMux I__4350 (
            .O(N__19472),
            .I(N__19467));
    CascadeMux I__4349 (
            .O(N__19471),
            .I(N__19464));
    InMux I__4348 (
            .O(N__19470),
            .I(N__19461));
    InMux I__4347 (
            .O(N__19467),
            .I(N__19456));
    InMux I__4346 (
            .O(N__19464),
            .I(N__19456));
    LocalMux I__4345 (
            .O(N__19461),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__4344 (
            .O(N__19456),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__4343 (
            .O(N__19451),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__4342 (
            .O(N__19448),
            .I(N__19443));
    InMux I__4341 (
            .O(N__19447),
            .I(N__19440));
    InMux I__4340 (
            .O(N__19446),
            .I(N__19437));
    LocalMux I__4339 (
            .O(N__19443),
            .I(N__19434));
    LocalMux I__4338 (
            .O(N__19440),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__4337 (
            .O(N__19437),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__4336 (
            .O(N__19434),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__4335 (
            .O(N__19427),
            .I(bfn_9_28_0_));
    InMux I__4334 (
            .O(N__19424),
            .I(N__19419));
    InMux I__4333 (
            .O(N__19423),
            .I(N__19416));
    InMux I__4332 (
            .O(N__19422),
            .I(N__19413));
    LocalMux I__4331 (
            .O(N__19419),
            .I(N__19410));
    LocalMux I__4330 (
            .O(N__19416),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__4329 (
            .O(N__19413),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__4328 (
            .O(N__19410),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__4327 (
            .O(N__19403),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    CascadeMux I__4326 (
            .O(N__19400),
            .I(N__19395));
    CascadeMux I__4325 (
            .O(N__19399),
            .I(N__19392));
    InMux I__4324 (
            .O(N__19398),
            .I(N__19389));
    InMux I__4323 (
            .O(N__19395),
            .I(N__19384));
    InMux I__4322 (
            .O(N__19392),
            .I(N__19384));
    LocalMux I__4321 (
            .O(N__19389),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__4320 (
            .O(N__19384),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__4319 (
            .O(N__19379),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    CascadeMux I__4318 (
            .O(N__19376),
            .I(N__19371));
    CascadeMux I__4317 (
            .O(N__19375),
            .I(N__19368));
    InMux I__4316 (
            .O(N__19374),
            .I(N__19365));
    InMux I__4315 (
            .O(N__19371),
            .I(N__19360));
    InMux I__4314 (
            .O(N__19368),
            .I(N__19360));
    LocalMux I__4313 (
            .O(N__19365),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__4312 (
            .O(N__19360),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__4311 (
            .O(N__19355),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__4310 (
            .O(N__19352),
            .I(N__19347));
    InMux I__4309 (
            .O(N__19351),
            .I(N__19342));
    InMux I__4308 (
            .O(N__19350),
            .I(N__19342));
    LocalMux I__4307 (
            .O(N__19347),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__4306 (
            .O(N__19342),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__4305 (
            .O(N__19337),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__4304 (
            .O(N__19334),
            .I(N__19329));
    InMux I__4303 (
            .O(N__19333),
            .I(N__19324));
    InMux I__4302 (
            .O(N__19332),
            .I(N__19324));
    LocalMux I__4301 (
            .O(N__19329),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__4300 (
            .O(N__19324),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__4299 (
            .O(N__19319),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__4298 (
            .O(N__19316),
            .I(N__19311));
    InMux I__4297 (
            .O(N__19315),
            .I(N__19306));
    InMux I__4296 (
            .O(N__19314),
            .I(N__19306));
    LocalMux I__4295 (
            .O(N__19311),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__4294 (
            .O(N__19306),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__4293 (
            .O(N__19301),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    CascadeMux I__4292 (
            .O(N__19298),
            .I(N__19293));
    CascadeMux I__4291 (
            .O(N__19297),
            .I(N__19290));
    InMux I__4290 (
            .O(N__19296),
            .I(N__19287));
    InMux I__4289 (
            .O(N__19293),
            .I(N__19282));
    InMux I__4288 (
            .O(N__19290),
            .I(N__19282));
    LocalMux I__4287 (
            .O(N__19287),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__4286 (
            .O(N__19282),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__4285 (
            .O(N__19277),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    CascadeMux I__4284 (
            .O(N__19274),
            .I(N__19269));
    CascadeMux I__4283 (
            .O(N__19273),
            .I(N__19266));
    InMux I__4282 (
            .O(N__19272),
            .I(N__19263));
    InMux I__4281 (
            .O(N__19269),
            .I(N__19258));
    InMux I__4280 (
            .O(N__19266),
            .I(N__19258));
    LocalMux I__4279 (
            .O(N__19263),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__4278 (
            .O(N__19258),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__4277 (
            .O(N__19253),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__4276 (
            .O(N__19250),
            .I(N__19245));
    InMux I__4275 (
            .O(N__19249),
            .I(N__19242));
    InMux I__4274 (
            .O(N__19248),
            .I(N__19239));
    LocalMux I__4273 (
            .O(N__19245),
            .I(N__19236));
    LocalMux I__4272 (
            .O(N__19242),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__4271 (
            .O(N__19239),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__4270 (
            .O(N__19236),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__4269 (
            .O(N__19229),
            .I(bfn_9_27_0_));
    InMux I__4268 (
            .O(N__19226),
            .I(N__19221));
    InMux I__4267 (
            .O(N__19225),
            .I(N__19218));
    InMux I__4266 (
            .O(N__19224),
            .I(N__19215));
    LocalMux I__4265 (
            .O(N__19221),
            .I(N__19212));
    LocalMux I__4264 (
            .O(N__19218),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__4263 (
            .O(N__19215),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__4262 (
            .O(N__19212),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__4261 (
            .O(N__19205),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    CascadeMux I__4260 (
            .O(N__19202),
            .I(N__19197));
    CascadeMux I__4259 (
            .O(N__19201),
            .I(N__19194));
    InMux I__4258 (
            .O(N__19200),
            .I(N__19191));
    InMux I__4257 (
            .O(N__19197),
            .I(N__19186));
    InMux I__4256 (
            .O(N__19194),
            .I(N__19186));
    LocalMux I__4255 (
            .O(N__19191),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__4254 (
            .O(N__19186),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__4253 (
            .O(N__19181),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    CascadeMux I__4252 (
            .O(N__19178),
            .I(N__19173));
    CascadeMux I__4251 (
            .O(N__19177),
            .I(N__19170));
    InMux I__4250 (
            .O(N__19176),
            .I(N__19167));
    InMux I__4249 (
            .O(N__19173),
            .I(N__19162));
    InMux I__4248 (
            .O(N__19170),
            .I(N__19162));
    LocalMux I__4247 (
            .O(N__19167),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__4246 (
            .O(N__19162),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__4245 (
            .O(N__19157),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__4244 (
            .O(N__19154),
            .I(N__19149));
    InMux I__4243 (
            .O(N__19153),
            .I(N__19144));
    InMux I__4242 (
            .O(N__19152),
            .I(N__19144));
    LocalMux I__4241 (
            .O(N__19149),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__4240 (
            .O(N__19144),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__4239 (
            .O(N__19139),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__4238 (
            .O(N__19136),
            .I(N__19131));
    InMux I__4237 (
            .O(N__19135),
            .I(N__19126));
    InMux I__4236 (
            .O(N__19134),
            .I(N__19126));
    LocalMux I__4235 (
            .O(N__19131),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__4234 (
            .O(N__19126),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__4233 (
            .O(N__19121),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    CascadeMux I__4232 (
            .O(N__19118),
            .I(N__19089));
    CascadeMux I__4231 (
            .O(N__19117),
            .I(N__19085));
    CascadeMux I__4230 (
            .O(N__19116),
            .I(N__19082));
    CascadeMux I__4229 (
            .O(N__19115),
            .I(N__19078));
    CascadeMux I__4228 (
            .O(N__19114),
            .I(N__19074));
    InMux I__4227 (
            .O(N__19113),
            .I(N__19055));
    InMux I__4226 (
            .O(N__19112),
            .I(N__19055));
    InMux I__4225 (
            .O(N__19111),
            .I(N__19055));
    InMux I__4224 (
            .O(N__19110),
            .I(N__19055));
    InMux I__4223 (
            .O(N__19109),
            .I(N__19055));
    InMux I__4222 (
            .O(N__19108),
            .I(N__19055));
    InMux I__4221 (
            .O(N__19107),
            .I(N__19055));
    InMux I__4220 (
            .O(N__19106),
            .I(N__19055));
    InMux I__4219 (
            .O(N__19105),
            .I(N__19038));
    InMux I__4218 (
            .O(N__19104),
            .I(N__19038));
    InMux I__4217 (
            .O(N__19103),
            .I(N__19038));
    InMux I__4216 (
            .O(N__19102),
            .I(N__19038));
    InMux I__4215 (
            .O(N__19101),
            .I(N__19038));
    InMux I__4214 (
            .O(N__19100),
            .I(N__19038));
    InMux I__4213 (
            .O(N__19099),
            .I(N__19038));
    InMux I__4212 (
            .O(N__19098),
            .I(N__19038));
    InMux I__4211 (
            .O(N__19097),
            .I(N__19021));
    InMux I__4210 (
            .O(N__19096),
            .I(N__19021));
    InMux I__4209 (
            .O(N__19095),
            .I(N__19021));
    InMux I__4208 (
            .O(N__19094),
            .I(N__19021));
    InMux I__4207 (
            .O(N__19093),
            .I(N__19021));
    InMux I__4206 (
            .O(N__19092),
            .I(N__19021));
    InMux I__4205 (
            .O(N__19089),
            .I(N__19021));
    InMux I__4204 (
            .O(N__19088),
            .I(N__19021));
    InMux I__4203 (
            .O(N__19085),
            .I(N__19004));
    InMux I__4202 (
            .O(N__19082),
            .I(N__19004));
    InMux I__4201 (
            .O(N__19081),
            .I(N__19004));
    InMux I__4200 (
            .O(N__19078),
            .I(N__19004));
    InMux I__4199 (
            .O(N__19077),
            .I(N__19004));
    InMux I__4198 (
            .O(N__19074),
            .I(N__19004));
    InMux I__4197 (
            .O(N__19073),
            .I(N__19004));
    InMux I__4196 (
            .O(N__19072),
            .I(N__19004));
    LocalMux I__4195 (
            .O(N__19055),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    LocalMux I__4194 (
            .O(N__19038),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    LocalMux I__4193 (
            .O(N__19021),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    LocalMux I__4192 (
            .O(N__19004),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    InMux I__4191 (
            .O(N__18995),
            .I(N__18965));
    InMux I__4190 (
            .O(N__18994),
            .I(N__18965));
    InMux I__4189 (
            .O(N__18993),
            .I(N__18965));
    InMux I__4188 (
            .O(N__18992),
            .I(N__18965));
    InMux I__4187 (
            .O(N__18991),
            .I(N__18965));
    InMux I__4186 (
            .O(N__18990),
            .I(N__18965));
    InMux I__4185 (
            .O(N__18989),
            .I(N__18954));
    InMux I__4184 (
            .O(N__18988),
            .I(N__18954));
    InMux I__4183 (
            .O(N__18987),
            .I(N__18954));
    InMux I__4182 (
            .O(N__18986),
            .I(N__18954));
    InMux I__4181 (
            .O(N__18985),
            .I(N__18954));
    InMux I__4180 (
            .O(N__18984),
            .I(N__18949));
    InMux I__4179 (
            .O(N__18983),
            .I(N__18949));
    InMux I__4178 (
            .O(N__18982),
            .I(N__18938));
    InMux I__4177 (
            .O(N__18981),
            .I(N__18938));
    InMux I__4176 (
            .O(N__18980),
            .I(N__18938));
    InMux I__4175 (
            .O(N__18979),
            .I(N__18938));
    InMux I__4174 (
            .O(N__18978),
            .I(N__18938));
    LocalMux I__4173 (
            .O(N__18965),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    LocalMux I__4172 (
            .O(N__18954),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    LocalMux I__4171 (
            .O(N__18949),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    LocalMux I__4170 (
            .O(N__18938),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    CascadeMux I__4169 (
            .O(N__18929),
            .I(N__18925));
    InMux I__4168 (
            .O(N__18928),
            .I(N__18922));
    InMux I__4167 (
            .O(N__18925),
            .I(N__18919));
    LocalMux I__4166 (
            .O(N__18922),
            .I(measured_delay_hc_26));
    LocalMux I__4165 (
            .O(N__18919),
            .I(measured_delay_hc_26));
    InMux I__4164 (
            .O(N__18914),
            .I(N__18911));
    LocalMux I__4163 (
            .O(N__18911),
            .I(N__18908));
    Span4Mux_v I__4162 (
            .O(N__18908),
            .I(N__18904));
    InMux I__4161 (
            .O(N__18907),
            .I(N__18901));
    Odrv4 I__4160 (
            .O(N__18904),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    LocalMux I__4159 (
            .O(N__18901),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    CascadeMux I__4158 (
            .O(N__18896),
            .I(N__18893));
    InMux I__4157 (
            .O(N__18893),
            .I(N__18889));
    CascadeMux I__4156 (
            .O(N__18892),
            .I(N__18885));
    LocalMux I__4155 (
            .O(N__18889),
            .I(N__18882));
    InMux I__4154 (
            .O(N__18888),
            .I(N__18879));
    InMux I__4153 (
            .O(N__18885),
            .I(N__18876));
    Odrv4 I__4152 (
            .O(N__18882),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    LocalMux I__4151 (
            .O(N__18879),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    LocalMux I__4150 (
            .O(N__18876),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    CEMux I__4149 (
            .O(N__18869),
            .I(N__18854));
    CEMux I__4148 (
            .O(N__18868),
            .I(N__18854));
    CEMux I__4147 (
            .O(N__18867),
            .I(N__18854));
    CEMux I__4146 (
            .O(N__18866),
            .I(N__18854));
    CEMux I__4145 (
            .O(N__18865),
            .I(N__18854));
    GlobalMux I__4144 (
            .O(N__18854),
            .I(N__18851));
    gio2CtrlBuf I__4143 (
            .O(N__18851),
            .I(\delay_measurement_inst.delay_hc_timer.N_136_i_g ));
    InMux I__4142 (
            .O(N__18848),
            .I(N__18843));
    InMux I__4141 (
            .O(N__18847),
            .I(N__18840));
    InMux I__4140 (
            .O(N__18846),
            .I(N__18837));
    LocalMux I__4139 (
            .O(N__18843),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__4138 (
            .O(N__18840),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__4137 (
            .O(N__18837),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__4136 (
            .O(N__18830),
            .I(bfn_9_26_0_));
    InMux I__4135 (
            .O(N__18827),
            .I(N__18822));
    InMux I__4134 (
            .O(N__18826),
            .I(N__18819));
    InMux I__4133 (
            .O(N__18825),
            .I(N__18816));
    LocalMux I__4132 (
            .O(N__18822),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__4131 (
            .O(N__18819),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__4130 (
            .O(N__18816),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__4129 (
            .O(N__18809),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    CascadeMux I__4128 (
            .O(N__18806),
            .I(N__18801));
    CascadeMux I__4127 (
            .O(N__18805),
            .I(N__18798));
    InMux I__4126 (
            .O(N__18804),
            .I(N__18795));
    InMux I__4125 (
            .O(N__18801),
            .I(N__18790));
    InMux I__4124 (
            .O(N__18798),
            .I(N__18790));
    LocalMux I__4123 (
            .O(N__18795),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__4122 (
            .O(N__18790),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__4121 (
            .O(N__18785),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    CascadeMux I__4120 (
            .O(N__18782),
            .I(N__18777));
    CascadeMux I__4119 (
            .O(N__18781),
            .I(N__18774));
    InMux I__4118 (
            .O(N__18780),
            .I(N__18771));
    InMux I__4117 (
            .O(N__18777),
            .I(N__18766));
    InMux I__4116 (
            .O(N__18774),
            .I(N__18766));
    LocalMux I__4115 (
            .O(N__18771),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__4114 (
            .O(N__18766),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__4113 (
            .O(N__18761),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__4112 (
            .O(N__18758),
            .I(N__18753));
    InMux I__4111 (
            .O(N__18757),
            .I(N__18748));
    InMux I__4110 (
            .O(N__18756),
            .I(N__18748));
    LocalMux I__4109 (
            .O(N__18753),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__4108 (
            .O(N__18748),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__4107 (
            .O(N__18743),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__4106 (
            .O(N__18740),
            .I(N__18737));
    LocalMux I__4105 (
            .O(N__18737),
            .I(N__18732));
    InMux I__4104 (
            .O(N__18736),
            .I(N__18729));
    InMux I__4103 (
            .O(N__18735),
            .I(N__18726));
    Span4Mux_v I__4102 (
            .O(N__18732),
            .I(N__18721));
    LocalMux I__4101 (
            .O(N__18729),
            .I(N__18721));
    LocalMux I__4100 (
            .O(N__18726),
            .I(N__18718));
    Span4Mux_h I__4099 (
            .O(N__18721),
            .I(N__18715));
    Odrv12 I__4098 (
            .O(N__18718),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_5 ));
    Odrv4 I__4097 (
            .O(N__18715),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_5 ));
    InMux I__4096 (
            .O(N__18710),
            .I(N__18706));
    CascadeMux I__4095 (
            .O(N__18709),
            .I(N__18703));
    LocalMux I__4094 (
            .O(N__18706),
            .I(N__18700));
    InMux I__4093 (
            .O(N__18703),
            .I(N__18697));
    Span4Mux_v I__4092 (
            .O(N__18700),
            .I(N__18692));
    LocalMux I__4091 (
            .O(N__18697),
            .I(N__18692));
    Span4Mux_h I__4090 (
            .O(N__18692),
            .I(N__18688));
    InMux I__4089 (
            .O(N__18691),
            .I(N__18685));
    Span4Mux_h I__4088 (
            .O(N__18688),
            .I(N__18682));
    LocalMux I__4087 (
            .O(N__18685),
            .I(N__18679));
    Odrv4 I__4086 (
            .O(N__18682),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4 ));
    Odrv12 I__4085 (
            .O(N__18679),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4 ));
    CascadeMux I__4084 (
            .O(N__18674),
            .I(N__18670));
    InMux I__4083 (
            .O(N__18673),
            .I(N__18667));
    InMux I__4082 (
            .O(N__18670),
            .I(N__18664));
    LocalMux I__4081 (
            .O(N__18667),
            .I(measured_delay_hc_30));
    LocalMux I__4080 (
            .O(N__18664),
            .I(measured_delay_hc_30));
    InMux I__4079 (
            .O(N__18659),
            .I(N__18655));
    InMux I__4078 (
            .O(N__18658),
            .I(N__18652));
    LocalMux I__4077 (
            .O(N__18655),
            .I(measured_delay_hc_24));
    LocalMux I__4076 (
            .O(N__18652),
            .I(measured_delay_hc_24));
    InMux I__4075 (
            .O(N__18647),
            .I(N__18643));
    InMux I__4074 (
            .O(N__18646),
            .I(N__18640));
    LocalMux I__4073 (
            .O(N__18643),
            .I(measured_delay_hc_25));
    LocalMux I__4072 (
            .O(N__18640),
            .I(measured_delay_hc_25));
    InMux I__4071 (
            .O(N__18635),
            .I(N__18631));
    InMux I__4070 (
            .O(N__18634),
            .I(N__18628));
    LocalMux I__4069 (
            .O(N__18631),
            .I(measured_delay_hc_28));
    LocalMux I__4068 (
            .O(N__18628),
            .I(measured_delay_hc_28));
    InMux I__4067 (
            .O(N__18623),
            .I(N__18619));
    InMux I__4066 (
            .O(N__18622),
            .I(N__18616));
    LocalMux I__4065 (
            .O(N__18619),
            .I(measured_delay_hc_29));
    LocalMux I__4064 (
            .O(N__18616),
            .I(measured_delay_hc_29));
    InMux I__4063 (
            .O(N__18611),
            .I(N__18593));
    InMux I__4062 (
            .O(N__18610),
            .I(N__18593));
    InMux I__4061 (
            .O(N__18609),
            .I(N__18586));
    InMux I__4060 (
            .O(N__18608),
            .I(N__18586));
    InMux I__4059 (
            .O(N__18607),
            .I(N__18586));
    InMux I__4058 (
            .O(N__18606),
            .I(N__18573));
    InMux I__4057 (
            .O(N__18605),
            .I(N__18573));
    InMux I__4056 (
            .O(N__18604),
            .I(N__18573));
    InMux I__4055 (
            .O(N__18603),
            .I(N__18573));
    InMux I__4054 (
            .O(N__18602),
            .I(N__18573));
    InMux I__4053 (
            .O(N__18601),
            .I(N__18573));
    InMux I__4052 (
            .O(N__18600),
            .I(N__18566));
    InMux I__4051 (
            .O(N__18599),
            .I(N__18566));
    InMux I__4050 (
            .O(N__18598),
            .I(N__18566));
    LocalMux I__4049 (
            .O(N__18593),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__4048 (
            .O(N__18586),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__4047 (
            .O(N__18573),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__4046 (
            .O(N__18566),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    InMux I__4045 (
            .O(N__18557),
            .I(N__18553));
    InMux I__4044 (
            .O(N__18556),
            .I(N__18550));
    LocalMux I__4043 (
            .O(N__18553),
            .I(measured_delay_hc_23));
    LocalMux I__4042 (
            .O(N__18550),
            .I(measured_delay_hc_23));
    InMux I__4041 (
            .O(N__18545),
            .I(N__18541));
    InMux I__4040 (
            .O(N__18544),
            .I(N__18538));
    LocalMux I__4039 (
            .O(N__18541),
            .I(measured_delay_hc_27));
    LocalMux I__4038 (
            .O(N__18538),
            .I(measured_delay_hc_27));
    CascadeMux I__4037 (
            .O(N__18533),
            .I(N__18530));
    InMux I__4036 (
            .O(N__18530),
            .I(N__18527));
    LocalMux I__4035 (
            .O(N__18527),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ));
    InMux I__4034 (
            .O(N__18524),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__4033 (
            .O(N__18521),
            .I(N__18517));
    InMux I__4032 (
            .O(N__18520),
            .I(N__18514));
    LocalMux I__4031 (
            .O(N__18517),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__4030 (
            .O(N__18514),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__4029 (
            .O(N__18509),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__4028 (
            .O(N__18506),
            .I(N__18503));
    LocalMux I__4027 (
            .O(N__18503),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ));
    CEMux I__4026 (
            .O(N__18500),
            .I(N__18496));
    CEMux I__4025 (
            .O(N__18499),
            .I(N__18493));
    LocalMux I__4024 (
            .O(N__18496),
            .I(N__18488));
    LocalMux I__4023 (
            .O(N__18493),
            .I(N__18484));
    CEMux I__4022 (
            .O(N__18492),
            .I(N__18481));
    CEMux I__4021 (
            .O(N__18491),
            .I(N__18478));
    Span4Mux_v I__4020 (
            .O(N__18488),
            .I(N__18475));
    CEMux I__4019 (
            .O(N__18487),
            .I(N__18472));
    Span4Mux_h I__4018 (
            .O(N__18484),
            .I(N__18467));
    LocalMux I__4017 (
            .O(N__18481),
            .I(N__18467));
    LocalMux I__4016 (
            .O(N__18478),
            .I(N__18464));
    Span4Mux_h I__4015 (
            .O(N__18475),
            .I(N__18459));
    LocalMux I__4014 (
            .O(N__18472),
            .I(N__18459));
    Sp12to4 I__4013 (
            .O(N__18467),
            .I(N__18456));
    Span4Mux_h I__4012 (
            .O(N__18464),
            .I(N__18451));
    Span4Mux_h I__4011 (
            .O(N__18459),
            .I(N__18451));
    Odrv12 I__4010 (
            .O(N__18456),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__4009 (
            .O(N__18451),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    InMux I__4008 (
            .O(N__18446),
            .I(N__18443));
    LocalMux I__4007 (
            .O(N__18443),
            .I(N__18439));
    InMux I__4006 (
            .O(N__18442),
            .I(N__18435));
    Span4Mux_h I__4005 (
            .O(N__18439),
            .I(N__18432));
    InMux I__4004 (
            .O(N__18438),
            .I(N__18429));
    LocalMux I__4003 (
            .O(N__18435),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    Odrv4 I__4002 (
            .O(N__18432),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    LocalMux I__4001 (
            .O(N__18429),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    InMux I__4000 (
            .O(N__18422),
            .I(N__18419));
    LocalMux I__3999 (
            .O(N__18419),
            .I(N__18415));
    InMux I__3998 (
            .O(N__18418),
            .I(N__18411));
    Span4Mux_h I__3997 (
            .O(N__18415),
            .I(N__18408));
    InMux I__3996 (
            .O(N__18414),
            .I(N__18405));
    LocalMux I__3995 (
            .O(N__18411),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__3994 (
            .O(N__18408),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__3993 (
            .O(N__18405),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__3992 (
            .O(N__18398),
            .I(N__18395));
    LocalMux I__3991 (
            .O(N__18395),
            .I(N__18389));
    InMux I__3990 (
            .O(N__18394),
            .I(N__18384));
    InMux I__3989 (
            .O(N__18393),
            .I(N__18379));
    InMux I__3988 (
            .O(N__18392),
            .I(N__18379));
    Span4Mux_h I__3987 (
            .O(N__18389),
            .I(N__18376));
    InMux I__3986 (
            .O(N__18388),
            .I(N__18371));
    InMux I__3985 (
            .O(N__18387),
            .I(N__18371));
    LocalMux I__3984 (
            .O(N__18384),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__3983 (
            .O(N__18379),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__3982 (
            .O(N__18376),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__3981 (
            .O(N__18371),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__3980 (
            .O(N__18362),
            .I(N__18359));
    LocalMux I__3979 (
            .O(N__18359),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ));
    InMux I__3978 (
            .O(N__18356),
            .I(N__18353));
    LocalMux I__3977 (
            .O(N__18353),
            .I(\phase_controller_slave.start_timer_hc_0_sqmuxa ));
    CascadeMux I__3976 (
            .O(N__18350),
            .I(N__18344));
    CascadeMux I__3975 (
            .O(N__18349),
            .I(N__18341));
    CascadeMux I__3974 (
            .O(N__18348),
            .I(N__18338));
    InMux I__3973 (
            .O(N__18347),
            .I(N__18318));
    InMux I__3972 (
            .O(N__18344),
            .I(N__18309));
    InMux I__3971 (
            .O(N__18341),
            .I(N__18309));
    InMux I__3970 (
            .O(N__18338),
            .I(N__18309));
    InMux I__3969 (
            .O(N__18337),
            .I(N__18302));
    InMux I__3968 (
            .O(N__18336),
            .I(N__18302));
    InMux I__3967 (
            .O(N__18335),
            .I(N__18302));
    InMux I__3966 (
            .O(N__18334),
            .I(N__18285));
    InMux I__3965 (
            .O(N__18333),
            .I(N__18285));
    InMux I__3964 (
            .O(N__18332),
            .I(N__18285));
    InMux I__3963 (
            .O(N__18331),
            .I(N__18285));
    InMux I__3962 (
            .O(N__18330),
            .I(N__18285));
    InMux I__3961 (
            .O(N__18329),
            .I(N__18285));
    InMux I__3960 (
            .O(N__18328),
            .I(N__18285));
    InMux I__3959 (
            .O(N__18327),
            .I(N__18285));
    InMux I__3958 (
            .O(N__18326),
            .I(N__18274));
    InMux I__3957 (
            .O(N__18325),
            .I(N__18274));
    InMux I__3956 (
            .O(N__18324),
            .I(N__18274));
    InMux I__3955 (
            .O(N__18323),
            .I(N__18274));
    InMux I__3954 (
            .O(N__18322),
            .I(N__18274));
    InMux I__3953 (
            .O(N__18321),
            .I(N__18271));
    LocalMux I__3952 (
            .O(N__18318),
            .I(N__18268));
    InMux I__3951 (
            .O(N__18317),
            .I(N__18262));
    InMux I__3950 (
            .O(N__18316),
            .I(N__18262));
    LocalMux I__3949 (
            .O(N__18309),
            .I(N__18255));
    LocalMux I__3948 (
            .O(N__18302),
            .I(N__18255));
    LocalMux I__3947 (
            .O(N__18285),
            .I(N__18255));
    LocalMux I__3946 (
            .O(N__18274),
            .I(N__18248));
    LocalMux I__3945 (
            .O(N__18271),
            .I(N__18248));
    Span4Mux_h I__3944 (
            .O(N__18268),
            .I(N__18248));
    InMux I__3943 (
            .O(N__18267),
            .I(N__18245));
    LocalMux I__3942 (
            .O(N__18262),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv12 I__3941 (
            .O(N__18255),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__3940 (
            .O(N__18248),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__3939 (
            .O(N__18245),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    CascadeMux I__3938 (
            .O(N__18236),
            .I(N__18212));
    InMux I__3937 (
            .O(N__18235),
            .I(N__18198));
    InMux I__3936 (
            .O(N__18234),
            .I(N__18198));
    InMux I__3935 (
            .O(N__18233),
            .I(N__18198));
    InMux I__3934 (
            .O(N__18232),
            .I(N__18198));
    InMux I__3933 (
            .O(N__18231),
            .I(N__18198));
    InMux I__3932 (
            .O(N__18230),
            .I(N__18198));
    InMux I__3931 (
            .O(N__18229),
            .I(N__18181));
    InMux I__3930 (
            .O(N__18228),
            .I(N__18181));
    InMux I__3929 (
            .O(N__18227),
            .I(N__18181));
    InMux I__3928 (
            .O(N__18226),
            .I(N__18181));
    InMux I__3927 (
            .O(N__18225),
            .I(N__18181));
    InMux I__3926 (
            .O(N__18224),
            .I(N__18181));
    InMux I__3925 (
            .O(N__18223),
            .I(N__18181));
    InMux I__3924 (
            .O(N__18222),
            .I(N__18181));
    InMux I__3923 (
            .O(N__18221),
            .I(N__18170));
    InMux I__3922 (
            .O(N__18220),
            .I(N__18170));
    InMux I__3921 (
            .O(N__18219),
            .I(N__18170));
    InMux I__3920 (
            .O(N__18218),
            .I(N__18170));
    InMux I__3919 (
            .O(N__18217),
            .I(N__18170));
    InMux I__3918 (
            .O(N__18216),
            .I(N__18167));
    InMux I__3917 (
            .O(N__18215),
            .I(N__18164));
    InMux I__3916 (
            .O(N__18212),
            .I(N__18158));
    InMux I__3915 (
            .O(N__18211),
            .I(N__18158));
    LocalMux I__3914 (
            .O(N__18198),
            .I(N__18155));
    LocalMux I__3913 (
            .O(N__18181),
            .I(N__18146));
    LocalMux I__3912 (
            .O(N__18170),
            .I(N__18146));
    LocalMux I__3911 (
            .O(N__18167),
            .I(N__18146));
    LocalMux I__3910 (
            .O(N__18164),
            .I(N__18146));
    InMux I__3909 (
            .O(N__18163),
            .I(N__18143));
    LocalMux I__3908 (
            .O(N__18158),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv12 I__3907 (
            .O(N__18155),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__3906 (
            .O(N__18146),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__3905 (
            .O(N__18143),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    CascadeMux I__3904 (
            .O(N__18134),
            .I(N__18131));
    InMux I__3903 (
            .O(N__18131),
            .I(N__18128));
    LocalMux I__3902 (
            .O(N__18128),
            .I(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ));
    InMux I__3901 (
            .O(N__18125),
            .I(N__18122));
    LocalMux I__3900 (
            .O(N__18122),
            .I(\phase_controller_slave.N_21 ));
    IoInMux I__3899 (
            .O(N__18119),
            .I(N__18116));
    LocalMux I__3898 (
            .O(N__18116),
            .I(N__18113));
    Odrv12 I__3897 (
            .O(N__18113),
            .I(s3_phy_c));
    InMux I__3896 (
            .O(N__18110),
            .I(N__18106));
    CascadeMux I__3895 (
            .O(N__18109),
            .I(N__18103));
    LocalMux I__3894 (
            .O(N__18106),
            .I(N__18098));
    InMux I__3893 (
            .O(N__18103),
            .I(N__18091));
    InMux I__3892 (
            .O(N__18102),
            .I(N__18091));
    InMux I__3891 (
            .O(N__18101),
            .I(N__18091));
    Span4Mux_h I__3890 (
            .O(N__18098),
            .I(N__18088));
    LocalMux I__3889 (
            .O(N__18091),
            .I(N__18085));
    Span4Mux_h I__3888 (
            .O(N__18088),
            .I(N__18080));
    Span4Mux_h I__3887 (
            .O(N__18085),
            .I(N__18080));
    Odrv4 I__3886 (
            .O(N__18080),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    CascadeMux I__3885 (
            .O(N__18077),
            .I(N__18074));
    InMux I__3884 (
            .O(N__18074),
            .I(N__18071));
    LocalMux I__3883 (
            .O(N__18071),
            .I(N__18068));
    Span4Mux_h I__3882 (
            .O(N__18068),
            .I(N__18065));
    Odrv4 I__3881 (
            .O(N__18065),
            .I(\phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ));
    InMux I__3880 (
            .O(N__18062),
            .I(N__18057));
    InMux I__3879 (
            .O(N__18061),
            .I(N__18052));
    InMux I__3878 (
            .O(N__18060),
            .I(N__18052));
    LocalMux I__3877 (
            .O(N__18057),
            .I(N__18047));
    LocalMux I__3876 (
            .O(N__18052),
            .I(N__18044));
    InMux I__3875 (
            .O(N__18051),
            .I(N__18039));
    InMux I__3874 (
            .O(N__18050),
            .I(N__18039));
    Odrv12 I__3873 (
            .O(N__18047),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__3872 (
            .O(N__18044),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__3871 (
            .O(N__18039),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__3870 (
            .O(N__18032),
            .I(N__18028));
    InMux I__3869 (
            .O(N__18031),
            .I(N__18025));
    LocalMux I__3868 (
            .O(N__18028),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__3867 (
            .O(N__18025),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__3866 (
            .O(N__18020),
            .I(N__18017));
    LocalMux I__3865 (
            .O(N__18017),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ));
    InMux I__3864 (
            .O(N__18014),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__3863 (
            .O(N__18011),
            .I(N__18007));
    InMux I__3862 (
            .O(N__18010),
            .I(N__18004));
    LocalMux I__3861 (
            .O(N__18007),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__3860 (
            .O(N__18004),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__3859 (
            .O(N__17999),
            .I(N__17996));
    LocalMux I__3858 (
            .O(N__17996),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ));
    InMux I__3857 (
            .O(N__17993),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__3856 (
            .O(N__17990),
            .I(N__17986));
    InMux I__3855 (
            .O(N__17989),
            .I(N__17983));
    LocalMux I__3854 (
            .O(N__17986),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__3853 (
            .O(N__17983),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__3852 (
            .O(N__17978),
            .I(N__17975));
    LocalMux I__3851 (
            .O(N__17975),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ));
    InMux I__3850 (
            .O(N__17972),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__3849 (
            .O(N__17969),
            .I(N__17965));
    InMux I__3848 (
            .O(N__17968),
            .I(N__17962));
    LocalMux I__3847 (
            .O(N__17965),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__3846 (
            .O(N__17962),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__3845 (
            .O(N__17957),
            .I(N__17954));
    LocalMux I__3844 (
            .O(N__17954),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ));
    InMux I__3843 (
            .O(N__17951),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__3842 (
            .O(N__17948),
            .I(N__17944));
    InMux I__3841 (
            .O(N__17947),
            .I(N__17941));
    LocalMux I__3840 (
            .O(N__17944),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__3839 (
            .O(N__17941),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__3838 (
            .O(N__17936),
            .I(N__17933));
    LocalMux I__3837 (
            .O(N__17933),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ));
    InMux I__3836 (
            .O(N__17930),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__3835 (
            .O(N__17927),
            .I(N__17923));
    InMux I__3834 (
            .O(N__17926),
            .I(N__17920));
    LocalMux I__3833 (
            .O(N__17923),
            .I(N__17917));
    LocalMux I__3832 (
            .O(N__17920),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__3831 (
            .O(N__17917),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__3830 (
            .O(N__17912),
            .I(N__17909));
    LocalMux I__3829 (
            .O(N__17909),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ));
    InMux I__3828 (
            .O(N__17906),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__3827 (
            .O(N__17903),
            .I(N__17899));
    InMux I__3826 (
            .O(N__17902),
            .I(N__17896));
    LocalMux I__3825 (
            .O(N__17899),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__3824 (
            .O(N__17896),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__3823 (
            .O(N__17891),
            .I(N__17888));
    InMux I__3822 (
            .O(N__17888),
            .I(N__17885));
    LocalMux I__3821 (
            .O(N__17885),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ));
    InMux I__3820 (
            .O(N__17882),
            .I(bfn_9_19_0_));
    InMux I__3819 (
            .O(N__17879),
            .I(N__17875));
    InMux I__3818 (
            .O(N__17878),
            .I(N__17872));
    LocalMux I__3817 (
            .O(N__17875),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__3816 (
            .O(N__17872),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__3815 (
            .O(N__17867),
            .I(N__17863));
    InMux I__3814 (
            .O(N__17866),
            .I(N__17860));
    LocalMux I__3813 (
            .O(N__17863),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__3812 (
            .O(N__17860),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__3811 (
            .O(N__17855),
            .I(N__17852));
    InMux I__3810 (
            .O(N__17852),
            .I(N__17849));
    LocalMux I__3809 (
            .O(N__17849),
            .I(N__17846));
    Span4Mux_h I__3808 (
            .O(N__17846),
            .I(N__17843));
    Span4Mux_v I__3807 (
            .O(N__17843),
            .I(N__17840));
    Odrv4 I__3806 (
            .O(N__17840),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ));
    InMux I__3805 (
            .O(N__17837),
            .I(N__17834));
    LocalMux I__3804 (
            .O(N__17834),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ));
    InMux I__3803 (
            .O(N__17831),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__3802 (
            .O(N__17828),
            .I(N__17824));
    InMux I__3801 (
            .O(N__17827),
            .I(N__17821));
    LocalMux I__3800 (
            .O(N__17824),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__3799 (
            .O(N__17821),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__3798 (
            .O(N__17816),
            .I(N__17813));
    LocalMux I__3797 (
            .O(N__17813),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ));
    InMux I__3796 (
            .O(N__17810),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__3795 (
            .O(N__17807),
            .I(N__17803));
    InMux I__3794 (
            .O(N__17806),
            .I(N__17800));
    LocalMux I__3793 (
            .O(N__17803),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__3792 (
            .O(N__17800),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__3791 (
            .O(N__17795),
            .I(N__17792));
    LocalMux I__3790 (
            .O(N__17792),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ));
    InMux I__3789 (
            .O(N__17789),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__3788 (
            .O(N__17786),
            .I(N__17782));
    InMux I__3787 (
            .O(N__17785),
            .I(N__17779));
    LocalMux I__3786 (
            .O(N__17782),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__3785 (
            .O(N__17779),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__3784 (
            .O(N__17774),
            .I(N__17771));
    LocalMux I__3783 (
            .O(N__17771),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ));
    InMux I__3782 (
            .O(N__17768),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__3781 (
            .O(N__17765),
            .I(N__17761));
    InMux I__3780 (
            .O(N__17764),
            .I(N__17758));
    LocalMux I__3779 (
            .O(N__17761),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__3778 (
            .O(N__17758),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__3777 (
            .O(N__17753),
            .I(N__17750));
    LocalMux I__3776 (
            .O(N__17750),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ));
    InMux I__3775 (
            .O(N__17747),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__3774 (
            .O(N__17744),
            .I(N__17741));
    LocalMux I__3773 (
            .O(N__17741),
            .I(N__17738));
    Span4Mux_h I__3772 (
            .O(N__17738),
            .I(N__17734));
    InMux I__3771 (
            .O(N__17737),
            .I(N__17731));
    Odrv4 I__3770 (
            .O(N__17734),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__3769 (
            .O(N__17731),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__3768 (
            .O(N__17726),
            .I(N__17723));
    InMux I__3767 (
            .O(N__17723),
            .I(N__17720));
    LocalMux I__3766 (
            .O(N__17720),
            .I(N__17717));
    Odrv4 I__3765 (
            .O(N__17717),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ));
    InMux I__3764 (
            .O(N__17714),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__3763 (
            .O(N__17711),
            .I(N__17707));
    InMux I__3762 (
            .O(N__17710),
            .I(N__17704));
    LocalMux I__3761 (
            .O(N__17707),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__3760 (
            .O(N__17704),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__3759 (
            .O(N__17699),
            .I(N__17696));
    LocalMux I__3758 (
            .O(N__17696),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ));
    InMux I__3757 (
            .O(N__17693),
            .I(bfn_9_18_0_));
    InMux I__3756 (
            .O(N__17690),
            .I(N__17686));
    InMux I__3755 (
            .O(N__17689),
            .I(N__17683));
    LocalMux I__3754 (
            .O(N__17686),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__3753 (
            .O(N__17683),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__3752 (
            .O(N__17678),
            .I(N__17675));
    LocalMux I__3751 (
            .O(N__17675),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ));
    InMux I__3750 (
            .O(N__17672),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__3749 (
            .O(N__17669),
            .I(N__17665));
    InMux I__3748 (
            .O(N__17668),
            .I(N__17662));
    LocalMux I__3747 (
            .O(N__17665),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__3746 (
            .O(N__17662),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    CascadeMux I__3745 (
            .O(N__17657),
            .I(N__17654));
    InMux I__3744 (
            .O(N__17654),
            .I(N__17651));
    LocalMux I__3743 (
            .O(N__17651),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ));
    InMux I__3742 (
            .O(N__17648),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__3741 (
            .O(N__17645),
            .I(N__17641));
    InMux I__3740 (
            .O(N__17644),
            .I(N__17638));
    LocalMux I__3739 (
            .O(N__17641),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__3738 (
            .O(N__17638),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__3737 (
            .O(N__17633),
            .I(N__17630));
    LocalMux I__3736 (
            .O(N__17630),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ));
    InMux I__3735 (
            .O(N__17627),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__3734 (
            .O(N__17624),
            .I(N__17620));
    InMux I__3733 (
            .O(N__17623),
            .I(N__17617));
    LocalMux I__3732 (
            .O(N__17620),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__3731 (
            .O(N__17617),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__3730 (
            .O(N__17612),
            .I(N__17609));
    LocalMux I__3729 (
            .O(N__17609),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ));
    InMux I__3728 (
            .O(N__17606),
            .I(bfn_9_15_0_));
    InMux I__3727 (
            .O(N__17603),
            .I(N__17599));
    InMux I__3726 (
            .O(N__17602),
            .I(N__17596));
    LocalMux I__3725 (
            .O(N__17599),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__3724 (
            .O(N__17596),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__3723 (
            .O(N__17591),
            .I(N__17588));
    LocalMux I__3722 (
            .O(N__17588),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ));
    InMux I__3721 (
            .O(N__17585),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__3720 (
            .O(N__17582),
            .I(N__17578));
    InMux I__3719 (
            .O(N__17581),
            .I(N__17575));
    LocalMux I__3718 (
            .O(N__17578),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__3717 (
            .O(N__17575),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__3716 (
            .O(N__17570),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__3715 (
            .O(N__17567),
            .I(N__17564));
    LocalMux I__3714 (
            .O(N__17564),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ));
    CascadeMux I__3713 (
            .O(N__17561),
            .I(N__17553));
    CascadeMux I__3712 (
            .O(N__17560),
            .I(N__17550));
    CascadeMux I__3711 (
            .O(N__17559),
            .I(N__17547));
    CascadeMux I__3710 (
            .O(N__17558),
            .I(N__17544));
    CascadeMux I__3709 (
            .O(N__17557),
            .I(N__17536));
    CascadeMux I__3708 (
            .O(N__17556),
            .I(N__17533));
    InMux I__3707 (
            .O(N__17553),
            .I(N__17516));
    InMux I__3706 (
            .O(N__17550),
            .I(N__17516));
    InMux I__3705 (
            .O(N__17547),
            .I(N__17516));
    InMux I__3704 (
            .O(N__17544),
            .I(N__17516));
    InMux I__3703 (
            .O(N__17543),
            .I(N__17509));
    InMux I__3702 (
            .O(N__17542),
            .I(N__17509));
    InMux I__3701 (
            .O(N__17541),
            .I(N__17509));
    InMux I__3700 (
            .O(N__17540),
            .I(N__17501));
    InMux I__3699 (
            .O(N__17539),
            .I(N__17501));
    InMux I__3698 (
            .O(N__17536),
            .I(N__17496));
    InMux I__3697 (
            .O(N__17533),
            .I(N__17496));
    InMux I__3696 (
            .O(N__17532),
            .I(N__17479));
    InMux I__3695 (
            .O(N__17531),
            .I(N__17479));
    InMux I__3694 (
            .O(N__17530),
            .I(N__17479));
    InMux I__3693 (
            .O(N__17529),
            .I(N__17479));
    InMux I__3692 (
            .O(N__17528),
            .I(N__17479));
    InMux I__3691 (
            .O(N__17527),
            .I(N__17479));
    InMux I__3690 (
            .O(N__17526),
            .I(N__17479));
    InMux I__3689 (
            .O(N__17525),
            .I(N__17479));
    LocalMux I__3688 (
            .O(N__17516),
            .I(N__17474));
    LocalMux I__3687 (
            .O(N__17509),
            .I(N__17474));
    CascadeMux I__3686 (
            .O(N__17508),
            .I(N__17471));
    InMux I__3685 (
            .O(N__17507),
            .I(N__17466));
    InMux I__3684 (
            .O(N__17506),
            .I(N__17463));
    LocalMux I__3683 (
            .O(N__17501),
            .I(N__17460));
    LocalMux I__3682 (
            .O(N__17496),
            .I(N__17453));
    LocalMux I__3681 (
            .O(N__17479),
            .I(N__17453));
    Span4Mux_h I__3680 (
            .O(N__17474),
            .I(N__17453));
    InMux I__3679 (
            .O(N__17471),
            .I(N__17446));
    InMux I__3678 (
            .O(N__17470),
            .I(N__17446));
    InMux I__3677 (
            .O(N__17469),
            .I(N__17446));
    LocalMux I__3676 (
            .O(N__17466),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__3675 (
            .O(N__17463),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__3674 (
            .O(N__17460),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__3673 (
            .O(N__17453),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__3672 (
            .O(N__17446),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    CascadeMux I__3671 (
            .O(N__17435),
            .I(N__17432));
    InMux I__3670 (
            .O(N__17432),
            .I(N__17422));
    InMux I__3669 (
            .O(N__17431),
            .I(N__17407));
    InMux I__3668 (
            .O(N__17430),
            .I(N__17407));
    InMux I__3667 (
            .O(N__17429),
            .I(N__17407));
    InMux I__3666 (
            .O(N__17428),
            .I(N__17407));
    InMux I__3665 (
            .O(N__17427),
            .I(N__17407));
    InMux I__3664 (
            .O(N__17426),
            .I(N__17407));
    InMux I__3663 (
            .O(N__17425),
            .I(N__17407));
    LocalMux I__3662 (
            .O(N__17422),
            .I(N__17391));
    LocalMux I__3661 (
            .O(N__17407),
            .I(N__17388));
    InMux I__3660 (
            .O(N__17406),
            .I(N__17373));
    InMux I__3659 (
            .O(N__17405),
            .I(N__17373));
    InMux I__3658 (
            .O(N__17404),
            .I(N__17373));
    InMux I__3657 (
            .O(N__17403),
            .I(N__17373));
    InMux I__3656 (
            .O(N__17402),
            .I(N__17373));
    InMux I__3655 (
            .O(N__17401),
            .I(N__17373));
    InMux I__3654 (
            .O(N__17400),
            .I(N__17373));
    InMux I__3653 (
            .O(N__17399),
            .I(N__17367));
    InMux I__3652 (
            .O(N__17398),
            .I(N__17364));
    InMux I__3651 (
            .O(N__17397),
            .I(N__17355));
    InMux I__3650 (
            .O(N__17396),
            .I(N__17355));
    InMux I__3649 (
            .O(N__17395),
            .I(N__17355));
    InMux I__3648 (
            .O(N__17394),
            .I(N__17355));
    Span4Mux_v I__3647 (
            .O(N__17391),
            .I(N__17352));
    Span4Mux_h I__3646 (
            .O(N__17388),
            .I(N__17347));
    LocalMux I__3645 (
            .O(N__17373),
            .I(N__17347));
    InMux I__3644 (
            .O(N__17372),
            .I(N__17340));
    InMux I__3643 (
            .O(N__17371),
            .I(N__17340));
    InMux I__3642 (
            .O(N__17370),
            .I(N__17340));
    LocalMux I__3641 (
            .O(N__17367),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__3640 (
            .O(N__17364),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__3639 (
            .O(N__17355),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__3638 (
            .O(N__17352),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__3637 (
            .O(N__17347),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__3636 (
            .O(N__17340),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    CascadeMux I__3635 (
            .O(N__17327),
            .I(N__17324));
    InMux I__3634 (
            .O(N__17324),
            .I(N__17321));
    LocalMux I__3633 (
            .O(N__17321),
            .I(N__17318));
    Span4Mux_h I__3632 (
            .O(N__17318),
            .I(N__17315));
    Odrv4 I__3631 (
            .O(N__17315),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ));
    InMux I__3630 (
            .O(N__17312),
            .I(N__17308));
    InMux I__3629 (
            .O(N__17311),
            .I(N__17305));
    LocalMux I__3628 (
            .O(N__17308),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__3627 (
            .O(N__17305),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__3626 (
            .O(N__17300),
            .I(N__17297));
    LocalMux I__3625 (
            .O(N__17297),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ));
    InMux I__3624 (
            .O(N__17294),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__3623 (
            .O(N__17291),
            .I(N__17287));
    InMux I__3622 (
            .O(N__17290),
            .I(N__17284));
    LocalMux I__3621 (
            .O(N__17287),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__3620 (
            .O(N__17284),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__3619 (
            .O(N__17279),
            .I(N__17276));
    LocalMux I__3618 (
            .O(N__17276),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ));
    InMux I__3617 (
            .O(N__17273),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__3616 (
            .O(N__17270),
            .I(N__17266));
    InMux I__3615 (
            .O(N__17269),
            .I(N__17263));
    LocalMux I__3614 (
            .O(N__17266),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__3613 (
            .O(N__17263),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__3612 (
            .O(N__17258),
            .I(N__17255));
    LocalMux I__3611 (
            .O(N__17255),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ));
    InMux I__3610 (
            .O(N__17252),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__3609 (
            .O(N__17249),
            .I(N__17245));
    InMux I__3608 (
            .O(N__17248),
            .I(N__17242));
    LocalMux I__3607 (
            .O(N__17245),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__3606 (
            .O(N__17242),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__3605 (
            .O(N__17237),
            .I(N__17234));
    LocalMux I__3604 (
            .O(N__17234),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ));
    InMux I__3603 (
            .O(N__17231),
            .I(bfn_9_14_0_));
    InMux I__3602 (
            .O(N__17228),
            .I(N__17224));
    InMux I__3601 (
            .O(N__17227),
            .I(N__17221));
    LocalMux I__3600 (
            .O(N__17224),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__3599 (
            .O(N__17221),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    CascadeMux I__3598 (
            .O(N__17216),
            .I(N__17213));
    InMux I__3597 (
            .O(N__17213),
            .I(N__17210));
    LocalMux I__3596 (
            .O(N__17210),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ));
    InMux I__3595 (
            .O(N__17207),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__3594 (
            .O(N__17204),
            .I(N__17200));
    InMux I__3593 (
            .O(N__17203),
            .I(N__17197));
    LocalMux I__3592 (
            .O(N__17200),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__3591 (
            .O(N__17197),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__3590 (
            .O(N__17192),
            .I(N__17189));
    LocalMux I__3589 (
            .O(N__17189),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ));
    InMux I__3588 (
            .O(N__17186),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__3587 (
            .O(N__17183),
            .I(N__17180));
    LocalMux I__3586 (
            .O(N__17180),
            .I(N__17176));
    InMux I__3585 (
            .O(N__17179),
            .I(N__17173));
    Span4Mux_h I__3584 (
            .O(N__17176),
            .I(N__17170));
    LocalMux I__3583 (
            .O(N__17173),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__3582 (
            .O(N__17170),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__3581 (
            .O(N__17165),
            .I(N__17162));
    LocalMux I__3580 (
            .O(N__17162),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ));
    InMux I__3579 (
            .O(N__17159),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__3578 (
            .O(N__17156),
            .I(N__17152));
    InMux I__3577 (
            .O(N__17155),
            .I(N__17149));
    LocalMux I__3576 (
            .O(N__17152),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__3575 (
            .O(N__17149),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    CascadeMux I__3574 (
            .O(N__17144),
            .I(N__17141));
    InMux I__3573 (
            .O(N__17141),
            .I(N__17138));
    LocalMux I__3572 (
            .O(N__17138),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ));
    InMux I__3571 (
            .O(N__17135),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__3570 (
            .O(N__17132),
            .I(N__17128));
    InMux I__3569 (
            .O(N__17131),
            .I(N__17125));
    LocalMux I__3568 (
            .O(N__17128),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__3567 (
            .O(N__17125),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__3566 (
            .O(N__17120),
            .I(N__17117));
    LocalMux I__3565 (
            .O(N__17117),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ));
    InMux I__3564 (
            .O(N__17114),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ));
    CascadeMux I__3563 (
            .O(N__17111),
            .I(N__17108));
    InMux I__3562 (
            .O(N__17108),
            .I(N__17105));
    LocalMux I__3561 (
            .O(N__17105),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__3560 (
            .O(N__17102),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__3559 (
            .O(N__17099),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__3558 (
            .O(N__17096),
            .I(N__17092));
    InMux I__3557 (
            .O(N__17095),
            .I(N__17087));
    InMux I__3556 (
            .O(N__17092),
            .I(N__17087));
    LocalMux I__3555 (
            .O(N__17087),
            .I(N__17084));
    Span4Mux_v I__3554 (
            .O(N__17084),
            .I(N__17080));
    InMux I__3553 (
            .O(N__17083),
            .I(N__17077));
    Odrv4 I__3552 (
            .O(N__17080),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    LocalMux I__3551 (
            .O(N__17077),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__3550 (
            .O(N__17072),
            .I(N__17068));
    InMux I__3549 (
            .O(N__17071),
            .I(N__17064));
    LocalMux I__3548 (
            .O(N__17068),
            .I(N__17061));
    InMux I__3547 (
            .O(N__17067),
            .I(N__17058));
    LocalMux I__3546 (
            .O(N__17064),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__3545 (
            .O(N__17061),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__3544 (
            .O(N__17058),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__3543 (
            .O(N__17051),
            .I(N__17048));
    InMux I__3542 (
            .O(N__17048),
            .I(N__17045));
    LocalMux I__3541 (
            .O(N__17045),
            .I(N__17042));
    Span4Mux_v I__3540 (
            .O(N__17042),
            .I(N__17039));
    Odrv4 I__3539 (
            .O(N__17039),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ));
    InMux I__3538 (
            .O(N__17036),
            .I(N__17032));
    InMux I__3537 (
            .O(N__17035),
            .I(N__17029));
    LocalMux I__3536 (
            .O(N__17032),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__3535 (
            .O(N__17029),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__3534 (
            .O(N__17024),
            .I(N__17021));
    LocalMux I__3533 (
            .O(N__17021),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ));
    InMux I__3532 (
            .O(N__17018),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__3531 (
            .O(N__17015),
            .I(N__17011));
    InMux I__3530 (
            .O(N__17014),
            .I(N__17008));
    LocalMux I__3529 (
            .O(N__17011),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__3528 (
            .O(N__17008),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__3527 (
            .O(N__17003),
            .I(N__17000));
    InMux I__3526 (
            .O(N__17000),
            .I(N__16997));
    LocalMux I__3525 (
            .O(N__16997),
            .I(N__16994));
    Odrv4 I__3524 (
            .O(N__16994),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ));
    InMux I__3523 (
            .O(N__16991),
            .I(N__16988));
    LocalMux I__3522 (
            .O(N__16988),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ));
    InMux I__3521 (
            .O(N__16985),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__3520 (
            .O(N__16982),
            .I(N__16978));
    InMux I__3519 (
            .O(N__16981),
            .I(N__16975));
    LocalMux I__3518 (
            .O(N__16978),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__3517 (
            .O(N__16975),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__3516 (
            .O(N__16970),
            .I(N__16967));
    LocalMux I__3515 (
            .O(N__16967),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ));
    InMux I__3514 (
            .O(N__16964),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__3513 (
            .O(N__16961),
            .I(N__16957));
    InMux I__3512 (
            .O(N__16960),
            .I(N__16954));
    LocalMux I__3511 (
            .O(N__16957),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__3510 (
            .O(N__16954),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__3509 (
            .O(N__16949),
            .I(N__16946));
    LocalMux I__3508 (
            .O(N__16946),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ));
    InMux I__3507 (
            .O(N__16943),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__3506 (
            .O(N__16940),
            .I(N__16936));
    InMux I__3505 (
            .O(N__16939),
            .I(N__16933));
    LocalMux I__3504 (
            .O(N__16936),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__3503 (
            .O(N__16933),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__3502 (
            .O(N__16928),
            .I(N__16925));
    LocalMux I__3501 (
            .O(N__16925),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ));
    InMux I__3500 (
            .O(N__16922),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ));
    CascadeMux I__3499 (
            .O(N__16919),
            .I(N__16916));
    InMux I__3498 (
            .O(N__16916),
            .I(N__16910));
    InMux I__3497 (
            .O(N__16915),
            .I(N__16910));
    LocalMux I__3496 (
            .O(N__16910),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__3495 (
            .O(N__16907),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__3494 (
            .O(N__16904),
            .I(N__16901));
    LocalMux I__3493 (
            .O(N__16901),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__3492 (
            .O(N__16898),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__3491 (
            .O(N__16895),
            .I(N__16892));
    LocalMux I__3490 (
            .O(N__16892),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__3489 (
            .O(N__16889),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__3488 (
            .O(N__16886),
            .I(N__16883));
    LocalMux I__3487 (
            .O(N__16883),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__3486 (
            .O(N__16880),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__3485 (
            .O(N__16877),
            .I(N__16874));
    InMux I__3484 (
            .O(N__16874),
            .I(N__16871));
    LocalMux I__3483 (
            .O(N__16871),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__3482 (
            .O(N__16868),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__3481 (
            .O(N__16865),
            .I(N__16862));
    LocalMux I__3480 (
            .O(N__16862),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__3479 (
            .O(N__16859),
            .I(bfn_8_29_0_));
    InMux I__3478 (
            .O(N__16856),
            .I(N__16853));
    LocalMux I__3477 (
            .O(N__16853),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__3476 (
            .O(N__16850),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__3475 (
            .O(N__16847),
            .I(N__16844));
    LocalMux I__3474 (
            .O(N__16844),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__3473 (
            .O(N__16841),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__3472 (
            .O(N__16838),
            .I(N__16835));
    InMux I__3471 (
            .O(N__16835),
            .I(N__16829));
    InMux I__3470 (
            .O(N__16834),
            .I(N__16826));
    InMux I__3469 (
            .O(N__16833),
            .I(N__16823));
    InMux I__3468 (
            .O(N__16832),
            .I(N__16820));
    LocalMux I__3467 (
            .O(N__16829),
            .I(N__16813));
    LocalMux I__3466 (
            .O(N__16826),
            .I(N__16813));
    LocalMux I__3465 (
            .O(N__16823),
            .I(N__16813));
    LocalMux I__3464 (
            .O(N__16820),
            .I(N__16810));
    Span4Mux_v I__3463 (
            .O(N__16813),
            .I(N__16807));
    Odrv4 I__3462 (
            .O(N__16810),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    Odrv4 I__3461 (
            .O(N__16807),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    InMux I__3460 (
            .O(N__16802),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__3459 (
            .O(N__16799),
            .I(N__16789));
    InMux I__3458 (
            .O(N__16798),
            .I(N__16786));
    InMux I__3457 (
            .O(N__16797),
            .I(N__16783));
    InMux I__3456 (
            .O(N__16796),
            .I(N__16774));
    InMux I__3455 (
            .O(N__16795),
            .I(N__16774));
    InMux I__3454 (
            .O(N__16794),
            .I(N__16774));
    InMux I__3453 (
            .O(N__16793),
            .I(N__16774));
    InMux I__3452 (
            .O(N__16792),
            .I(N__16769));
    InMux I__3451 (
            .O(N__16789),
            .I(N__16769));
    LocalMux I__3450 (
            .O(N__16786),
            .I(N__16762));
    LocalMux I__3449 (
            .O(N__16783),
            .I(N__16762));
    LocalMux I__3448 (
            .O(N__16774),
            .I(N__16762));
    LocalMux I__3447 (
            .O(N__16769),
            .I(N__16759));
    Odrv4 I__3446 (
            .O(N__16762),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    Odrv4 I__3445 (
            .O(N__16759),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    InMux I__3444 (
            .O(N__16754),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__3443 (
            .O(N__16751),
            .I(N__16748));
    InMux I__3442 (
            .O(N__16748),
            .I(N__16743));
    InMux I__3441 (
            .O(N__16747),
            .I(N__16740));
    CascadeMux I__3440 (
            .O(N__16746),
            .I(N__16737));
    LocalMux I__3439 (
            .O(N__16743),
            .I(N__16732));
    LocalMux I__3438 (
            .O(N__16740),
            .I(N__16732));
    InMux I__3437 (
            .O(N__16737),
            .I(N__16729));
    Odrv4 I__3436 (
            .O(N__16732),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    LocalMux I__3435 (
            .O(N__16729),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    InMux I__3434 (
            .O(N__16724),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__3433 (
            .O(N__16721),
            .I(N__16718));
    LocalMux I__3432 (
            .O(N__16718),
            .I(N__16714));
    InMux I__3431 (
            .O(N__16717),
            .I(N__16711));
    Span4Mux_h I__3430 (
            .O(N__16714),
            .I(N__16705));
    LocalMux I__3429 (
            .O(N__16711),
            .I(N__16705));
    InMux I__3428 (
            .O(N__16710),
            .I(N__16702));
    Odrv4 I__3427 (
            .O(N__16705),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    LocalMux I__3426 (
            .O(N__16702),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    InMux I__3425 (
            .O(N__16697),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__3424 (
            .O(N__16694),
            .I(N__16691));
    LocalMux I__3423 (
            .O(N__16691),
            .I(N__16687));
    InMux I__3422 (
            .O(N__16690),
            .I(N__16684));
    Span4Mux_h I__3421 (
            .O(N__16687),
            .I(N__16678));
    LocalMux I__3420 (
            .O(N__16684),
            .I(N__16678));
    InMux I__3419 (
            .O(N__16683),
            .I(N__16675));
    Odrv4 I__3418 (
            .O(N__16678),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    LocalMux I__3417 (
            .O(N__16675),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    InMux I__3416 (
            .O(N__16670),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__3415 (
            .O(N__16667),
            .I(N__16663));
    CascadeMux I__3414 (
            .O(N__16666),
            .I(N__16659));
    LocalMux I__3413 (
            .O(N__16663),
            .I(N__16656));
    InMux I__3412 (
            .O(N__16662),
            .I(N__16653));
    InMux I__3411 (
            .O(N__16659),
            .I(N__16650));
    Span4Mux_h I__3410 (
            .O(N__16656),
            .I(N__16643));
    LocalMux I__3409 (
            .O(N__16653),
            .I(N__16643));
    LocalMux I__3408 (
            .O(N__16650),
            .I(N__16643));
    Odrv4 I__3407 (
            .O(N__16643),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    InMux I__3406 (
            .O(N__16640),
            .I(bfn_8_28_0_));
    CascadeMux I__3405 (
            .O(N__16637),
            .I(N__16634));
    InMux I__3404 (
            .O(N__16634),
            .I(N__16630));
    InMux I__3403 (
            .O(N__16633),
            .I(N__16627));
    LocalMux I__3402 (
            .O(N__16630),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    LocalMux I__3401 (
            .O(N__16627),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__3400 (
            .O(N__16622),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__3399 (
            .O(N__16619),
            .I(N__16613));
    InMux I__3398 (
            .O(N__16618),
            .I(N__16613));
    LocalMux I__3397 (
            .O(N__16613),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__3396 (
            .O(N__16610),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__3395 (
            .O(N__16607),
            .I(N__16603));
    InMux I__3394 (
            .O(N__16606),
            .I(N__16600));
    InMux I__3393 (
            .O(N__16603),
            .I(N__16597));
    LocalMux I__3392 (
            .O(N__16600),
            .I(N__16593));
    LocalMux I__3391 (
            .O(N__16597),
            .I(N__16590));
    InMux I__3390 (
            .O(N__16596),
            .I(N__16587));
    Odrv4 I__3389 (
            .O(N__16593),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    Odrv4 I__3388 (
            .O(N__16590),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    LocalMux I__3387 (
            .O(N__16587),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    InMux I__3386 (
            .O(N__16580),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__3385 (
            .O(N__16577),
            .I(N__16574));
    LocalMux I__3384 (
            .O(N__16574),
            .I(N__16569));
    InMux I__3383 (
            .O(N__16573),
            .I(N__16566));
    InMux I__3382 (
            .O(N__16572),
            .I(N__16563));
    Odrv4 I__3381 (
            .O(N__16569),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    LocalMux I__3380 (
            .O(N__16566),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    LocalMux I__3379 (
            .O(N__16563),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    InMux I__3378 (
            .O(N__16556),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__3377 (
            .O(N__16553),
            .I(N__16550));
    LocalMux I__3376 (
            .O(N__16550),
            .I(N__16545));
    InMux I__3375 (
            .O(N__16549),
            .I(N__16540));
    InMux I__3374 (
            .O(N__16548),
            .I(N__16540));
    Odrv4 I__3373 (
            .O(N__16545),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__3372 (
            .O(N__16540),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    InMux I__3371 (
            .O(N__16535),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__3370 (
            .O(N__16532),
            .I(N__16528));
    CascadeMux I__3369 (
            .O(N__16531),
            .I(N__16525));
    LocalMux I__3368 (
            .O(N__16528),
            .I(N__16521));
    InMux I__3367 (
            .O(N__16525),
            .I(N__16516));
    InMux I__3366 (
            .O(N__16524),
            .I(N__16516));
    Odrv4 I__3365 (
            .O(N__16521),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    LocalMux I__3364 (
            .O(N__16516),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    InMux I__3363 (
            .O(N__16511),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__3362 (
            .O(N__16508),
            .I(N__16504));
    InMux I__3361 (
            .O(N__16507),
            .I(N__16500));
    InMux I__3360 (
            .O(N__16504),
            .I(N__16497));
    InMux I__3359 (
            .O(N__16503),
            .I(N__16494));
    LocalMux I__3358 (
            .O(N__16500),
            .I(N__16490));
    LocalMux I__3357 (
            .O(N__16497),
            .I(N__16485));
    LocalMux I__3356 (
            .O(N__16494),
            .I(N__16485));
    InMux I__3355 (
            .O(N__16493),
            .I(N__16482));
    Odrv4 I__3354 (
            .O(N__16490),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    Odrv12 I__3353 (
            .O(N__16485),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    LocalMux I__3352 (
            .O(N__16482),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    InMux I__3351 (
            .O(N__16475),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__3350 (
            .O(N__16472),
            .I(N__16469));
    LocalMux I__3349 (
            .O(N__16469),
            .I(N__16464));
    InMux I__3348 (
            .O(N__16468),
            .I(N__16459));
    InMux I__3347 (
            .O(N__16467),
            .I(N__16459));
    Odrv12 I__3346 (
            .O(N__16464),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    LocalMux I__3345 (
            .O(N__16459),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    InMux I__3344 (
            .O(N__16454),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__3343 (
            .O(N__16451),
            .I(N__16446));
    InMux I__3342 (
            .O(N__16450),
            .I(N__16441));
    InMux I__3341 (
            .O(N__16449),
            .I(N__16441));
    LocalMux I__3340 (
            .O(N__16446),
            .I(N__16438));
    LocalMux I__3339 (
            .O(N__16441),
            .I(N__16435));
    Odrv12 I__3338 (
            .O(N__16438),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    Odrv4 I__3337 (
            .O(N__16435),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    InMux I__3336 (
            .O(N__16430),
            .I(bfn_8_27_0_));
    InMux I__3335 (
            .O(N__16427),
            .I(N__16422));
    InMux I__3334 (
            .O(N__16426),
            .I(N__16419));
    InMux I__3333 (
            .O(N__16425),
            .I(N__16416));
    LocalMux I__3332 (
            .O(N__16422),
            .I(N__16413));
    LocalMux I__3331 (
            .O(N__16419),
            .I(N__16408));
    LocalMux I__3330 (
            .O(N__16416),
            .I(N__16408));
    Odrv12 I__3329 (
            .O(N__16413),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    Odrv12 I__3328 (
            .O(N__16408),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    InMux I__3327 (
            .O(N__16403),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__3326 (
            .O(N__16400),
            .I(N__16396));
    CascadeMux I__3325 (
            .O(N__16399),
            .I(N__16393));
    LocalMux I__3324 (
            .O(N__16396),
            .I(N__16389));
    InMux I__3323 (
            .O(N__16393),
            .I(N__16386));
    InMux I__3322 (
            .O(N__16392),
            .I(N__16383));
    Span4Mux_h I__3321 (
            .O(N__16389),
            .I(N__16378));
    LocalMux I__3320 (
            .O(N__16386),
            .I(N__16378));
    LocalMux I__3319 (
            .O(N__16383),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    Odrv4 I__3318 (
            .O(N__16378),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    InMux I__3317 (
            .O(N__16373),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__3316 (
            .O(N__16370),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2Z0Z_6_cascade_ ));
    InMux I__3315 (
            .O(N__16367),
            .I(N__16361));
    InMux I__3314 (
            .O(N__16366),
            .I(N__16361));
    LocalMux I__3313 (
            .O(N__16361),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_3 ));
    InMux I__3312 (
            .O(N__16358),
            .I(N__16354));
    InMux I__3311 (
            .O(N__16357),
            .I(N__16351));
    LocalMux I__3310 (
            .O(N__16354),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0 ));
    LocalMux I__3309 (
            .O(N__16351),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0 ));
    InMux I__3308 (
            .O(N__16346),
            .I(N__16339));
    InMux I__3307 (
            .O(N__16345),
            .I(N__16339));
    InMux I__3306 (
            .O(N__16344),
            .I(N__16336));
    LocalMux I__3305 (
            .O(N__16339),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ));
    LocalMux I__3304 (
            .O(N__16336),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ));
    InMux I__3303 (
            .O(N__16331),
            .I(N__16328));
    LocalMux I__3302 (
            .O(N__16328),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6 ));
    CascadeMux I__3301 (
            .O(N__16325),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9_cascade_ ));
    InMux I__3300 (
            .O(N__16322),
            .I(N__16319));
    LocalMux I__3299 (
            .O(N__16319),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12 ));
    InMux I__3298 (
            .O(N__16316),
            .I(N__16312));
    InMux I__3297 (
            .O(N__16315),
            .I(N__16309));
    LocalMux I__3296 (
            .O(N__16312),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_2 ));
    LocalMux I__3295 (
            .O(N__16309),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_2 ));
    CascadeMux I__3294 (
            .O(N__16304),
            .I(N__16301));
    InMux I__3293 (
            .O(N__16301),
            .I(N__16297));
    InMux I__3292 (
            .O(N__16300),
            .I(N__16294));
    LocalMux I__3291 (
            .O(N__16297),
            .I(N__16290));
    LocalMux I__3290 (
            .O(N__16294),
            .I(N__16287));
    InMux I__3289 (
            .O(N__16293),
            .I(N__16284));
    Odrv4 I__3288 (
            .O(N__16290),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    Odrv4 I__3287 (
            .O(N__16287),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    LocalMux I__3286 (
            .O(N__16284),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    CascadeMux I__3285 (
            .O(N__16277),
            .I(N__16274));
    InMux I__3284 (
            .O(N__16274),
            .I(N__16271));
    LocalMux I__3283 (
            .O(N__16271),
            .I(N__16267));
    InMux I__3282 (
            .O(N__16270),
            .I(N__16264));
    Span4Mux_h I__3281 (
            .O(N__16267),
            .I(N__16258));
    LocalMux I__3280 (
            .O(N__16264),
            .I(N__16258));
    InMux I__3279 (
            .O(N__16263),
            .I(N__16255));
    Odrv4 I__3278 (
            .O(N__16258),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    LocalMux I__3277 (
            .O(N__16255),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    InMux I__3276 (
            .O(N__16250),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__3275 (
            .O(N__16247),
            .I(N__16244));
    LocalMux I__3274 (
            .O(N__16244),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5FBM1Z0Z_9 ));
    CascadeMux I__3273 (
            .O(N__16241),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_cascade_ ));
    InMux I__3272 (
            .O(N__16238),
            .I(N__16235));
    LocalMux I__3271 (
            .O(N__16235),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3 ));
    CascadeMux I__3270 (
            .O(N__16232),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3_cascade_ ));
    CascadeMux I__3269 (
            .O(N__16229),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_cascade_ ));
    InMux I__3268 (
            .O(N__16226),
            .I(N__16223));
    LocalMux I__3267 (
            .O(N__16223),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2 ));
    CascadeMux I__3266 (
            .O(N__16220),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_cascade_ ));
    InMux I__3265 (
            .O(N__16217),
            .I(N__16211));
    InMux I__3264 (
            .O(N__16216),
            .I(N__16211));
    LocalMux I__3263 (
            .O(N__16211),
            .I(N__16208));
    Span4Mux_h I__3262 (
            .O(N__16208),
            .I(N__16205));
    Odrv4 I__3261 (
            .O(N__16205),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_2 ));
    InMux I__3260 (
            .O(N__16202),
            .I(N__16199));
    LocalMux I__3259 (
            .O(N__16199),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2Z0Z_6 ));
    CascadeMux I__3258 (
            .O(N__16196),
            .I(N__16191));
    InMux I__3257 (
            .O(N__16195),
            .I(N__16187));
    InMux I__3256 (
            .O(N__16194),
            .I(N__16178));
    InMux I__3255 (
            .O(N__16191),
            .I(N__16178));
    InMux I__3254 (
            .O(N__16190),
            .I(N__16178));
    LocalMux I__3253 (
            .O(N__16187),
            .I(N__16175));
    InMux I__3252 (
            .O(N__16186),
            .I(N__16172));
    InMux I__3251 (
            .O(N__16185),
            .I(N__16169));
    LocalMux I__3250 (
            .O(N__16178),
            .I(N__16166));
    Span4Mux_h I__3249 (
            .O(N__16175),
            .I(N__16163));
    LocalMux I__3248 (
            .O(N__16172),
            .I(N__16160));
    LocalMux I__3247 (
            .O(N__16169),
            .I(N__16155));
    Span4Mux_h I__3246 (
            .O(N__16166),
            .I(N__16155));
    Odrv4 I__3245 (
            .O(N__16163),
            .I(measured_delay_hc_9));
    Odrv4 I__3244 (
            .O(N__16160),
            .I(measured_delay_hc_9));
    Odrv4 I__3243 (
            .O(N__16155),
            .I(measured_delay_hc_9));
    InMux I__3242 (
            .O(N__16148),
            .I(N__16143));
    InMux I__3241 (
            .O(N__16147),
            .I(N__16140));
    CascadeMux I__3240 (
            .O(N__16146),
            .I(N__16135));
    LocalMux I__3239 (
            .O(N__16143),
            .I(N__16130));
    LocalMux I__3238 (
            .O(N__16140),
            .I(N__16130));
    InMux I__3237 (
            .O(N__16139),
            .I(N__16127));
    InMux I__3236 (
            .O(N__16138),
            .I(N__16124));
    InMux I__3235 (
            .O(N__16135),
            .I(N__16121));
    Span4Mux_h I__3234 (
            .O(N__16130),
            .I(N__16118));
    LocalMux I__3233 (
            .O(N__16127),
            .I(N__16113));
    LocalMux I__3232 (
            .O(N__16124),
            .I(N__16113));
    LocalMux I__3231 (
            .O(N__16121),
            .I(measured_delay_hc_7));
    Odrv4 I__3230 (
            .O(N__16118),
            .I(measured_delay_hc_7));
    Odrv12 I__3229 (
            .O(N__16113),
            .I(measured_delay_hc_7));
    CascadeMux I__3228 (
            .O(N__16106),
            .I(N__16103));
    InMux I__3227 (
            .O(N__16103),
            .I(N__16099));
    InMux I__3226 (
            .O(N__16102),
            .I(N__16096));
    LocalMux I__3225 (
            .O(N__16099),
            .I(N__16090));
    LocalMux I__3224 (
            .O(N__16096),
            .I(N__16087));
    InMux I__3223 (
            .O(N__16095),
            .I(N__16082));
    InMux I__3222 (
            .O(N__16094),
            .I(N__16082));
    InMux I__3221 (
            .O(N__16093),
            .I(N__16079));
    Span4Mux_h I__3220 (
            .O(N__16090),
            .I(N__16076));
    Span4Mux_v I__3219 (
            .O(N__16087),
            .I(N__16073));
    LocalMux I__3218 (
            .O(N__16082),
            .I(N__16070));
    LocalMux I__3217 (
            .O(N__16079),
            .I(measured_delay_hc_2));
    Odrv4 I__3216 (
            .O(N__16076),
            .I(measured_delay_hc_2));
    Odrv4 I__3215 (
            .O(N__16073),
            .I(measured_delay_hc_2));
    Odrv4 I__3214 (
            .O(N__16070),
            .I(measured_delay_hc_2));
    CascadeMux I__3213 (
            .O(N__16061),
            .I(N__16056));
    CascadeMux I__3212 (
            .O(N__16060),
            .I(N__16052));
    InMux I__3211 (
            .O(N__16059),
            .I(N__16049));
    InMux I__3210 (
            .O(N__16056),
            .I(N__16046));
    InMux I__3209 (
            .O(N__16055),
            .I(N__16042));
    InMux I__3208 (
            .O(N__16052),
            .I(N__16039));
    LocalMux I__3207 (
            .O(N__16049),
            .I(N__16036));
    LocalMux I__3206 (
            .O(N__16046),
            .I(N__16033));
    InMux I__3205 (
            .O(N__16045),
            .I(N__16030));
    LocalMux I__3204 (
            .O(N__16042),
            .I(N__16027));
    LocalMux I__3203 (
            .O(N__16039),
            .I(N__16018));
    Span4Mux_v I__3202 (
            .O(N__16036),
            .I(N__16018));
    Span4Mux_h I__3201 (
            .O(N__16033),
            .I(N__16018));
    LocalMux I__3200 (
            .O(N__16030),
            .I(N__16018));
    Odrv4 I__3199 (
            .O(N__16027),
            .I(measured_delay_hc_8));
    Odrv4 I__3198 (
            .O(N__16018),
            .I(measured_delay_hc_8));
    InMux I__3197 (
            .O(N__16013),
            .I(N__16010));
    LocalMux I__3196 (
            .O(N__16010),
            .I(N__16003));
    InMux I__3195 (
            .O(N__16009),
            .I(N__16000));
    CascadeMux I__3194 (
            .O(N__16008),
            .I(N__15997));
    InMux I__3193 (
            .O(N__16007),
            .I(N__15994));
    InMux I__3192 (
            .O(N__16006),
            .I(N__15991));
    Span4Mux_v I__3191 (
            .O(N__16003),
            .I(N__15986));
    LocalMux I__3190 (
            .O(N__16000),
            .I(N__15986));
    InMux I__3189 (
            .O(N__15997),
            .I(N__15983));
    LocalMux I__3188 (
            .O(N__15994),
            .I(N__15980));
    LocalMux I__3187 (
            .O(N__15991),
            .I(N__15977));
    Span4Mux_h I__3186 (
            .O(N__15986),
            .I(N__15974));
    LocalMux I__3185 (
            .O(N__15983),
            .I(measured_delay_hc_12));
    Odrv4 I__3184 (
            .O(N__15980),
            .I(measured_delay_hc_12));
    Odrv12 I__3183 (
            .O(N__15977),
            .I(measured_delay_hc_12));
    Odrv4 I__3182 (
            .O(N__15974),
            .I(measured_delay_hc_12));
    InMux I__3181 (
            .O(N__15965),
            .I(N__15962));
    LocalMux I__3180 (
            .O(N__15962),
            .I(N__15956));
    InMux I__3179 (
            .O(N__15961),
            .I(N__15953));
    InMux I__3178 (
            .O(N__15960),
            .I(N__15949));
    InMux I__3177 (
            .O(N__15959),
            .I(N__15946));
    Span4Mux_v I__3176 (
            .O(N__15956),
            .I(N__15941));
    LocalMux I__3175 (
            .O(N__15953),
            .I(N__15941));
    InMux I__3174 (
            .O(N__15952),
            .I(N__15938));
    LocalMux I__3173 (
            .O(N__15949),
            .I(N__15935));
    LocalMux I__3172 (
            .O(N__15946),
            .I(N__15932));
    Span4Mux_h I__3171 (
            .O(N__15941),
            .I(N__15929));
    LocalMux I__3170 (
            .O(N__15938),
            .I(measured_delay_hc_10));
    Odrv4 I__3169 (
            .O(N__15935),
            .I(measured_delay_hc_10));
    Odrv12 I__3168 (
            .O(N__15932),
            .I(measured_delay_hc_10));
    Odrv4 I__3167 (
            .O(N__15929),
            .I(measured_delay_hc_10));
    CascadeMux I__3166 (
            .O(N__15920),
            .I(N__15917));
    InMux I__3165 (
            .O(N__15917),
            .I(N__15908));
    InMux I__3164 (
            .O(N__15916),
            .I(N__15908));
    InMux I__3163 (
            .O(N__15915),
            .I(N__15908));
    LocalMux I__3162 (
            .O(N__15908),
            .I(N__15900));
    InMux I__3161 (
            .O(N__15907),
            .I(N__15897));
    CascadeMux I__3160 (
            .O(N__15906),
            .I(N__15889));
    CascadeMux I__3159 (
            .O(N__15905),
            .I(N__15886));
    InMux I__3158 (
            .O(N__15904),
            .I(N__15877));
    InMux I__3157 (
            .O(N__15903),
            .I(N__15877));
    Span4Mux_h I__3156 (
            .O(N__15900),
            .I(N__15866));
    LocalMux I__3155 (
            .O(N__15897),
            .I(N__15866));
    InMux I__3154 (
            .O(N__15896),
            .I(N__15861));
    InMux I__3153 (
            .O(N__15895),
            .I(N__15861));
    InMux I__3152 (
            .O(N__15894),
            .I(N__15856));
    InMux I__3151 (
            .O(N__15893),
            .I(N__15856));
    InMux I__3150 (
            .O(N__15892),
            .I(N__15847));
    InMux I__3149 (
            .O(N__15889),
            .I(N__15847));
    InMux I__3148 (
            .O(N__15886),
            .I(N__15847));
    InMux I__3147 (
            .O(N__15885),
            .I(N__15847));
    InMux I__3146 (
            .O(N__15884),
            .I(N__15844));
    InMux I__3145 (
            .O(N__15883),
            .I(N__15839));
    InMux I__3144 (
            .O(N__15882),
            .I(N__15839));
    LocalMux I__3143 (
            .O(N__15877),
            .I(N__15835));
    InMux I__3142 (
            .O(N__15876),
            .I(N__15824));
    InMux I__3141 (
            .O(N__15875),
            .I(N__15824));
    InMux I__3140 (
            .O(N__15874),
            .I(N__15824));
    InMux I__3139 (
            .O(N__15873),
            .I(N__15824));
    InMux I__3138 (
            .O(N__15872),
            .I(N__15824));
    InMux I__3137 (
            .O(N__15871),
            .I(N__15821));
    Span4Mux_h I__3136 (
            .O(N__15866),
            .I(N__15814));
    LocalMux I__3135 (
            .O(N__15861),
            .I(N__15814));
    LocalMux I__3134 (
            .O(N__15856),
            .I(N__15814));
    LocalMux I__3133 (
            .O(N__15847),
            .I(N__15807));
    LocalMux I__3132 (
            .O(N__15844),
            .I(N__15807));
    LocalMux I__3131 (
            .O(N__15839),
            .I(N__15807));
    InMux I__3130 (
            .O(N__15838),
            .I(N__15804));
    Span4Mux_v I__3129 (
            .O(N__15835),
            .I(N__15797));
    LocalMux I__3128 (
            .O(N__15824),
            .I(N__15797));
    LocalMux I__3127 (
            .O(N__15821),
            .I(N__15797));
    Span4Mux_v I__3126 (
            .O(N__15814),
            .I(N__15792));
    Span4Mux_v I__3125 (
            .O(N__15807),
            .I(N__15792));
    LocalMux I__3124 (
            .O(N__15804),
            .I(measured_delay_hc_31));
    Odrv4 I__3123 (
            .O(N__15797),
            .I(measured_delay_hc_31));
    Odrv4 I__3122 (
            .O(N__15792),
            .I(measured_delay_hc_31));
    InMux I__3121 (
            .O(N__15785),
            .I(N__15780));
    InMux I__3120 (
            .O(N__15784),
            .I(N__15775));
    CascadeMux I__3119 (
            .O(N__15783),
            .I(N__15772));
    LocalMux I__3118 (
            .O(N__15780),
            .I(N__15769));
    InMux I__3117 (
            .O(N__15779),
            .I(N__15766));
    InMux I__3116 (
            .O(N__15778),
            .I(N__15763));
    LocalMux I__3115 (
            .O(N__15775),
            .I(N__15760));
    InMux I__3114 (
            .O(N__15772),
            .I(N__15757));
    Span4Mux_h I__3113 (
            .O(N__15769),
            .I(N__15752));
    LocalMux I__3112 (
            .O(N__15766),
            .I(N__15752));
    LocalMux I__3111 (
            .O(N__15763),
            .I(N__15749));
    Span4Mux_h I__3110 (
            .O(N__15760),
            .I(N__15746));
    LocalMux I__3109 (
            .O(N__15757),
            .I(measured_delay_hc_11));
    Odrv4 I__3108 (
            .O(N__15752),
            .I(measured_delay_hc_11));
    Odrv12 I__3107 (
            .O(N__15749),
            .I(measured_delay_hc_11));
    Odrv4 I__3106 (
            .O(N__15746),
            .I(measured_delay_hc_11));
    CascadeMux I__3105 (
            .O(N__15737),
            .I(N__15726));
    CascadeMux I__3104 (
            .O(N__15736),
            .I(N__15723));
    CascadeMux I__3103 (
            .O(N__15735),
            .I(N__15720));
    CascadeMux I__3102 (
            .O(N__15734),
            .I(N__15717));
    CascadeMux I__3101 (
            .O(N__15733),
            .I(N__15711));
    CascadeMux I__3100 (
            .O(N__15732),
            .I(N__15707));
    CascadeMux I__3099 (
            .O(N__15731),
            .I(N__15704));
    InMux I__3098 (
            .O(N__15730),
            .I(N__15691));
    InMux I__3097 (
            .O(N__15729),
            .I(N__15691));
    InMux I__3096 (
            .O(N__15726),
            .I(N__15691));
    InMux I__3095 (
            .O(N__15723),
            .I(N__15678));
    InMux I__3094 (
            .O(N__15720),
            .I(N__15678));
    InMux I__3093 (
            .O(N__15717),
            .I(N__15678));
    InMux I__3092 (
            .O(N__15716),
            .I(N__15678));
    InMux I__3091 (
            .O(N__15715),
            .I(N__15678));
    InMux I__3090 (
            .O(N__15714),
            .I(N__15678));
    InMux I__3089 (
            .O(N__15711),
            .I(N__15673));
    InMux I__3088 (
            .O(N__15710),
            .I(N__15673));
    InMux I__3087 (
            .O(N__15707),
            .I(N__15666));
    InMux I__3086 (
            .O(N__15704),
            .I(N__15666));
    InMux I__3085 (
            .O(N__15703),
            .I(N__15666));
    CascadeMux I__3084 (
            .O(N__15702),
            .I(N__15662));
    CascadeMux I__3083 (
            .O(N__15701),
            .I(N__15659));
    CascadeMux I__3082 (
            .O(N__15700),
            .I(N__15656));
    CascadeMux I__3081 (
            .O(N__15699),
            .I(N__15653));
    InMux I__3080 (
            .O(N__15698),
            .I(N__15647));
    LocalMux I__3079 (
            .O(N__15691),
            .I(N__15644));
    LocalMux I__3078 (
            .O(N__15678),
            .I(N__15637));
    LocalMux I__3077 (
            .O(N__15673),
            .I(N__15637));
    LocalMux I__3076 (
            .O(N__15666),
            .I(N__15637));
    InMux I__3075 (
            .O(N__15665),
            .I(N__15634));
    InMux I__3074 (
            .O(N__15662),
            .I(N__15618));
    InMux I__3073 (
            .O(N__15659),
            .I(N__15618));
    InMux I__3072 (
            .O(N__15656),
            .I(N__15618));
    InMux I__3071 (
            .O(N__15653),
            .I(N__15618));
    InMux I__3070 (
            .O(N__15652),
            .I(N__15618));
    InMux I__3069 (
            .O(N__15651),
            .I(N__15618));
    InMux I__3068 (
            .O(N__15650),
            .I(N__15618));
    LocalMux I__3067 (
            .O(N__15647),
            .I(N__15615));
    Span4Mux_h I__3066 (
            .O(N__15644),
            .I(N__15608));
    Span4Mux_v I__3065 (
            .O(N__15637),
            .I(N__15608));
    LocalMux I__3064 (
            .O(N__15634),
            .I(N__15608));
    InMux I__3063 (
            .O(N__15633),
            .I(N__15605));
    LocalMux I__3062 (
            .O(N__15618),
            .I(N__15602));
    Span4Mux_h I__3061 (
            .O(N__15615),
            .I(N__15599));
    Span4Mux_h I__3060 (
            .O(N__15608),
            .I(N__15596));
    LocalMux I__3059 (
            .O(N__15605),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv12 I__3058 (
            .O(N__15602),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__3057 (
            .O(N__15599),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__3056 (
            .O(N__15596),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    InMux I__3055 (
            .O(N__15587),
            .I(N__15581));
    InMux I__3054 (
            .O(N__15586),
            .I(N__15581));
    LocalMux I__3053 (
            .O(N__15581),
            .I(N__15573));
    InMux I__3052 (
            .O(N__15580),
            .I(N__15566));
    InMux I__3051 (
            .O(N__15579),
            .I(N__15566));
    InMux I__3050 (
            .O(N__15578),
            .I(N__15566));
    InMux I__3049 (
            .O(N__15577),
            .I(N__15563));
    InMux I__3048 (
            .O(N__15576),
            .I(N__15555));
    Span4Mux_h I__3047 (
            .O(N__15573),
            .I(N__15548));
    LocalMux I__3046 (
            .O(N__15566),
            .I(N__15548));
    LocalMux I__3045 (
            .O(N__15563),
            .I(N__15545));
    InMux I__3044 (
            .O(N__15562),
            .I(N__15534));
    InMux I__3043 (
            .O(N__15561),
            .I(N__15534));
    InMux I__3042 (
            .O(N__15560),
            .I(N__15534));
    InMux I__3041 (
            .O(N__15559),
            .I(N__15534));
    InMux I__3040 (
            .O(N__15558),
            .I(N__15534));
    LocalMux I__3039 (
            .O(N__15555),
            .I(N__15527));
    InMux I__3038 (
            .O(N__15554),
            .I(N__15522));
    InMux I__3037 (
            .O(N__15553),
            .I(N__15522));
    Span4Mux_v I__3036 (
            .O(N__15548),
            .I(N__15515));
    Span4Mux_v I__3035 (
            .O(N__15545),
            .I(N__15515));
    LocalMux I__3034 (
            .O(N__15534),
            .I(N__15515));
    InMux I__3033 (
            .O(N__15533),
            .I(N__15506));
    InMux I__3032 (
            .O(N__15532),
            .I(N__15506));
    InMux I__3031 (
            .O(N__15531),
            .I(N__15506));
    InMux I__3030 (
            .O(N__15530),
            .I(N__15506));
    Odrv12 I__3029 (
            .O(N__15527),
            .I(\phase_controller_inst1.stoper_hc.un1_start ));
    LocalMux I__3028 (
            .O(N__15522),
            .I(\phase_controller_inst1.stoper_hc.un1_start ));
    Odrv4 I__3027 (
            .O(N__15515),
            .I(\phase_controller_inst1.stoper_hc.un1_start ));
    LocalMux I__3026 (
            .O(N__15506),
            .I(\phase_controller_inst1.stoper_hc.un1_start ));
    InMux I__3025 (
            .O(N__15497),
            .I(N__15494));
    LocalMux I__3024 (
            .O(N__15494),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__3023 (
            .O(N__15491),
            .I(N__15488));
    LocalMux I__3022 (
            .O(N__15488),
            .I(N__15485));
    Odrv4 I__3021 (
            .O(N__15485),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__3020 (
            .O(N__15482),
            .I(N__15479));
    LocalMux I__3019 (
            .O(N__15479),
            .I(N__15476));
    Odrv4 I__3018 (
            .O(N__15476),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    InMux I__3017 (
            .O(N__15473),
            .I(N__15470));
    LocalMux I__3016 (
            .O(N__15470),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    InMux I__3015 (
            .O(N__15467),
            .I(N__15457));
    InMux I__3014 (
            .O(N__15466),
            .I(N__15457));
    InMux I__3013 (
            .O(N__15465),
            .I(N__15440));
    InMux I__3012 (
            .O(N__15464),
            .I(N__15440));
    InMux I__3011 (
            .O(N__15463),
            .I(N__15440));
    InMux I__3010 (
            .O(N__15462),
            .I(N__15440));
    LocalMux I__3009 (
            .O(N__15457),
            .I(N__15431));
    InMux I__3008 (
            .O(N__15456),
            .I(N__15420));
    InMux I__3007 (
            .O(N__15455),
            .I(N__15420));
    InMux I__3006 (
            .O(N__15454),
            .I(N__15420));
    InMux I__3005 (
            .O(N__15453),
            .I(N__15420));
    InMux I__3004 (
            .O(N__15452),
            .I(N__15420));
    InMux I__3003 (
            .O(N__15451),
            .I(N__15413));
    InMux I__3002 (
            .O(N__15450),
            .I(N__15413));
    InMux I__3001 (
            .O(N__15449),
            .I(N__15413));
    LocalMux I__3000 (
            .O(N__15440),
            .I(N__15408));
    InMux I__2999 (
            .O(N__15439),
            .I(N__15395));
    InMux I__2998 (
            .O(N__15438),
            .I(N__15395));
    InMux I__2997 (
            .O(N__15437),
            .I(N__15395));
    InMux I__2996 (
            .O(N__15436),
            .I(N__15395));
    InMux I__2995 (
            .O(N__15435),
            .I(N__15395));
    InMux I__2994 (
            .O(N__15434),
            .I(N__15395));
    Span4Mux_h I__2993 (
            .O(N__15431),
            .I(N__15388));
    LocalMux I__2992 (
            .O(N__15420),
            .I(N__15388));
    LocalMux I__2991 (
            .O(N__15413),
            .I(N__15388));
    InMux I__2990 (
            .O(N__15412),
            .I(N__15383));
    InMux I__2989 (
            .O(N__15411),
            .I(N__15383));
    Odrv4 I__2988 (
            .O(N__15408),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_d ));
    LocalMux I__2987 (
            .O(N__15395),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_d ));
    Odrv4 I__2986 (
            .O(N__15388),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_d ));
    LocalMux I__2985 (
            .O(N__15383),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_d ));
    CascadeMux I__2984 (
            .O(N__15374),
            .I(N__15370));
    CascadeMux I__2983 (
            .O(N__15373),
            .I(N__15367));
    InMux I__2982 (
            .O(N__15370),
            .I(N__15362));
    InMux I__2981 (
            .O(N__15367),
            .I(N__15362));
    LocalMux I__2980 (
            .O(N__15362),
            .I(N__15346));
    InMux I__2979 (
            .O(N__15361),
            .I(N__15337));
    InMux I__2978 (
            .O(N__15360),
            .I(N__15337));
    InMux I__2977 (
            .O(N__15359),
            .I(N__15337));
    InMux I__2976 (
            .O(N__15358),
            .I(N__15337));
    CascadeMux I__2975 (
            .O(N__15357),
            .I(N__15334));
    InMux I__2974 (
            .O(N__15356),
            .I(N__15318));
    InMux I__2973 (
            .O(N__15355),
            .I(N__15318));
    InMux I__2972 (
            .O(N__15354),
            .I(N__15318));
    InMux I__2971 (
            .O(N__15353),
            .I(N__15318));
    InMux I__2970 (
            .O(N__15352),
            .I(N__15318));
    InMux I__2969 (
            .O(N__15351),
            .I(N__15311));
    InMux I__2968 (
            .O(N__15350),
            .I(N__15311));
    InMux I__2967 (
            .O(N__15349),
            .I(N__15311));
    Span4Mux_v I__2966 (
            .O(N__15346),
            .I(N__15306));
    LocalMux I__2965 (
            .O(N__15337),
            .I(N__15303));
    InMux I__2964 (
            .O(N__15334),
            .I(N__15290));
    InMux I__2963 (
            .O(N__15333),
            .I(N__15290));
    InMux I__2962 (
            .O(N__15332),
            .I(N__15290));
    InMux I__2961 (
            .O(N__15331),
            .I(N__15290));
    InMux I__2960 (
            .O(N__15330),
            .I(N__15290));
    InMux I__2959 (
            .O(N__15329),
            .I(N__15290));
    LocalMux I__2958 (
            .O(N__15318),
            .I(N__15285));
    LocalMux I__2957 (
            .O(N__15311),
            .I(N__15285));
    InMux I__2956 (
            .O(N__15310),
            .I(N__15280));
    InMux I__2955 (
            .O(N__15309),
            .I(N__15280));
    Odrv4 I__2954 (
            .O(N__15306),
            .I(\phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0 ));
    Odrv4 I__2953 (
            .O(N__15303),
            .I(\phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0 ));
    LocalMux I__2952 (
            .O(N__15290),
            .I(\phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0 ));
    Odrv4 I__2951 (
            .O(N__15285),
            .I(\phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0 ));
    LocalMux I__2950 (
            .O(N__15280),
            .I(\phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0 ));
    InMux I__2949 (
            .O(N__15269),
            .I(N__15266));
    LocalMux I__2948 (
            .O(N__15266),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__2947 (
            .O(N__15263),
            .I(N__15251));
    CascadeMux I__2946 (
            .O(N__15262),
            .I(N__15248));
    CascadeMux I__2945 (
            .O(N__15261),
            .I(N__15245));
    CascadeMux I__2944 (
            .O(N__15260),
            .I(N__15242));
    CascadeMux I__2943 (
            .O(N__15259),
            .I(N__15239));
    InMux I__2942 (
            .O(N__15258),
            .I(N__15224));
    InMux I__2941 (
            .O(N__15257),
            .I(N__15215));
    InMux I__2940 (
            .O(N__15256),
            .I(N__15215));
    InMux I__2939 (
            .O(N__15255),
            .I(N__15215));
    InMux I__2938 (
            .O(N__15254),
            .I(N__15215));
    InMux I__2937 (
            .O(N__15251),
            .I(N__15212));
    InMux I__2936 (
            .O(N__15248),
            .I(N__15203));
    InMux I__2935 (
            .O(N__15245),
            .I(N__15203));
    InMux I__2934 (
            .O(N__15242),
            .I(N__15203));
    InMux I__2933 (
            .O(N__15239),
            .I(N__15203));
    InMux I__2932 (
            .O(N__15238),
            .I(N__15200));
    InMux I__2931 (
            .O(N__15237),
            .I(N__15197));
    InMux I__2930 (
            .O(N__15236),
            .I(N__15190));
    InMux I__2929 (
            .O(N__15235),
            .I(N__15190));
    InMux I__2928 (
            .O(N__15234),
            .I(N__15190));
    InMux I__2927 (
            .O(N__15233),
            .I(N__15175));
    InMux I__2926 (
            .O(N__15232),
            .I(N__15175));
    InMux I__2925 (
            .O(N__15231),
            .I(N__15175));
    InMux I__2924 (
            .O(N__15230),
            .I(N__15175));
    InMux I__2923 (
            .O(N__15229),
            .I(N__15175));
    InMux I__2922 (
            .O(N__15228),
            .I(N__15175));
    InMux I__2921 (
            .O(N__15227),
            .I(N__15175));
    LocalMux I__2920 (
            .O(N__15224),
            .I(N__15172));
    LocalMux I__2919 (
            .O(N__15215),
            .I(N__15165));
    LocalMux I__2918 (
            .O(N__15212),
            .I(N__15165));
    LocalMux I__2917 (
            .O(N__15203),
            .I(N__15158));
    LocalMux I__2916 (
            .O(N__15200),
            .I(N__15158));
    LocalMux I__2915 (
            .O(N__15197),
            .I(N__15158));
    LocalMux I__2914 (
            .O(N__15190),
            .I(N__15153));
    LocalMux I__2913 (
            .O(N__15175),
            .I(N__15153));
    Span4Mux_h I__2912 (
            .O(N__15172),
            .I(N__15150));
    InMux I__2911 (
            .O(N__15171),
            .I(N__15147));
    InMux I__2910 (
            .O(N__15170),
            .I(N__15144));
    Span4Mux_v I__2909 (
            .O(N__15165),
            .I(N__15141));
    Span12Mux_h I__2908 (
            .O(N__15158),
            .I(N__15138));
    Span4Mux_v I__2907 (
            .O(N__15153),
            .I(N__15131));
    Span4Mux_h I__2906 (
            .O(N__15150),
            .I(N__15131));
    LocalMux I__2905 (
            .O(N__15147),
            .I(N__15131));
    LocalMux I__2904 (
            .O(N__15144),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__2903 (
            .O(N__15141),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv12 I__2902 (
            .O(N__15138),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__2901 (
            .O(N__15131),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    InMux I__2900 (
            .O(N__15122),
            .I(N__15119));
    LocalMux I__2899 (
            .O(N__15119),
            .I(N__15115));
    InMux I__2898 (
            .O(N__15118),
            .I(N__15112));
    Span4Mux_v I__2897 (
            .O(N__15115),
            .I(N__15106));
    LocalMux I__2896 (
            .O(N__15112),
            .I(N__15106));
    InMux I__2895 (
            .O(N__15111),
            .I(N__15103));
    Span4Mux_h I__2894 (
            .O(N__15106),
            .I(N__15098));
    LocalMux I__2893 (
            .O(N__15103),
            .I(N__15095));
    InMux I__2892 (
            .O(N__15102),
            .I(N__15090));
    InMux I__2891 (
            .O(N__15101),
            .I(N__15090));
    Odrv4 I__2890 (
            .O(N__15098),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__2889 (
            .O(N__15095),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__2888 (
            .O(N__15090),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__2887 (
            .O(N__15083),
            .I(N__15080));
    InMux I__2886 (
            .O(N__15080),
            .I(N__15058));
    InMux I__2885 (
            .O(N__15079),
            .I(N__15053));
    InMux I__2884 (
            .O(N__15078),
            .I(N__15053));
    InMux I__2883 (
            .O(N__15077),
            .I(N__15036));
    InMux I__2882 (
            .O(N__15076),
            .I(N__15036));
    InMux I__2881 (
            .O(N__15075),
            .I(N__15036));
    InMux I__2880 (
            .O(N__15074),
            .I(N__15036));
    InMux I__2879 (
            .O(N__15073),
            .I(N__15036));
    InMux I__2878 (
            .O(N__15072),
            .I(N__15036));
    InMux I__2877 (
            .O(N__15071),
            .I(N__15036));
    InMux I__2876 (
            .O(N__15070),
            .I(N__15036));
    InMux I__2875 (
            .O(N__15069),
            .I(N__15033));
    InMux I__2874 (
            .O(N__15068),
            .I(N__15016));
    InMux I__2873 (
            .O(N__15067),
            .I(N__15016));
    InMux I__2872 (
            .O(N__15066),
            .I(N__15016));
    InMux I__2871 (
            .O(N__15065),
            .I(N__15016));
    InMux I__2870 (
            .O(N__15064),
            .I(N__15016));
    InMux I__2869 (
            .O(N__15063),
            .I(N__15016));
    InMux I__2868 (
            .O(N__15062),
            .I(N__15016));
    InMux I__2867 (
            .O(N__15061),
            .I(N__15016));
    LocalMux I__2866 (
            .O(N__15058),
            .I(N__15009));
    LocalMux I__2865 (
            .O(N__15053),
            .I(N__15009));
    LocalMux I__2864 (
            .O(N__15036),
            .I(N__15009));
    LocalMux I__2863 (
            .O(N__15033),
            .I(N__15003));
    LocalMux I__2862 (
            .O(N__15016),
            .I(N__15003));
    Span4Mux_v I__2861 (
            .O(N__15009),
            .I(N__14998));
    CascadeMux I__2860 (
            .O(N__15008),
            .I(N__14994));
    Span4Mux_v I__2859 (
            .O(N__15003),
            .I(N__14991));
    InMux I__2858 (
            .O(N__15002),
            .I(N__14988));
    InMux I__2857 (
            .O(N__15001),
            .I(N__14985));
    Span4Mux_h I__2856 (
            .O(N__14998),
            .I(N__14982));
    InMux I__2855 (
            .O(N__14997),
            .I(N__14979));
    InMux I__2854 (
            .O(N__14994),
            .I(N__14976));
    Sp12to4 I__2853 (
            .O(N__14991),
            .I(N__14971));
    LocalMux I__2852 (
            .O(N__14988),
            .I(N__14971));
    LocalMux I__2851 (
            .O(N__14985),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__2850 (
            .O(N__14982),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__2849 (
            .O(N__14979),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__2848 (
            .O(N__14976),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv12 I__2847 (
            .O(N__14971),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    InMux I__2846 (
            .O(N__14960),
            .I(N__14957));
    LocalMux I__2845 (
            .O(N__14957),
            .I(N__14954));
    Span4Mux_h I__2844 (
            .O(N__14954),
            .I(N__14950));
    CascadeMux I__2843 (
            .O(N__14953),
            .I(N__14947));
    Span4Mux_h I__2842 (
            .O(N__14950),
            .I(N__14942));
    InMux I__2841 (
            .O(N__14947),
            .I(N__14937));
    InMux I__2840 (
            .O(N__14946),
            .I(N__14937));
    InMux I__2839 (
            .O(N__14945),
            .I(N__14934));
    Odrv4 I__2838 (
            .O(N__14942),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    LocalMux I__2837 (
            .O(N__14937),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    LocalMux I__2836 (
            .O(N__14934),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    InMux I__2835 (
            .O(N__14927),
            .I(N__14924));
    LocalMux I__2834 (
            .O(N__14924),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ));
    CascadeMux I__2833 (
            .O(N__14921),
            .I(\phase_controller_inst1.stoper_tr.time_passed11_cascade_ ));
    CascadeMux I__2832 (
            .O(N__14918),
            .I(N__14915));
    InMux I__2831 (
            .O(N__14915),
            .I(N__14912));
    LocalMux I__2830 (
            .O(N__14912),
            .I(\phase_controller_slave.stoper_tr.time_passed_1_sqmuxa ));
    InMux I__2829 (
            .O(N__14909),
            .I(N__14906));
    LocalMux I__2828 (
            .O(N__14906),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_0_0 ));
    InMux I__2827 (
            .O(N__14903),
            .I(N__14897));
    InMux I__2826 (
            .O(N__14902),
            .I(N__14897));
    LocalMux I__2825 (
            .O(N__14897),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ));
    InMux I__2824 (
            .O(N__14894),
            .I(N__14891));
    LocalMux I__2823 (
            .O(N__14891),
            .I(N__14888));
    Span4Mux_v I__2822 (
            .O(N__14888),
            .I(N__14885));
    Sp12to4 I__2821 (
            .O(N__14885),
            .I(N__14882));
    Span12Mux_h I__2820 (
            .O(N__14882),
            .I(N__14879));
    Odrv12 I__2819 (
            .O(N__14879),
            .I(il_min_comp2_c));
    InMux I__2818 (
            .O(N__14876),
            .I(N__14870));
    InMux I__2817 (
            .O(N__14875),
            .I(N__14867));
    InMux I__2816 (
            .O(N__14874),
            .I(N__14864));
    InMux I__2815 (
            .O(N__14873),
            .I(N__14860));
    LocalMux I__2814 (
            .O(N__14870),
            .I(N__14857));
    LocalMux I__2813 (
            .O(N__14867),
            .I(N__14852));
    LocalMux I__2812 (
            .O(N__14864),
            .I(N__14852));
    InMux I__2811 (
            .O(N__14863),
            .I(N__14849));
    LocalMux I__2810 (
            .O(N__14860),
            .I(N__14846));
    Span4Mux_h I__2809 (
            .O(N__14857),
            .I(N__14843));
    Span4Mux_h I__2808 (
            .O(N__14852),
            .I(N__14840));
    LocalMux I__2807 (
            .O(N__14849),
            .I(measured_delay_hc_16));
    Odrv4 I__2806 (
            .O(N__14846),
            .I(measured_delay_hc_16));
    Odrv4 I__2805 (
            .O(N__14843),
            .I(measured_delay_hc_16));
    Odrv4 I__2804 (
            .O(N__14840),
            .I(measured_delay_hc_16));
    InMux I__2803 (
            .O(N__14831),
            .I(N__14825));
    InMux I__2802 (
            .O(N__14830),
            .I(N__14821));
    InMux I__2801 (
            .O(N__14829),
            .I(N__14818));
    InMux I__2800 (
            .O(N__14828),
            .I(N__14815));
    LocalMux I__2799 (
            .O(N__14825),
            .I(N__14811));
    InMux I__2798 (
            .O(N__14824),
            .I(N__14808));
    LocalMux I__2797 (
            .O(N__14821),
            .I(N__14803));
    LocalMux I__2796 (
            .O(N__14818),
            .I(N__14803));
    LocalMux I__2795 (
            .O(N__14815),
            .I(N__14800));
    InMux I__2794 (
            .O(N__14814),
            .I(N__14797));
    Span4Mux_h I__2793 (
            .O(N__14811),
            .I(N__14794));
    LocalMux I__2792 (
            .O(N__14808),
            .I(N__14789));
    Span4Mux_h I__2791 (
            .O(N__14803),
            .I(N__14789));
    Span4Mux_h I__2790 (
            .O(N__14800),
            .I(N__14786));
    LocalMux I__2789 (
            .O(N__14797),
            .I(measured_delay_hc_14));
    Odrv4 I__2788 (
            .O(N__14794),
            .I(measured_delay_hc_14));
    Odrv4 I__2787 (
            .O(N__14789),
            .I(measured_delay_hc_14));
    Odrv4 I__2786 (
            .O(N__14786),
            .I(measured_delay_hc_14));
    CascadeMux I__2785 (
            .O(N__14777),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_ ));
    InMux I__2784 (
            .O(N__14774),
            .I(N__14771));
    LocalMux I__2783 (
            .O(N__14771),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ));
    InMux I__2782 (
            .O(N__14768),
            .I(N__14765));
    LocalMux I__2781 (
            .O(N__14765),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2 ));
    CascadeMux I__2780 (
            .O(N__14762),
            .I(N__14759));
    InMux I__2779 (
            .O(N__14759),
            .I(N__14756));
    LocalMux I__2778 (
            .O(N__14756),
            .I(N__14753));
    Odrv4 I__2777 (
            .O(N__14753),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_0_1 ));
    InMux I__2776 (
            .O(N__14750),
            .I(N__14747));
    LocalMux I__2775 (
            .O(N__14747),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ));
    CascadeMux I__2774 (
            .O(N__14744),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8_cascade_ ));
    InMux I__2773 (
            .O(N__14741),
            .I(N__14738));
    LocalMux I__2772 (
            .O(N__14738),
            .I(N__14735));
    Odrv4 I__2771 (
            .O(N__14735),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1 ));
    InMux I__2770 (
            .O(N__14732),
            .I(N__14726));
    InMux I__2769 (
            .O(N__14731),
            .I(N__14723));
    CascadeMux I__2768 (
            .O(N__14730),
            .I(N__14719));
    CascadeMux I__2767 (
            .O(N__14729),
            .I(N__14716));
    LocalMux I__2766 (
            .O(N__14726),
            .I(N__14711));
    LocalMux I__2765 (
            .O(N__14723),
            .I(N__14711));
    InMux I__2764 (
            .O(N__14722),
            .I(N__14708));
    InMux I__2763 (
            .O(N__14719),
            .I(N__14705));
    InMux I__2762 (
            .O(N__14716),
            .I(N__14702));
    Span4Mux_h I__2761 (
            .O(N__14711),
            .I(N__14699));
    LocalMux I__2760 (
            .O(N__14708),
            .I(N__14696));
    LocalMux I__2759 (
            .O(N__14705),
            .I(N__14693));
    LocalMux I__2758 (
            .O(N__14702),
            .I(measured_delay_hc_5));
    Odrv4 I__2757 (
            .O(N__14699),
            .I(measured_delay_hc_5));
    Odrv4 I__2756 (
            .O(N__14696),
            .I(measured_delay_hc_5));
    Odrv4 I__2755 (
            .O(N__14693),
            .I(measured_delay_hc_5));
    InMux I__2754 (
            .O(N__14684),
            .I(N__14677));
    InMux I__2753 (
            .O(N__14683),
            .I(N__14677));
    InMux I__2752 (
            .O(N__14682),
            .I(N__14674));
    LocalMux I__2751 (
            .O(N__14677),
            .I(N__14671));
    LocalMux I__2750 (
            .O(N__14674),
            .I(measured_delay_hc_20));
    Odrv4 I__2749 (
            .O(N__14671),
            .I(measured_delay_hc_20));
    CascadeMux I__2748 (
            .O(N__14666),
            .I(N__14662));
    InMux I__2747 (
            .O(N__14665),
            .I(N__14659));
    InMux I__2746 (
            .O(N__14662),
            .I(N__14656));
    LocalMux I__2745 (
            .O(N__14659),
            .I(N__14653));
    LocalMux I__2744 (
            .O(N__14656),
            .I(N__14647));
    Span4Mux_h I__2743 (
            .O(N__14653),
            .I(N__14644));
    InMux I__2742 (
            .O(N__14652),
            .I(N__14641));
    InMux I__2741 (
            .O(N__14651),
            .I(N__14638));
    InMux I__2740 (
            .O(N__14650),
            .I(N__14635));
    Span4Mux_v I__2739 (
            .O(N__14647),
            .I(N__14632));
    Span4Mux_v I__2738 (
            .O(N__14644),
            .I(N__14625));
    LocalMux I__2737 (
            .O(N__14641),
            .I(N__14625));
    LocalMux I__2736 (
            .O(N__14638),
            .I(N__14625));
    LocalMux I__2735 (
            .O(N__14635),
            .I(measured_delay_hc_3));
    Odrv4 I__2734 (
            .O(N__14632),
            .I(measured_delay_hc_3));
    Odrv4 I__2733 (
            .O(N__14625),
            .I(measured_delay_hc_3));
    CascadeMux I__2732 (
            .O(N__14618),
            .I(N__14611));
    InMux I__2731 (
            .O(N__14617),
            .I(N__14608));
    InMux I__2730 (
            .O(N__14616),
            .I(N__14605));
    InMux I__2729 (
            .O(N__14615),
            .I(N__14602));
    InMux I__2728 (
            .O(N__14614),
            .I(N__14599));
    InMux I__2727 (
            .O(N__14611),
            .I(N__14596));
    LocalMux I__2726 (
            .O(N__14608),
            .I(N__14593));
    LocalMux I__2725 (
            .O(N__14605),
            .I(N__14588));
    LocalMux I__2724 (
            .O(N__14602),
            .I(N__14588));
    LocalMux I__2723 (
            .O(N__14599),
            .I(N__14585));
    LocalMux I__2722 (
            .O(N__14596),
            .I(N__14580));
    Span4Mux_v I__2721 (
            .O(N__14593),
            .I(N__14580));
    Span4Mux_h I__2720 (
            .O(N__14588),
            .I(N__14577));
    Odrv4 I__2719 (
            .O(N__14585),
            .I(measured_delay_hc_17));
    Odrv4 I__2718 (
            .O(N__14580),
            .I(measured_delay_hc_17));
    Odrv4 I__2717 (
            .O(N__14577),
            .I(measured_delay_hc_17));
    CascadeMux I__2716 (
            .O(N__14570),
            .I(N__14566));
    InMux I__2715 (
            .O(N__14569),
            .I(N__14562));
    InMux I__2714 (
            .O(N__14566),
            .I(N__14559));
    InMux I__2713 (
            .O(N__14565),
            .I(N__14555));
    LocalMux I__2712 (
            .O(N__14562),
            .I(N__14551));
    LocalMux I__2711 (
            .O(N__14559),
            .I(N__14548));
    CascadeMux I__2710 (
            .O(N__14558),
            .I(N__14545));
    LocalMux I__2709 (
            .O(N__14555),
            .I(N__14542));
    InMux I__2708 (
            .O(N__14554),
            .I(N__14539));
    Span4Mux_v I__2707 (
            .O(N__14551),
            .I(N__14536));
    Span4Mux_v I__2706 (
            .O(N__14548),
            .I(N__14533));
    InMux I__2705 (
            .O(N__14545),
            .I(N__14530));
    Span4Mux_v I__2704 (
            .O(N__14542),
            .I(N__14525));
    LocalMux I__2703 (
            .O(N__14539),
            .I(N__14525));
    Span4Mux_v I__2702 (
            .O(N__14536),
            .I(N__14520));
    Span4Mux_h I__2701 (
            .O(N__14533),
            .I(N__14520));
    LocalMux I__2700 (
            .O(N__14530),
            .I(N__14515));
    Span4Mux_v I__2699 (
            .O(N__14525),
            .I(N__14515));
    Odrv4 I__2698 (
            .O(N__14520),
            .I(measured_delay_hc_6));
    Odrv4 I__2697 (
            .O(N__14515),
            .I(measured_delay_hc_6));
    InMux I__2696 (
            .O(N__14510),
            .I(N__14504));
    InMux I__2695 (
            .O(N__14509),
            .I(N__14501));
    CascadeMux I__2694 (
            .O(N__14508),
            .I(N__14498));
    InMux I__2693 (
            .O(N__14507),
            .I(N__14494));
    LocalMux I__2692 (
            .O(N__14504),
            .I(N__14489));
    LocalMux I__2691 (
            .O(N__14501),
            .I(N__14489));
    InMux I__2690 (
            .O(N__14498),
            .I(N__14486));
    CascadeMux I__2689 (
            .O(N__14497),
            .I(N__14483));
    LocalMux I__2688 (
            .O(N__14494),
            .I(N__14480));
    Span4Mux_h I__2687 (
            .O(N__14489),
            .I(N__14475));
    LocalMux I__2686 (
            .O(N__14486),
            .I(N__14475));
    InMux I__2685 (
            .O(N__14483),
            .I(N__14472));
    Span4Mux_h I__2684 (
            .O(N__14480),
            .I(N__14469));
    Span4Mux_v I__2683 (
            .O(N__14475),
            .I(N__14466));
    LocalMux I__2682 (
            .O(N__14472),
            .I(measured_delay_hc_13));
    Odrv4 I__2681 (
            .O(N__14469),
            .I(measured_delay_hc_13));
    Odrv4 I__2680 (
            .O(N__14466),
            .I(measured_delay_hc_13));
    CascadeMux I__2679 (
            .O(N__14459),
            .I(N__14454));
    CascadeMux I__2678 (
            .O(N__14458),
            .I(N__14451));
    InMux I__2677 (
            .O(N__14457),
            .I(N__14446));
    InMux I__2676 (
            .O(N__14454),
            .I(N__14443));
    InMux I__2675 (
            .O(N__14451),
            .I(N__14440));
    CascadeMux I__2674 (
            .O(N__14450),
            .I(N__14437));
    InMux I__2673 (
            .O(N__14449),
            .I(N__14434));
    LocalMux I__2672 (
            .O(N__14446),
            .I(N__14431));
    LocalMux I__2671 (
            .O(N__14443),
            .I(N__14428));
    LocalMux I__2670 (
            .O(N__14440),
            .I(N__14425));
    InMux I__2669 (
            .O(N__14437),
            .I(N__14422));
    LocalMux I__2668 (
            .O(N__14434),
            .I(N__14419));
    Span4Mux_v I__2667 (
            .O(N__14431),
            .I(N__14416));
    Span4Mux_h I__2666 (
            .O(N__14428),
            .I(N__14413));
    Span4Mux_v I__2665 (
            .O(N__14425),
            .I(N__14410));
    LocalMux I__2664 (
            .O(N__14422),
            .I(measured_delay_hc_19));
    Odrv4 I__2663 (
            .O(N__14419),
            .I(measured_delay_hc_19));
    Odrv4 I__2662 (
            .O(N__14416),
            .I(measured_delay_hc_19));
    Odrv4 I__2661 (
            .O(N__14413),
            .I(measured_delay_hc_19));
    Odrv4 I__2660 (
            .O(N__14410),
            .I(measured_delay_hc_19));
    InMux I__2659 (
            .O(N__14399),
            .I(N__14394));
    InMux I__2658 (
            .O(N__14398),
            .I(N__14389));
    CascadeMux I__2657 (
            .O(N__14397),
            .I(N__14386));
    LocalMux I__2656 (
            .O(N__14394),
            .I(N__14382));
    InMux I__2655 (
            .O(N__14393),
            .I(N__14379));
    InMux I__2654 (
            .O(N__14392),
            .I(N__14376));
    LocalMux I__2653 (
            .O(N__14389),
            .I(N__14373));
    InMux I__2652 (
            .O(N__14386),
            .I(N__14370));
    CascadeMux I__2651 (
            .O(N__14385),
            .I(N__14367));
    Span4Mux_h I__2650 (
            .O(N__14382),
            .I(N__14360));
    LocalMux I__2649 (
            .O(N__14379),
            .I(N__14360));
    LocalMux I__2648 (
            .O(N__14376),
            .I(N__14360));
    Span4Mux_v I__2647 (
            .O(N__14373),
            .I(N__14355));
    LocalMux I__2646 (
            .O(N__14370),
            .I(N__14355));
    InMux I__2645 (
            .O(N__14367),
            .I(N__14352));
    Span4Mux_v I__2644 (
            .O(N__14360),
            .I(N__14349));
    Span4Mux_h I__2643 (
            .O(N__14355),
            .I(N__14346));
    LocalMux I__2642 (
            .O(N__14352),
            .I(measured_delay_hc_15));
    Odrv4 I__2641 (
            .O(N__14349),
            .I(measured_delay_hc_15));
    Odrv4 I__2640 (
            .O(N__14346),
            .I(measured_delay_hc_15));
    InMux I__2639 (
            .O(N__14339),
            .I(N__14334));
    InMux I__2638 (
            .O(N__14338),
            .I(N__14329));
    InMux I__2637 (
            .O(N__14337),
            .I(N__14326));
    LocalMux I__2636 (
            .O(N__14334),
            .I(N__14323));
    InMux I__2635 (
            .O(N__14333),
            .I(N__14320));
    CascadeMux I__2634 (
            .O(N__14332),
            .I(N__14317));
    LocalMux I__2633 (
            .O(N__14329),
            .I(N__14308));
    LocalMux I__2632 (
            .O(N__14326),
            .I(N__14308));
    Span4Mux_v I__2631 (
            .O(N__14323),
            .I(N__14308));
    LocalMux I__2630 (
            .O(N__14320),
            .I(N__14308));
    InMux I__2629 (
            .O(N__14317),
            .I(N__14305));
    Span4Mux_h I__2628 (
            .O(N__14308),
            .I(N__14302));
    LocalMux I__2627 (
            .O(N__14305),
            .I(measured_delay_hc_18));
    Odrv4 I__2626 (
            .O(N__14302),
            .I(measured_delay_hc_18));
    InMux I__2625 (
            .O(N__14297),
            .I(N__14294));
    LocalMux I__2624 (
            .O(N__14294),
            .I(N__14291));
    Odrv4 I__2623 (
            .O(N__14291),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    InMux I__2622 (
            .O(N__14288),
            .I(N__14285));
    LocalMux I__2621 (
            .O(N__14285),
            .I(N__14282));
    Odrv4 I__2620 (
            .O(N__14282),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    InMux I__2619 (
            .O(N__14279),
            .I(N__14276));
    LocalMux I__2618 (
            .O(N__14276),
            .I(N__14273));
    Odrv4 I__2617 (
            .O(N__14273),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__2616 (
            .O(N__14270),
            .I(N__14267));
    LocalMux I__2615 (
            .O(N__14267),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    InMux I__2614 (
            .O(N__14264),
            .I(N__14259));
    InMux I__2613 (
            .O(N__14263),
            .I(N__14256));
    InMux I__2612 (
            .O(N__14262),
            .I(N__14253));
    LocalMux I__2611 (
            .O(N__14259),
            .I(N__14246));
    LocalMux I__2610 (
            .O(N__14256),
            .I(N__14246));
    LocalMux I__2609 (
            .O(N__14253),
            .I(N__14243));
    InMux I__2608 (
            .O(N__14252),
            .I(N__14240));
    InMux I__2607 (
            .O(N__14251),
            .I(N__14237));
    Span4Mux_h I__2606 (
            .O(N__14246),
            .I(N__14234));
    Span4Mux_h I__2605 (
            .O(N__14243),
            .I(N__14229));
    LocalMux I__2604 (
            .O(N__14240),
            .I(N__14229));
    LocalMux I__2603 (
            .O(N__14237),
            .I(measured_delay_hc_4));
    Odrv4 I__2602 (
            .O(N__14234),
            .I(measured_delay_hc_4));
    Odrv4 I__2601 (
            .O(N__14229),
            .I(measured_delay_hc_4));
    CascadeMux I__2600 (
            .O(N__14222),
            .I(N__14218));
    CascadeMux I__2599 (
            .O(N__14221),
            .I(N__14215));
    InMux I__2598 (
            .O(N__14218),
            .I(N__14211));
    InMux I__2597 (
            .O(N__14215),
            .I(N__14208));
    CascadeMux I__2596 (
            .O(N__14214),
            .I(N__14203));
    LocalMux I__2595 (
            .O(N__14211),
            .I(N__14200));
    LocalMux I__2594 (
            .O(N__14208),
            .I(N__14197));
    InMux I__2593 (
            .O(N__14207),
            .I(N__14192));
    InMux I__2592 (
            .O(N__14206),
            .I(N__14192));
    InMux I__2591 (
            .O(N__14203),
            .I(N__14189));
    Span4Mux_h I__2590 (
            .O(N__14200),
            .I(N__14186));
    Span4Mux_v I__2589 (
            .O(N__14197),
            .I(N__14183));
    LocalMux I__2588 (
            .O(N__14192),
            .I(N__14180));
    LocalMux I__2587 (
            .O(N__14189),
            .I(measured_delay_hc_1));
    Odrv4 I__2586 (
            .O(N__14186),
            .I(measured_delay_hc_1));
    Odrv4 I__2585 (
            .O(N__14183),
            .I(measured_delay_hc_1));
    Odrv4 I__2584 (
            .O(N__14180),
            .I(measured_delay_hc_1));
    InMux I__2583 (
            .O(N__14171),
            .I(N__14164));
    InMux I__2582 (
            .O(N__14170),
            .I(N__14164));
    InMux I__2581 (
            .O(N__14169),
            .I(N__14161));
    LocalMux I__2580 (
            .O(N__14164),
            .I(N__14158));
    LocalMux I__2579 (
            .O(N__14161),
            .I(N__14153));
    Span4Mux_h I__2578 (
            .O(N__14158),
            .I(N__14153));
    Odrv4 I__2577 (
            .O(N__14153),
            .I(measured_delay_hc_22));
    InMux I__2576 (
            .O(N__14150),
            .I(N__14143));
    InMux I__2575 (
            .O(N__14149),
            .I(N__14143));
    InMux I__2574 (
            .O(N__14148),
            .I(N__14140));
    LocalMux I__2573 (
            .O(N__14143),
            .I(N__14137));
    LocalMux I__2572 (
            .O(N__14140),
            .I(N__14132));
    Span4Mux_h I__2571 (
            .O(N__14137),
            .I(N__14132));
    Odrv4 I__2570 (
            .O(N__14132),
            .I(measured_delay_hc_21));
    CascadeMux I__2569 (
            .O(N__14129),
            .I(N__14126));
    InMux I__2568 (
            .O(N__14126),
            .I(N__14123));
    LocalMux I__2567 (
            .O(N__14123),
            .I(N__14117));
    InMux I__2566 (
            .O(N__14122),
            .I(N__14114));
    InMux I__2565 (
            .O(N__14121),
            .I(N__14111));
    InMux I__2564 (
            .O(N__14120),
            .I(N__14108));
    Span4Mux_h I__2563 (
            .O(N__14117),
            .I(N__14105));
    LocalMux I__2562 (
            .O(N__14114),
            .I(N__14102));
    LocalMux I__2561 (
            .O(N__14111),
            .I(N__14099));
    LocalMux I__2560 (
            .O(N__14108),
            .I(measured_delay_hc_0));
    Odrv4 I__2559 (
            .O(N__14105),
            .I(measured_delay_hc_0));
    Odrv12 I__2558 (
            .O(N__14102),
            .I(measured_delay_hc_0));
    Odrv4 I__2557 (
            .O(N__14099),
            .I(measured_delay_hc_0));
    CascadeMux I__2556 (
            .O(N__14090),
            .I(N__14087));
    InMux I__2555 (
            .O(N__14087),
            .I(N__14084));
    LocalMux I__2554 (
            .O(N__14084),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ));
    CascadeMux I__2553 (
            .O(N__14081),
            .I(N__14078));
    InMux I__2552 (
            .O(N__14078),
            .I(N__14075));
    LocalMux I__2551 (
            .O(N__14075),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ));
    CascadeMux I__2550 (
            .O(N__14072),
            .I(N__14069));
    InMux I__2549 (
            .O(N__14069),
            .I(N__14066));
    LocalMux I__2548 (
            .O(N__14066),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ));
    CascadeMux I__2547 (
            .O(N__14063),
            .I(N__14060));
    InMux I__2546 (
            .O(N__14060),
            .I(N__14057));
    LocalMux I__2545 (
            .O(N__14057),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ));
    InMux I__2544 (
            .O(N__14054),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__2543 (
            .O(N__14051),
            .I(\phase_controller_inst1.stoper_hc.time_passed11_cascade_ ));
    InMux I__2542 (
            .O(N__14048),
            .I(N__14045));
    LocalMux I__2541 (
            .O(N__14045),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__2540 (
            .O(N__14042),
            .I(N__14039));
    InMux I__2539 (
            .O(N__14039),
            .I(N__14036));
    LocalMux I__2538 (
            .O(N__14036),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__2537 (
            .O(N__14033),
            .I(N__14030));
    InMux I__2536 (
            .O(N__14030),
            .I(N__14027));
    LocalMux I__2535 (
            .O(N__14027),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__2534 (
            .O(N__14024),
            .I(N__14021));
    InMux I__2533 (
            .O(N__14021),
            .I(N__14018));
    LocalMux I__2532 (
            .O(N__14018),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__2531 (
            .O(N__14015),
            .I(N__14012));
    InMux I__2530 (
            .O(N__14012),
            .I(N__14009));
    LocalMux I__2529 (
            .O(N__14009),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__2528 (
            .O(N__14006),
            .I(N__14003));
    InMux I__2527 (
            .O(N__14003),
            .I(N__14000));
    LocalMux I__2526 (
            .O(N__14000),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__2525 (
            .O(N__13997),
            .I(N__13994));
    LocalMux I__2524 (
            .O(N__13994),
            .I(N__13991));
    Odrv4 I__2523 (
            .O(N__13991),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    CascadeMux I__2522 (
            .O(N__13988),
            .I(N__13985));
    InMux I__2521 (
            .O(N__13985),
            .I(N__13982));
    LocalMux I__2520 (
            .O(N__13982),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__2519 (
            .O(N__13979),
            .I(N__13976));
    InMux I__2518 (
            .O(N__13976),
            .I(N__13973));
    LocalMux I__2517 (
            .O(N__13973),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__2516 (
            .O(N__13970),
            .I(N__13967));
    LocalMux I__2515 (
            .O(N__13967),
            .I(N__13964));
    Span4Mux_h I__2514 (
            .O(N__13964),
            .I(N__13961));
    Odrv4 I__2513 (
            .O(N__13961),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__2512 (
            .O(N__13958),
            .I(N__13955));
    InMux I__2511 (
            .O(N__13955),
            .I(N__13952));
    LocalMux I__2510 (
            .O(N__13952),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    CascadeMux I__2509 (
            .O(N__13949),
            .I(N__13946));
    InMux I__2508 (
            .O(N__13946),
            .I(N__13943));
    LocalMux I__2507 (
            .O(N__13943),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ));
    InMux I__2506 (
            .O(N__13940),
            .I(N__13937));
    LocalMux I__2505 (
            .O(N__13937),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__2504 (
            .O(N__13934),
            .I(N__13931));
    InMux I__2503 (
            .O(N__13931),
            .I(N__13928));
    LocalMux I__2502 (
            .O(N__13928),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__2501 (
            .O(N__13925),
            .I(N__13922));
    LocalMux I__2500 (
            .O(N__13922),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__2499 (
            .O(N__13919),
            .I(N__13916));
    InMux I__2498 (
            .O(N__13916),
            .I(N__13913));
    LocalMux I__2497 (
            .O(N__13913),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__2496 (
            .O(N__13910),
            .I(N__13907));
    LocalMux I__2495 (
            .O(N__13907),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__2494 (
            .O(N__13904),
            .I(N__13901));
    InMux I__2493 (
            .O(N__13901),
            .I(N__13898));
    LocalMux I__2492 (
            .O(N__13898),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__2491 (
            .O(N__13895),
            .I(N__13892));
    LocalMux I__2490 (
            .O(N__13892),
            .I(N__13889));
    Odrv4 I__2489 (
            .O(N__13889),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__2488 (
            .O(N__13886),
            .I(N__13883));
    InMux I__2487 (
            .O(N__13883),
            .I(N__13880));
    LocalMux I__2486 (
            .O(N__13880),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__2485 (
            .O(N__13877),
            .I(N__13874));
    LocalMux I__2484 (
            .O(N__13874),
            .I(N__13871));
    Odrv4 I__2483 (
            .O(N__13871),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__2482 (
            .O(N__13868),
            .I(N__13865));
    InMux I__2481 (
            .O(N__13865),
            .I(N__13862));
    LocalMux I__2480 (
            .O(N__13862),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__2479 (
            .O(N__13859),
            .I(N__13856));
    LocalMux I__2478 (
            .O(N__13856),
            .I(N__13853));
    Odrv4 I__2477 (
            .O(N__13853),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ));
    CascadeMux I__2476 (
            .O(N__13850),
            .I(N__13847));
    InMux I__2475 (
            .O(N__13847),
            .I(N__13844));
    LocalMux I__2474 (
            .O(N__13844),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__2473 (
            .O(N__13841),
            .I(N__13838));
    LocalMux I__2472 (
            .O(N__13838),
            .I(N__13835));
    Odrv4 I__2471 (
            .O(N__13835),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    CascadeMux I__2470 (
            .O(N__13832),
            .I(N__13829));
    InMux I__2469 (
            .O(N__13829),
            .I(N__13826));
    LocalMux I__2468 (
            .O(N__13826),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    CEMux I__2467 (
            .O(N__13823),
            .I(N__13819));
    CEMux I__2466 (
            .O(N__13822),
            .I(N__13816));
    LocalMux I__2465 (
            .O(N__13819),
            .I(N__13813));
    LocalMux I__2464 (
            .O(N__13816),
            .I(N__13809));
    Span4Mux_v I__2463 (
            .O(N__13813),
            .I(N__13806));
    CEMux I__2462 (
            .O(N__13812),
            .I(N__13803));
    Span4Mux_h I__2461 (
            .O(N__13809),
            .I(N__13800));
    Span4Mux_s2_h I__2460 (
            .O(N__13806),
            .I(N__13795));
    LocalMux I__2459 (
            .O(N__13803),
            .I(N__13795));
    Span4Mux_h I__2458 (
            .O(N__13800),
            .I(N__13792));
    Sp12to4 I__2457 (
            .O(N__13795),
            .I(N__13789));
    Odrv4 I__2456 (
            .O(N__13792),
            .I(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv12 I__2455 (
            .O(N__13789),
            .I(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ));
    CascadeMux I__2454 (
            .O(N__13784),
            .I(N__13779));
    InMux I__2453 (
            .O(N__13783),
            .I(N__13776));
    InMux I__2452 (
            .O(N__13782),
            .I(N__13773));
    InMux I__2451 (
            .O(N__13779),
            .I(N__13770));
    LocalMux I__2450 (
            .O(N__13776),
            .I(N__13766));
    LocalMux I__2449 (
            .O(N__13773),
            .I(N__13763));
    LocalMux I__2448 (
            .O(N__13770),
            .I(N__13760));
    CascadeMux I__2447 (
            .O(N__13769),
            .I(N__13757));
    Span4Mux_h I__2446 (
            .O(N__13766),
            .I(N__13754));
    Span4Mux_h I__2445 (
            .O(N__13763),
            .I(N__13749));
    Span4Mux_h I__2444 (
            .O(N__13760),
            .I(N__13749));
    InMux I__2443 (
            .O(N__13757),
            .I(N__13746));
    Odrv4 I__2442 (
            .O(N__13754),
            .I(measured_delay_tr_19));
    Odrv4 I__2441 (
            .O(N__13749),
            .I(measured_delay_tr_19));
    LocalMux I__2440 (
            .O(N__13746),
            .I(measured_delay_tr_19));
    InMux I__2439 (
            .O(N__13739),
            .I(N__13736));
    LocalMux I__2438 (
            .O(N__13736),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__2437 (
            .O(N__13733),
            .I(N__13729));
    InMux I__2436 (
            .O(N__13732),
            .I(N__13726));
    LocalMux I__2435 (
            .O(N__13729),
            .I(N__13723));
    LocalMux I__2434 (
            .O(N__13726),
            .I(N__13720));
    Span4Mux_h I__2433 (
            .O(N__13723),
            .I(N__13715));
    Span4Mux_h I__2432 (
            .O(N__13720),
            .I(N__13712));
    InMux I__2431 (
            .O(N__13719),
            .I(N__13709));
    InMux I__2430 (
            .O(N__13718),
            .I(N__13706));
    Odrv4 I__2429 (
            .O(N__13715),
            .I(measured_delay_tr_17));
    Odrv4 I__2428 (
            .O(N__13712),
            .I(measured_delay_tr_17));
    LocalMux I__2427 (
            .O(N__13709),
            .I(measured_delay_tr_17));
    LocalMux I__2426 (
            .O(N__13706),
            .I(measured_delay_tr_17));
    InMux I__2425 (
            .O(N__13697),
            .I(N__13694));
    LocalMux I__2424 (
            .O(N__13694),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__2423 (
            .O(N__13691),
            .I(N__13687));
    InMux I__2422 (
            .O(N__13690),
            .I(N__13684));
    LocalMux I__2421 (
            .O(N__13687),
            .I(N__13681));
    LocalMux I__2420 (
            .O(N__13684),
            .I(N__13678));
    Span4Mux_v I__2419 (
            .O(N__13681),
            .I(N__13671));
    Span4Mux_v I__2418 (
            .O(N__13678),
            .I(N__13671));
    InMux I__2417 (
            .O(N__13677),
            .I(N__13668));
    InMux I__2416 (
            .O(N__13676),
            .I(N__13665));
    Odrv4 I__2415 (
            .O(N__13671),
            .I(measured_delay_tr_18));
    LocalMux I__2414 (
            .O(N__13668),
            .I(measured_delay_tr_18));
    LocalMux I__2413 (
            .O(N__13665),
            .I(measured_delay_tr_18));
    InMux I__2412 (
            .O(N__13658),
            .I(N__13655));
    LocalMux I__2411 (
            .O(N__13655),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    InMux I__2410 (
            .O(N__13652),
            .I(N__13649));
    LocalMux I__2409 (
            .O(N__13649),
            .I(N__13645));
    InMux I__2408 (
            .O(N__13648),
            .I(N__13641));
    Span4Mux_h I__2407 (
            .O(N__13645),
            .I(N__13637));
    InMux I__2406 (
            .O(N__13644),
            .I(N__13634));
    LocalMux I__2405 (
            .O(N__13641),
            .I(N__13631));
    InMux I__2404 (
            .O(N__13640),
            .I(N__13628));
    Span4Mux_v I__2403 (
            .O(N__13637),
            .I(N__13623));
    LocalMux I__2402 (
            .O(N__13634),
            .I(N__13623));
    Odrv4 I__2401 (
            .O(N__13631),
            .I(measured_delay_tr_16));
    LocalMux I__2400 (
            .O(N__13628),
            .I(measured_delay_tr_16));
    Odrv4 I__2399 (
            .O(N__13623),
            .I(measured_delay_tr_16));
    InMux I__2398 (
            .O(N__13616),
            .I(N__13613));
    LocalMux I__2397 (
            .O(N__13613),
            .I(N__13610));
    Odrv12 I__2396 (
            .O(N__13610),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__2395 (
            .O(N__13607),
            .I(N__13595));
    InMux I__2394 (
            .O(N__13606),
            .I(N__13595));
    InMux I__2393 (
            .O(N__13605),
            .I(N__13595));
    InMux I__2392 (
            .O(N__13604),
            .I(N__13595));
    LocalMux I__2391 (
            .O(N__13595),
            .I(N__13592));
    Span4Mux_h I__2390 (
            .O(N__13592),
            .I(N__13585));
    InMux I__2389 (
            .O(N__13591),
            .I(N__13576));
    InMux I__2388 (
            .O(N__13590),
            .I(N__13576));
    InMux I__2387 (
            .O(N__13589),
            .I(N__13576));
    InMux I__2386 (
            .O(N__13588),
            .I(N__13576));
    Span4Mux_v I__2385 (
            .O(N__13585),
            .I(N__13573));
    LocalMux I__2384 (
            .O(N__13576),
            .I(N__13570));
    Odrv4 I__2383 (
            .O(N__13573),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    Odrv12 I__2382 (
            .O(N__13570),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    CascadeMux I__2381 (
            .O(N__13565),
            .I(N__13562));
    InMux I__2380 (
            .O(N__13562),
            .I(N__13559));
    LocalMux I__2379 (
            .O(N__13559),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    InMux I__2378 (
            .O(N__13556),
            .I(N__13553));
    LocalMux I__2377 (
            .O(N__13553),
            .I(N__13550));
    Odrv4 I__2376 (
            .O(N__13550),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__2375 (
            .O(N__13547),
            .I(N__13544));
    InMux I__2374 (
            .O(N__13544),
            .I(N__13541));
    LocalMux I__2373 (
            .O(N__13541),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__2372 (
            .O(N__13538),
            .I(N__13535));
    InMux I__2371 (
            .O(N__13535),
            .I(N__13532));
    LocalMux I__2370 (
            .O(N__13532),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__2369 (
            .O(N__13529),
            .I(N__13526));
    InMux I__2368 (
            .O(N__13526),
            .I(N__13523));
    LocalMux I__2367 (
            .O(N__13523),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ));
    CascadeMux I__2366 (
            .O(N__13520),
            .I(N__13517));
    InMux I__2365 (
            .O(N__13517),
            .I(N__13514));
    LocalMux I__2364 (
            .O(N__13514),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ));
    CascadeMux I__2363 (
            .O(N__13511),
            .I(N__13508));
    InMux I__2362 (
            .O(N__13508),
            .I(N__13505));
    LocalMux I__2361 (
            .O(N__13505),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ));
    CascadeMux I__2360 (
            .O(N__13502),
            .I(N__13499));
    InMux I__2359 (
            .O(N__13499),
            .I(N__13496));
    LocalMux I__2358 (
            .O(N__13496),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ));
    InMux I__2357 (
            .O(N__13493),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__2356 (
            .O(N__13490),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_ ));
    InMux I__2355 (
            .O(N__13487),
            .I(N__13484));
    LocalMux I__2354 (
            .O(N__13484),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__2353 (
            .O(N__13481),
            .I(N__13478));
    InMux I__2352 (
            .O(N__13478),
            .I(N__13475));
    LocalMux I__2351 (
            .O(N__13475),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    InMux I__2350 (
            .O(N__13472),
            .I(N__13469));
    LocalMux I__2349 (
            .O(N__13469),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__2348 (
            .O(N__13466),
            .I(N__13463));
    InMux I__2347 (
            .O(N__13463),
            .I(N__13460));
    LocalMux I__2346 (
            .O(N__13460),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__2345 (
            .O(N__13457),
            .I(N__13454));
    LocalMux I__2344 (
            .O(N__13454),
            .I(N__13451));
    Odrv4 I__2343 (
            .O(N__13451),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__2342 (
            .O(N__13448),
            .I(N__13445));
    InMux I__2341 (
            .O(N__13445),
            .I(N__13442));
    LocalMux I__2340 (
            .O(N__13442),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__2339 (
            .O(N__13439),
            .I(N__13436));
    LocalMux I__2338 (
            .O(N__13436),
            .I(N__13433));
    Odrv4 I__2337 (
            .O(N__13433),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__2336 (
            .O(N__13430),
            .I(N__13427));
    InMux I__2335 (
            .O(N__13427),
            .I(N__13424));
    LocalMux I__2334 (
            .O(N__13424),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__2333 (
            .O(N__13421),
            .I(N__13418));
    LocalMux I__2332 (
            .O(N__13418),
            .I(N__13415));
    Odrv4 I__2331 (
            .O(N__13415),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__2330 (
            .O(N__13412),
            .I(N__13409));
    InMux I__2329 (
            .O(N__13409),
            .I(N__13406));
    LocalMux I__2328 (
            .O(N__13406),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__2327 (
            .O(N__13403),
            .I(N__13400));
    LocalMux I__2326 (
            .O(N__13400),
            .I(N__13397));
    Odrv4 I__2325 (
            .O(N__13397),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__2324 (
            .O(N__13394),
            .I(N__13391));
    InMux I__2323 (
            .O(N__13391),
            .I(N__13388));
    LocalMux I__2322 (
            .O(N__13388),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__2321 (
            .O(N__13385),
            .I(N__13382));
    LocalMux I__2320 (
            .O(N__13382),
            .I(N__13379));
    Odrv12 I__2319 (
            .O(N__13379),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__2318 (
            .O(N__13376),
            .I(N__13373));
    InMux I__2317 (
            .O(N__13373),
            .I(N__13370));
    LocalMux I__2316 (
            .O(N__13370),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__2315 (
            .O(N__13367),
            .I(N__13364));
    LocalMux I__2314 (
            .O(N__13364),
            .I(N__13361));
    Odrv4 I__2313 (
            .O(N__13361),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__2312 (
            .O(N__13358),
            .I(N__13355));
    LocalMux I__2311 (
            .O(N__13355),
            .I(N__13350));
    InMux I__2310 (
            .O(N__13354),
            .I(N__13347));
    InMux I__2309 (
            .O(N__13353),
            .I(N__13344));
    Odrv12 I__2308 (
            .O(N__13350),
            .I(measured_delay_tr_2));
    LocalMux I__2307 (
            .O(N__13347),
            .I(measured_delay_tr_2));
    LocalMux I__2306 (
            .O(N__13344),
            .I(measured_delay_tr_2));
    InMux I__2305 (
            .O(N__13337),
            .I(N__13331));
    InMux I__2304 (
            .O(N__13336),
            .I(N__13331));
    LocalMux I__2303 (
            .O(N__13331),
            .I(N__13328));
    Span4Mux_h I__2302 (
            .O(N__13328),
            .I(N__13322));
    InMux I__2301 (
            .O(N__13327),
            .I(N__13317));
    InMux I__2300 (
            .O(N__13326),
            .I(N__13317));
    InMux I__2299 (
            .O(N__13325),
            .I(N__13314));
    Odrv4 I__2298 (
            .O(N__13322),
            .I(measured_delay_tr_3));
    LocalMux I__2297 (
            .O(N__13317),
            .I(measured_delay_tr_3));
    LocalMux I__2296 (
            .O(N__13314),
            .I(measured_delay_tr_3));
    CascadeMux I__2295 (
            .O(N__13307),
            .I(N__13303));
    InMux I__2294 (
            .O(N__13306),
            .I(N__13294));
    InMux I__2293 (
            .O(N__13303),
            .I(N__13294));
    InMux I__2292 (
            .O(N__13302),
            .I(N__13294));
    CascadeMux I__2291 (
            .O(N__13301),
            .I(N__13290));
    LocalMux I__2290 (
            .O(N__13294),
            .I(N__13286));
    InMux I__2289 (
            .O(N__13293),
            .I(N__13279));
    InMux I__2288 (
            .O(N__13290),
            .I(N__13279));
    InMux I__2287 (
            .O(N__13289),
            .I(N__13279));
    Span4Mux_v I__2286 (
            .O(N__13286),
            .I(N__13276));
    LocalMux I__2285 (
            .O(N__13279),
            .I(N__13273));
    Odrv4 I__2284 (
            .O(N__13276),
            .I(\phase_controller_inst1.stoper_tr.N_109 ));
    Odrv4 I__2283 (
            .O(N__13273),
            .I(\phase_controller_inst1.stoper_tr.N_109 ));
    InMux I__2282 (
            .O(N__13268),
            .I(N__13256));
    InMux I__2281 (
            .O(N__13267),
            .I(N__13256));
    InMux I__2280 (
            .O(N__13266),
            .I(N__13256));
    InMux I__2279 (
            .O(N__13265),
            .I(N__13249));
    InMux I__2278 (
            .O(N__13264),
            .I(N__13249));
    InMux I__2277 (
            .O(N__13263),
            .I(N__13249));
    LocalMux I__2276 (
            .O(N__13256),
            .I(N__13246));
    LocalMux I__2275 (
            .O(N__13249),
            .I(N__13243));
    Span4Mux_h I__2274 (
            .O(N__13246),
            .I(N__13240));
    Odrv4 I__2273 (
            .O(N__13243),
            .I(\phase_controller_inst1.stoper_tr.N_110 ));
    Odrv4 I__2272 (
            .O(N__13240),
            .I(\phase_controller_inst1.stoper_tr.N_110 ));
    CascadeMux I__2271 (
            .O(N__13235),
            .I(N__13228));
    CascadeMux I__2270 (
            .O(N__13234),
            .I(N__13225));
    CascadeMux I__2269 (
            .O(N__13233),
            .I(N__13221));
    InMux I__2268 (
            .O(N__13232),
            .I(N__13218));
    InMux I__2267 (
            .O(N__13231),
            .I(N__13213));
    InMux I__2266 (
            .O(N__13228),
            .I(N__13213));
    InMux I__2265 (
            .O(N__13225),
            .I(N__13208));
    InMux I__2264 (
            .O(N__13224),
            .I(N__13208));
    InMux I__2263 (
            .O(N__13221),
            .I(N__13205));
    LocalMux I__2262 (
            .O(N__13218),
            .I(N__13200));
    LocalMux I__2261 (
            .O(N__13213),
            .I(N__13200));
    LocalMux I__2260 (
            .O(N__13208),
            .I(N__13195));
    LocalMux I__2259 (
            .O(N__13205),
            .I(N__13195));
    Span4Mux_h I__2258 (
            .O(N__13200),
            .I(N__13192));
    Odrv4 I__2257 (
            .O(N__13195),
            .I(\phase_controller_inst1.stoper_tr.N_92 ));
    Odrv4 I__2256 (
            .O(N__13192),
            .I(\phase_controller_inst1.stoper_tr.N_92 ));
    CascadeMux I__2255 (
            .O(N__13187),
            .I(N__13184));
    InMux I__2254 (
            .O(N__13184),
            .I(N__13180));
    CascadeMux I__2253 (
            .O(N__13183),
            .I(N__13176));
    LocalMux I__2252 (
            .O(N__13180),
            .I(N__13173));
    InMux I__2251 (
            .O(N__13179),
            .I(N__13170));
    InMux I__2250 (
            .O(N__13176),
            .I(N__13167));
    Span4Mux_h I__2249 (
            .O(N__13173),
            .I(N__13162));
    LocalMux I__2248 (
            .O(N__13170),
            .I(N__13162));
    LocalMux I__2247 (
            .O(N__13167),
            .I(measured_delay_tr_6));
    Odrv4 I__2246 (
            .O(N__13162),
            .I(measured_delay_tr_6));
    InMux I__2245 (
            .O(N__13157),
            .I(N__13146));
    InMux I__2244 (
            .O(N__13156),
            .I(N__13146));
    InMux I__2243 (
            .O(N__13155),
            .I(N__13146));
    InMux I__2242 (
            .O(N__13154),
            .I(N__13141));
    InMux I__2241 (
            .O(N__13153),
            .I(N__13141));
    LocalMux I__2240 (
            .O(N__13146),
            .I(N__13133));
    LocalMux I__2239 (
            .O(N__13141),
            .I(N__13130));
    InMux I__2238 (
            .O(N__13140),
            .I(N__13119));
    InMux I__2237 (
            .O(N__13139),
            .I(N__13119));
    InMux I__2236 (
            .O(N__13138),
            .I(N__13119));
    InMux I__2235 (
            .O(N__13137),
            .I(N__13119));
    InMux I__2234 (
            .O(N__13136),
            .I(N__13119));
    Span4Mux_h I__2233 (
            .O(N__13133),
            .I(N__13115));
    Span4Mux_v I__2232 (
            .O(N__13130),
            .I(N__13110));
    LocalMux I__2231 (
            .O(N__13119),
            .I(N__13110));
    InMux I__2230 (
            .O(N__13118),
            .I(N__13107));
    Odrv4 I__2229 (
            .O(N__13115),
            .I(\phase_controller_inst1.stoper_tr.N_95 ));
    Odrv4 I__2228 (
            .O(N__13110),
            .I(\phase_controller_inst1.stoper_tr.N_95 ));
    LocalMux I__2227 (
            .O(N__13107),
            .I(\phase_controller_inst1.stoper_tr.N_95 ));
    InMux I__2226 (
            .O(N__13100),
            .I(N__13097));
    LocalMux I__2225 (
            .O(N__13097),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__2224 (
            .O(N__13094),
            .I(N__13091));
    InMux I__2223 (
            .O(N__13091),
            .I(N__13088));
    LocalMux I__2222 (
            .O(N__13088),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__2221 (
            .O(N__13085),
            .I(N__13082));
    LocalMux I__2220 (
            .O(N__13082),
            .I(N__13079));
    Odrv4 I__2219 (
            .O(N__13079),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__2218 (
            .O(N__13076),
            .I(N__13073));
    InMux I__2217 (
            .O(N__13073),
            .I(N__13070));
    LocalMux I__2216 (
            .O(N__13070),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__2215 (
            .O(N__13067),
            .I(N__13064));
    LocalMux I__2214 (
            .O(N__13064),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__2213 (
            .O(N__13061),
            .I(N__13058));
    InMux I__2212 (
            .O(N__13058),
            .I(N__13055));
    LocalMux I__2211 (
            .O(N__13055),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__2210 (
            .O(N__13052),
            .I(N__13049));
    LocalMux I__2209 (
            .O(N__13049),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__2208 (
            .O(N__13046),
            .I(N__13043));
    InMux I__2207 (
            .O(N__13043),
            .I(N__13040));
    LocalMux I__2206 (
            .O(N__13040),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__2205 (
            .O(N__13037),
            .I(N__13034));
    LocalMux I__2204 (
            .O(N__13034),
            .I(N__13031));
    Odrv4 I__2203 (
            .O(N__13031),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__2202 (
            .O(N__13028),
            .I(N__13025));
    InMux I__2201 (
            .O(N__13025),
            .I(N__13022));
    LocalMux I__2200 (
            .O(N__13022),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__2199 (
            .O(N__13019),
            .I(N__13016));
    LocalMux I__2198 (
            .O(N__13016),
            .I(N__13012));
    InMux I__2197 (
            .O(N__13015),
            .I(N__13009));
    Span4Mux_v I__2196 (
            .O(N__13012),
            .I(N__13003));
    LocalMux I__2195 (
            .O(N__13009),
            .I(N__13003));
    InMux I__2194 (
            .O(N__13008),
            .I(N__13000));
    Odrv4 I__2193 (
            .O(N__13003),
            .I(measured_delay_tr_12));
    LocalMux I__2192 (
            .O(N__13000),
            .I(measured_delay_tr_12));
    InMux I__2191 (
            .O(N__12995),
            .I(N__12991));
    InMux I__2190 (
            .O(N__12994),
            .I(N__12988));
    LocalMux I__2189 (
            .O(N__12991),
            .I(N__12984));
    LocalMux I__2188 (
            .O(N__12988),
            .I(N__12981));
    CascadeMux I__2187 (
            .O(N__12987),
            .I(N__12978));
    Span4Mux_h I__2186 (
            .O(N__12984),
            .I(N__12975));
    Span4Mux_h I__2185 (
            .O(N__12981),
            .I(N__12972));
    InMux I__2184 (
            .O(N__12978),
            .I(N__12969));
    Odrv4 I__2183 (
            .O(N__12975),
            .I(measured_delay_tr_13));
    Odrv4 I__2182 (
            .O(N__12972),
            .I(measured_delay_tr_13));
    LocalMux I__2181 (
            .O(N__12969),
            .I(measured_delay_tr_13));
    InMux I__2180 (
            .O(N__12962),
            .I(N__12958));
    InMux I__2179 (
            .O(N__12961),
            .I(N__12953));
    LocalMux I__2178 (
            .O(N__12958),
            .I(N__12949));
    InMux I__2177 (
            .O(N__12957),
            .I(N__12944));
    InMux I__2176 (
            .O(N__12956),
            .I(N__12944));
    LocalMux I__2175 (
            .O(N__12953),
            .I(N__12941));
    InMux I__2174 (
            .O(N__12952),
            .I(N__12938));
    Span4Mux_v I__2173 (
            .O(N__12949),
            .I(N__12933));
    LocalMux I__2172 (
            .O(N__12944),
            .I(N__12933));
    Odrv4 I__2171 (
            .O(N__12941),
            .I(measured_delay_tr_14));
    LocalMux I__2170 (
            .O(N__12938),
            .I(measured_delay_tr_14));
    Odrv4 I__2169 (
            .O(N__12933),
            .I(measured_delay_tr_14));
    InMux I__2168 (
            .O(N__12926),
            .I(N__12911));
    InMux I__2167 (
            .O(N__12925),
            .I(N__12911));
    InMux I__2166 (
            .O(N__12924),
            .I(N__12911));
    InMux I__2165 (
            .O(N__12923),
            .I(N__12911));
    InMux I__2164 (
            .O(N__12922),
            .I(N__12911));
    LocalMux I__2163 (
            .O(N__12911),
            .I(N__12907));
    CascadeMux I__2162 (
            .O(N__12910),
            .I(N__12900));
    Span4Mux_v I__2161 (
            .O(N__12907),
            .I(N__12897));
    InMux I__2160 (
            .O(N__12906),
            .I(N__12886));
    InMux I__2159 (
            .O(N__12905),
            .I(N__12886));
    InMux I__2158 (
            .O(N__12904),
            .I(N__12886));
    InMux I__2157 (
            .O(N__12903),
            .I(N__12886));
    InMux I__2156 (
            .O(N__12900),
            .I(N__12886));
    Odrv4 I__2155 (
            .O(N__12897),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ));
    LocalMux I__2154 (
            .O(N__12886),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ));
    InMux I__2153 (
            .O(N__12881),
            .I(N__12877));
    InMux I__2152 (
            .O(N__12880),
            .I(N__12874));
    LocalMux I__2151 (
            .O(N__12877),
            .I(N__12870));
    LocalMux I__2150 (
            .O(N__12874),
            .I(N__12867));
    InMux I__2149 (
            .O(N__12873),
            .I(N__12864));
    Odrv4 I__2148 (
            .O(N__12870),
            .I(measured_delay_tr_10));
    Odrv4 I__2147 (
            .O(N__12867),
            .I(measured_delay_tr_10));
    LocalMux I__2146 (
            .O(N__12864),
            .I(measured_delay_tr_10));
    CascadeMux I__2145 (
            .O(N__12857),
            .I(N__12853));
    InMux I__2144 (
            .O(N__12856),
            .I(N__12850));
    InMux I__2143 (
            .O(N__12853),
            .I(N__12847));
    LocalMux I__2142 (
            .O(N__12850),
            .I(N__12844));
    LocalMux I__2141 (
            .O(N__12847),
            .I(N__12840));
    Span4Mux_h I__2140 (
            .O(N__12844),
            .I(N__12837));
    InMux I__2139 (
            .O(N__12843),
            .I(N__12834));
    Odrv12 I__2138 (
            .O(N__12840),
            .I(measured_delay_tr_4));
    Odrv4 I__2137 (
            .O(N__12837),
            .I(measured_delay_tr_4));
    LocalMux I__2136 (
            .O(N__12834),
            .I(measured_delay_tr_4));
    InMux I__2135 (
            .O(N__12827),
            .I(N__12824));
    LocalMux I__2134 (
            .O(N__12824),
            .I(N__12819));
    InMux I__2133 (
            .O(N__12823),
            .I(N__12812));
    InMux I__2132 (
            .O(N__12822),
            .I(N__12812));
    Span4Mux_v I__2131 (
            .O(N__12819),
            .I(N__12809));
    InMux I__2130 (
            .O(N__12818),
            .I(N__12806));
    CascadeMux I__2129 (
            .O(N__12817),
            .I(N__12803));
    LocalMux I__2128 (
            .O(N__12812),
            .I(N__12800));
    Span4Mux_h I__2127 (
            .O(N__12809),
            .I(N__12795));
    LocalMux I__2126 (
            .O(N__12806),
            .I(N__12795));
    InMux I__2125 (
            .O(N__12803),
            .I(N__12792));
    Span4Mux_v I__2124 (
            .O(N__12800),
            .I(N__12789));
    Odrv4 I__2123 (
            .O(N__12795),
            .I(measured_delay_tr_7));
    LocalMux I__2122 (
            .O(N__12792),
            .I(measured_delay_tr_7));
    Odrv4 I__2121 (
            .O(N__12789),
            .I(measured_delay_tr_7));
    InMux I__2120 (
            .O(N__12782),
            .I(N__12779));
    LocalMux I__2119 (
            .O(N__12779),
            .I(N__12773));
    InMux I__2118 (
            .O(N__12778),
            .I(N__12770));
    InMux I__2117 (
            .O(N__12777),
            .I(N__12767));
    CascadeMux I__2116 (
            .O(N__12776),
            .I(N__12764));
    Span4Mux_h I__2115 (
            .O(N__12773),
            .I(N__12759));
    LocalMux I__2114 (
            .O(N__12770),
            .I(N__12759));
    LocalMux I__2113 (
            .O(N__12767),
            .I(N__12756));
    InMux I__2112 (
            .O(N__12764),
            .I(N__12753));
    Span4Mux_h I__2111 (
            .O(N__12759),
            .I(N__12750));
    Odrv12 I__2110 (
            .O(N__12756),
            .I(measured_delay_tr_8));
    LocalMux I__2109 (
            .O(N__12753),
            .I(measured_delay_tr_8));
    Odrv4 I__2108 (
            .O(N__12750),
            .I(measured_delay_tr_8));
    InMux I__2107 (
            .O(N__12743),
            .I(N__12740));
    LocalMux I__2106 (
            .O(N__12740),
            .I(N__12735));
    InMux I__2105 (
            .O(N__12739),
            .I(N__12732));
    InMux I__2104 (
            .O(N__12738),
            .I(N__12729));
    Span4Mux_h I__2103 (
            .O(N__12735),
            .I(N__12724));
    LocalMux I__2102 (
            .O(N__12732),
            .I(N__12724));
    LocalMux I__2101 (
            .O(N__12729),
            .I(measured_delay_tr_5));
    Odrv4 I__2100 (
            .O(N__12724),
            .I(measured_delay_tr_5));
    InMux I__2099 (
            .O(N__12719),
            .I(N__12716));
    LocalMux I__2098 (
            .O(N__12716),
            .I(N__12713));
    Span4Mux_h I__2097 (
            .O(N__12713),
            .I(N__12709));
    InMux I__2096 (
            .O(N__12712),
            .I(N__12706));
    Odrv4 I__2095 (
            .O(N__12709),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ));
    LocalMux I__2094 (
            .O(N__12706),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ));
    CascadeMux I__2093 (
            .O(N__12701),
            .I(N__12697));
    CascadeMux I__2092 (
            .O(N__12700),
            .I(N__12694));
    InMux I__2091 (
            .O(N__12697),
            .I(N__12691));
    InMux I__2090 (
            .O(N__12694),
            .I(N__12688));
    LocalMux I__2089 (
            .O(N__12691),
            .I(N__12685));
    LocalMux I__2088 (
            .O(N__12688),
            .I(measured_delay_tr_1));
    Odrv12 I__2087 (
            .O(N__12685),
            .I(measured_delay_tr_1));
    CascadeMux I__2086 (
            .O(N__12680),
            .I(\phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_3_cascade_ ));
    InMux I__2085 (
            .O(N__12677),
            .I(N__12674));
    LocalMux I__2084 (
            .O(N__12674),
            .I(\phase_controller_inst1.stoper_hc.un1_m2_eZ0 ));
    CascadeMux I__2083 (
            .O(N__12671),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_ ));
    InMux I__2082 (
            .O(N__12668),
            .I(N__12665));
    LocalMux I__2081 (
            .O(N__12665),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11 ));
    CascadeMux I__2080 (
            .O(N__12662),
            .I(N__12659));
    InMux I__2079 (
            .O(N__12659),
            .I(N__12656));
    LocalMux I__2078 (
            .O(N__12656),
            .I(N__12652));
    InMux I__2077 (
            .O(N__12655),
            .I(N__12649));
    Odrv4 I__2076 (
            .O(N__12652),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_2_0Z0Z_0 ));
    LocalMux I__2075 (
            .O(N__12649),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_2_0Z0Z_0 ));
    InMux I__2074 (
            .O(N__12644),
            .I(N__12641));
    LocalMux I__2073 (
            .O(N__12641),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ));
    InMux I__2072 (
            .O(N__12638),
            .I(N__12635));
    LocalMux I__2071 (
            .O(N__12635),
            .I(N__12632));
    Glb2LocalMux I__2070 (
            .O(N__12632),
            .I(N__12629));
    GlobalMux I__2069 (
            .O(N__12629),
            .I(clk_12mhz));
    IoInMux I__2068 (
            .O(N__12626),
            .I(N__12623));
    LocalMux I__2067 (
            .O(N__12623),
            .I(N__12620));
    IoSpan4Mux I__2066 (
            .O(N__12620),
            .I(N__12617));
    Span4Mux_s0_v I__2065 (
            .O(N__12617),
            .I(N__12614));
    Odrv4 I__2064 (
            .O(N__12614),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__2063 (
            .O(N__12611),
            .I(N__12607));
    InMux I__2062 (
            .O(N__12610),
            .I(N__12604));
    LocalMux I__2061 (
            .O(N__12607),
            .I(N__12600));
    LocalMux I__2060 (
            .O(N__12604),
            .I(N__12597));
    InMux I__2059 (
            .O(N__12603),
            .I(N__12594));
    Odrv4 I__2058 (
            .O(N__12600),
            .I(measured_delay_tr_11));
    Odrv4 I__2057 (
            .O(N__12597),
            .I(measured_delay_tr_11));
    LocalMux I__2056 (
            .O(N__12594),
            .I(measured_delay_tr_11));
    CascadeMux I__2055 (
            .O(N__12587),
            .I(N__12583));
    CascadeMux I__2054 (
            .O(N__12586),
            .I(N__12580));
    InMux I__2053 (
            .O(N__12583),
            .I(N__12577));
    InMux I__2052 (
            .O(N__12580),
            .I(N__12574));
    LocalMux I__2051 (
            .O(N__12577),
            .I(N__12571));
    LocalMux I__2050 (
            .O(N__12574),
            .I(N__12568));
    Span4Mux_h I__2049 (
            .O(N__12571),
            .I(N__12563));
    Span4Mux_h I__2048 (
            .O(N__12568),
            .I(N__12560));
    InMux I__2047 (
            .O(N__12567),
            .I(N__12555));
    InMux I__2046 (
            .O(N__12566),
            .I(N__12555));
    Odrv4 I__2045 (
            .O(N__12563),
            .I(measured_delay_tr_9));
    Odrv4 I__2044 (
            .O(N__12560),
            .I(measured_delay_tr_9));
    LocalMux I__2043 (
            .O(N__12555),
            .I(measured_delay_tr_9));
    InMux I__2042 (
            .O(N__12548),
            .I(N__12545));
    LocalMux I__2041 (
            .O(N__12545),
            .I(N__12541));
    InMux I__2040 (
            .O(N__12544),
            .I(N__12538));
    Span4Mux_h I__2039 (
            .O(N__12541),
            .I(N__12532));
    LocalMux I__2038 (
            .O(N__12538),
            .I(N__12529));
    InMux I__2037 (
            .O(N__12537),
            .I(N__12522));
    InMux I__2036 (
            .O(N__12536),
            .I(N__12522));
    InMux I__2035 (
            .O(N__12535),
            .I(N__12522));
    Odrv4 I__2034 (
            .O(N__12532),
            .I(\phase_controller_inst1.stoper_tr.N_98 ));
    Odrv4 I__2033 (
            .O(N__12529),
            .I(\phase_controller_inst1.stoper_tr.N_98 ));
    LocalMux I__2032 (
            .O(N__12522),
            .I(\phase_controller_inst1.stoper_tr.N_98 ));
    InMux I__2031 (
            .O(N__12515),
            .I(N__12511));
    InMux I__2030 (
            .O(N__12514),
            .I(N__12508));
    LocalMux I__2029 (
            .O(N__12511),
            .I(phase_controller_inst1_stoper_hc_un1_startlto19_2));
    LocalMux I__2028 (
            .O(N__12508),
            .I(phase_controller_inst1_stoper_hc_un1_startlto19_2));
    CascadeMux I__2027 (
            .O(N__12503),
            .I(phase_controller_inst1_stoper_hc_un1_startlto19_2_cascade_));
    CascadeMux I__2026 (
            .O(N__12500),
            .I(N__12492));
    CascadeMux I__2025 (
            .O(N__12499),
            .I(N__12489));
    CascadeMux I__2024 (
            .O(N__12498),
            .I(N__12486));
    CascadeMux I__2023 (
            .O(N__12497),
            .I(N__12476));
    CascadeMux I__2022 (
            .O(N__12496),
            .I(N__12473));
    CascadeMux I__2021 (
            .O(N__12495),
            .I(N__12470));
    InMux I__2020 (
            .O(N__12492),
            .I(N__12457));
    InMux I__2019 (
            .O(N__12489),
            .I(N__12457));
    InMux I__2018 (
            .O(N__12486),
            .I(N__12457));
    InMux I__2017 (
            .O(N__12485),
            .I(N__12448));
    InMux I__2016 (
            .O(N__12484),
            .I(N__12448));
    InMux I__2015 (
            .O(N__12483),
            .I(N__12448));
    InMux I__2014 (
            .O(N__12482),
            .I(N__12448));
    InMux I__2013 (
            .O(N__12481),
            .I(N__12441));
    InMux I__2012 (
            .O(N__12480),
            .I(N__12441));
    InMux I__2011 (
            .O(N__12479),
            .I(N__12441));
    InMux I__2010 (
            .O(N__12476),
            .I(N__12434));
    InMux I__2009 (
            .O(N__12473),
            .I(N__12434));
    InMux I__2008 (
            .O(N__12470),
            .I(N__12434));
    InMux I__2007 (
            .O(N__12469),
            .I(N__12427));
    InMux I__2006 (
            .O(N__12468),
            .I(N__12427));
    InMux I__2005 (
            .O(N__12467),
            .I(N__12427));
    InMux I__2004 (
            .O(N__12466),
            .I(N__12424));
    InMux I__2003 (
            .O(N__12465),
            .I(N__12421));
    CascadeMux I__2002 (
            .O(N__12464),
            .I(N__12418));
    LocalMux I__2001 (
            .O(N__12457),
            .I(N__12407));
    LocalMux I__2000 (
            .O(N__12448),
            .I(N__12407));
    LocalMux I__1999 (
            .O(N__12441),
            .I(N__12407));
    LocalMux I__1998 (
            .O(N__12434),
            .I(N__12400));
    LocalMux I__1997 (
            .O(N__12427),
            .I(N__12400));
    LocalMux I__1996 (
            .O(N__12424),
            .I(N__12400));
    LocalMux I__1995 (
            .O(N__12421),
            .I(N__12397));
    InMux I__1994 (
            .O(N__12418),
            .I(N__12393));
    InMux I__1993 (
            .O(N__12417),
            .I(N__12388));
    InMux I__1992 (
            .O(N__12416),
            .I(N__12388));
    InMux I__1991 (
            .O(N__12415),
            .I(N__12383));
    InMux I__1990 (
            .O(N__12414),
            .I(N__12383));
    Span4Mux_v I__1989 (
            .O(N__12407),
            .I(N__12378));
    Span4Mux_h I__1988 (
            .O(N__12400),
            .I(N__12378));
    Span4Mux_h I__1987 (
            .O(N__12397),
            .I(N__12375));
    InMux I__1986 (
            .O(N__12396),
            .I(N__12372));
    LocalMux I__1985 (
            .O(N__12393),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__1984 (
            .O(N__12388),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__1983 (
            .O(N__12383),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__1982 (
            .O(N__12378),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__1981 (
            .O(N__12375),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__1980 (
            .O(N__12372),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    InMux I__1979 (
            .O(N__12359),
            .I(N__12326));
    InMux I__1978 (
            .O(N__12358),
            .I(N__12326));
    InMux I__1977 (
            .O(N__12357),
            .I(N__12326));
    InMux I__1976 (
            .O(N__12356),
            .I(N__12326));
    InMux I__1975 (
            .O(N__12355),
            .I(N__12326));
    InMux I__1974 (
            .O(N__12354),
            .I(N__12326));
    InMux I__1973 (
            .O(N__12353),
            .I(N__12326));
    InMux I__1972 (
            .O(N__12352),
            .I(N__12319));
    InMux I__1971 (
            .O(N__12351),
            .I(N__12319));
    InMux I__1970 (
            .O(N__12350),
            .I(N__12319));
    InMux I__1969 (
            .O(N__12349),
            .I(N__12306));
    InMux I__1968 (
            .O(N__12348),
            .I(N__12306));
    InMux I__1967 (
            .O(N__12347),
            .I(N__12306));
    InMux I__1966 (
            .O(N__12346),
            .I(N__12306));
    InMux I__1965 (
            .O(N__12345),
            .I(N__12306));
    InMux I__1964 (
            .O(N__12344),
            .I(N__12306));
    InMux I__1963 (
            .O(N__12343),
            .I(N__12303));
    InMux I__1962 (
            .O(N__12342),
            .I(N__12300));
    CascadeMux I__1961 (
            .O(N__12341),
            .I(N__12297));
    LocalMux I__1960 (
            .O(N__12326),
            .I(N__12288));
    LocalMux I__1959 (
            .O(N__12319),
            .I(N__12288));
    LocalMux I__1958 (
            .O(N__12306),
            .I(N__12283));
    LocalMux I__1957 (
            .O(N__12303),
            .I(N__12283));
    LocalMux I__1956 (
            .O(N__12300),
            .I(N__12280));
    InMux I__1955 (
            .O(N__12297),
            .I(N__12274));
    InMux I__1954 (
            .O(N__12296),
            .I(N__12274));
    InMux I__1953 (
            .O(N__12295),
            .I(N__12267));
    InMux I__1952 (
            .O(N__12294),
            .I(N__12267));
    InMux I__1951 (
            .O(N__12293),
            .I(N__12267));
    Span4Mux_v I__1950 (
            .O(N__12288),
            .I(N__12262));
    Span4Mux_h I__1949 (
            .O(N__12283),
            .I(N__12262));
    Span4Mux_h I__1948 (
            .O(N__12280),
            .I(N__12259));
    InMux I__1947 (
            .O(N__12279),
            .I(N__12256));
    LocalMux I__1946 (
            .O(N__12274),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__1945 (
            .O(N__12267),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__1944 (
            .O(N__12262),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__1943 (
            .O(N__12259),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    LocalMux I__1942 (
            .O(N__12256),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    CEMux I__1941 (
            .O(N__12245),
            .I(N__12242));
    LocalMux I__1940 (
            .O(N__12242),
            .I(N__12236));
    CEMux I__1939 (
            .O(N__12241),
            .I(N__12233));
    CEMux I__1938 (
            .O(N__12240),
            .I(N__12230));
    CEMux I__1937 (
            .O(N__12239),
            .I(N__12227));
    Span4Mux_v I__1936 (
            .O(N__12236),
            .I(N__12224));
    LocalMux I__1935 (
            .O(N__12233),
            .I(N__12221));
    LocalMux I__1934 (
            .O(N__12230),
            .I(N__12218));
    LocalMux I__1933 (
            .O(N__12227),
            .I(N__12215));
    Span4Mux_h I__1932 (
            .O(N__12224),
            .I(N__12212));
    Span4Mux_h I__1931 (
            .O(N__12221),
            .I(N__12209));
    Span4Mux_h I__1930 (
            .O(N__12218),
            .I(N__12206));
    Span4Mux_h I__1929 (
            .O(N__12215),
            .I(N__12203));
    Odrv4 I__1928 (
            .O(N__12212),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__1927 (
            .O(N__12209),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__1926 (
            .O(N__12206),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__1925 (
            .O(N__12203),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    InMux I__1924 (
            .O(N__12194),
            .I(N__12191));
    LocalMux I__1923 (
            .O(N__12191),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_a0Z0Z_1 ));
    CascadeMux I__1922 (
            .O(N__12188),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto31_aZ0Z2_cascade_ ));
    InMux I__1921 (
            .O(N__12185),
            .I(N__12181));
    InMux I__1920 (
            .O(N__12184),
            .I(N__12178));
    LocalMux I__1919 (
            .O(N__12181),
            .I(d_N_5_mux));
    LocalMux I__1918 (
            .O(N__12178),
            .I(d_N_5_mux));
    InMux I__1917 (
            .O(N__12173),
            .I(N__12170));
    LocalMux I__1916 (
            .O(N__12170),
            .I(N__12167));
    Odrv4 I__1915 (
            .O(N__12167),
            .I(\phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_1 ));
    CascadeMux I__1914 (
            .O(N__12164),
            .I(\phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_2_cascade_ ));
    InMux I__1913 (
            .O(N__12161),
            .I(N__12157));
    InMux I__1912 (
            .O(N__12160),
            .I(N__12154));
    LocalMux I__1911 (
            .O(N__12157),
            .I(N__12151));
    LocalMux I__1910 (
            .O(N__12154),
            .I(\phase_controller_inst1.stoper_hc.un1_N_6_mux ));
    Odrv4 I__1909 (
            .O(N__12151),
            .I(\phase_controller_inst1.stoper_hc.un1_N_6_mux ));
    CascadeMux I__1908 (
            .O(N__12146),
            .I(N__12143));
    InMux I__1907 (
            .O(N__12143),
            .I(N__12140));
    LocalMux I__1906 (
            .O(N__12140),
            .I(\phase_controller_inst1.stoper_hc.un1_m3_eZ0Z_1 ));
    InMux I__1905 (
            .O(N__12137),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    CascadeMux I__1904 (
            .O(N__12134),
            .I(N__12129));
    CascadeMux I__1903 (
            .O(N__12133),
            .I(N__12126));
    InMux I__1902 (
            .O(N__12132),
            .I(N__12123));
    InMux I__1901 (
            .O(N__12129),
            .I(N__12118));
    InMux I__1900 (
            .O(N__12126),
            .I(N__12118));
    LocalMux I__1899 (
            .O(N__12123),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__1898 (
            .O(N__12118),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__1897 (
            .O(N__12113),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    CascadeMux I__1896 (
            .O(N__12110),
            .I(N__12105));
    CascadeMux I__1895 (
            .O(N__12109),
            .I(N__12102));
    InMux I__1894 (
            .O(N__12108),
            .I(N__12099));
    InMux I__1893 (
            .O(N__12105),
            .I(N__12094));
    InMux I__1892 (
            .O(N__12102),
            .I(N__12094));
    LocalMux I__1891 (
            .O(N__12099),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__1890 (
            .O(N__12094),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__1889 (
            .O(N__12089),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__1888 (
            .O(N__12086),
            .I(N__12081));
    InMux I__1887 (
            .O(N__12085),
            .I(N__12078));
    InMux I__1886 (
            .O(N__12084),
            .I(N__12075));
    LocalMux I__1885 (
            .O(N__12081),
            .I(N__12072));
    LocalMux I__1884 (
            .O(N__12078),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__1883 (
            .O(N__12075),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__1882 (
            .O(N__12072),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__1881 (
            .O(N__12065),
            .I(bfn_5_18_0_));
    InMux I__1880 (
            .O(N__12062),
            .I(N__12057));
    InMux I__1879 (
            .O(N__12061),
            .I(N__12054));
    InMux I__1878 (
            .O(N__12060),
            .I(N__12051));
    LocalMux I__1877 (
            .O(N__12057),
            .I(N__12048));
    LocalMux I__1876 (
            .O(N__12054),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__1875 (
            .O(N__12051),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv4 I__1874 (
            .O(N__12048),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__1873 (
            .O(N__12041),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    CascadeMux I__1872 (
            .O(N__12038),
            .I(N__12033));
    CascadeMux I__1871 (
            .O(N__12037),
            .I(N__12030));
    InMux I__1870 (
            .O(N__12036),
            .I(N__12027));
    InMux I__1869 (
            .O(N__12033),
            .I(N__12022));
    InMux I__1868 (
            .O(N__12030),
            .I(N__12022));
    LocalMux I__1867 (
            .O(N__12027),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__1866 (
            .O(N__12022),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__1865 (
            .O(N__12017),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    CascadeMux I__1864 (
            .O(N__12014),
            .I(N__12009));
    CascadeMux I__1863 (
            .O(N__12013),
            .I(N__12006));
    InMux I__1862 (
            .O(N__12012),
            .I(N__12003));
    InMux I__1861 (
            .O(N__12009),
            .I(N__11998));
    InMux I__1860 (
            .O(N__12006),
            .I(N__11998));
    LocalMux I__1859 (
            .O(N__12003),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__1858 (
            .O(N__11998),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__1857 (
            .O(N__11993),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__1856 (
            .O(N__11990),
            .I(N__11986));
    InMux I__1855 (
            .O(N__11989),
            .I(N__11983));
    LocalMux I__1854 (
            .O(N__11986),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__1853 (
            .O(N__11983),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__1852 (
            .O(N__11978),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__1851 (
            .O(N__11975),
            .I(N__11937));
    InMux I__1850 (
            .O(N__11974),
            .I(N__11937));
    InMux I__1849 (
            .O(N__11973),
            .I(N__11937));
    InMux I__1848 (
            .O(N__11972),
            .I(N__11937));
    InMux I__1847 (
            .O(N__11971),
            .I(N__11928));
    InMux I__1846 (
            .O(N__11970),
            .I(N__11928));
    InMux I__1845 (
            .O(N__11969),
            .I(N__11928));
    InMux I__1844 (
            .O(N__11968),
            .I(N__11928));
    InMux I__1843 (
            .O(N__11967),
            .I(N__11923));
    InMux I__1842 (
            .O(N__11966),
            .I(N__11923));
    InMux I__1841 (
            .O(N__11965),
            .I(N__11914));
    InMux I__1840 (
            .O(N__11964),
            .I(N__11914));
    InMux I__1839 (
            .O(N__11963),
            .I(N__11914));
    InMux I__1838 (
            .O(N__11962),
            .I(N__11914));
    InMux I__1837 (
            .O(N__11961),
            .I(N__11905));
    InMux I__1836 (
            .O(N__11960),
            .I(N__11905));
    InMux I__1835 (
            .O(N__11959),
            .I(N__11905));
    InMux I__1834 (
            .O(N__11958),
            .I(N__11905));
    InMux I__1833 (
            .O(N__11957),
            .I(N__11896));
    InMux I__1832 (
            .O(N__11956),
            .I(N__11896));
    InMux I__1831 (
            .O(N__11955),
            .I(N__11896));
    InMux I__1830 (
            .O(N__11954),
            .I(N__11896));
    InMux I__1829 (
            .O(N__11953),
            .I(N__11887));
    InMux I__1828 (
            .O(N__11952),
            .I(N__11887));
    InMux I__1827 (
            .O(N__11951),
            .I(N__11887));
    InMux I__1826 (
            .O(N__11950),
            .I(N__11887));
    InMux I__1825 (
            .O(N__11949),
            .I(N__11878));
    InMux I__1824 (
            .O(N__11948),
            .I(N__11878));
    InMux I__1823 (
            .O(N__11947),
            .I(N__11878));
    InMux I__1822 (
            .O(N__11946),
            .I(N__11878));
    LocalMux I__1821 (
            .O(N__11937),
            .I(N__11875));
    LocalMux I__1820 (
            .O(N__11928),
            .I(N__11860));
    LocalMux I__1819 (
            .O(N__11923),
            .I(N__11860));
    LocalMux I__1818 (
            .O(N__11914),
            .I(N__11860));
    LocalMux I__1817 (
            .O(N__11905),
            .I(N__11860));
    LocalMux I__1816 (
            .O(N__11896),
            .I(N__11860));
    LocalMux I__1815 (
            .O(N__11887),
            .I(N__11860));
    LocalMux I__1814 (
            .O(N__11878),
            .I(N__11860));
    Odrv4 I__1813 (
            .O(N__11875),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv12 I__1812 (
            .O(N__11860),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__1811 (
            .O(N__11855),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    InMux I__1810 (
            .O(N__11852),
            .I(N__11848));
    InMux I__1809 (
            .O(N__11851),
            .I(N__11845));
    LocalMux I__1808 (
            .O(N__11848),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__1807 (
            .O(N__11845),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CEMux I__1806 (
            .O(N__11840),
            .I(N__11828));
    CEMux I__1805 (
            .O(N__11839),
            .I(N__11828));
    CEMux I__1804 (
            .O(N__11838),
            .I(N__11828));
    CEMux I__1803 (
            .O(N__11837),
            .I(N__11828));
    GlobalMux I__1802 (
            .O(N__11828),
            .I(N__11825));
    gio2CtrlBuf I__1801 (
            .O(N__11825),
            .I(\delay_measurement_inst.delay_tr_timer.N_139_i_g ));
    InMux I__1800 (
            .O(N__11822),
            .I(N__11817));
    InMux I__1799 (
            .O(N__11821),
            .I(N__11812));
    InMux I__1798 (
            .O(N__11820),
            .I(N__11812));
    LocalMux I__1797 (
            .O(N__11817),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__1796 (
            .O(N__11812),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__1795 (
            .O(N__11807),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    CascadeMux I__1794 (
            .O(N__11804),
            .I(N__11799));
    CascadeMux I__1793 (
            .O(N__11803),
            .I(N__11796));
    InMux I__1792 (
            .O(N__11802),
            .I(N__11793));
    InMux I__1791 (
            .O(N__11799),
            .I(N__11788));
    InMux I__1790 (
            .O(N__11796),
            .I(N__11788));
    LocalMux I__1789 (
            .O(N__11793),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__1788 (
            .O(N__11788),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__1787 (
            .O(N__11783),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    CascadeMux I__1786 (
            .O(N__11780),
            .I(N__11775));
    CascadeMux I__1785 (
            .O(N__11779),
            .I(N__11772));
    InMux I__1784 (
            .O(N__11778),
            .I(N__11769));
    InMux I__1783 (
            .O(N__11775),
            .I(N__11764));
    InMux I__1782 (
            .O(N__11772),
            .I(N__11764));
    LocalMux I__1781 (
            .O(N__11769),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__1780 (
            .O(N__11764),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__1779 (
            .O(N__11759),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__1778 (
            .O(N__11756),
            .I(N__11751));
    InMux I__1777 (
            .O(N__11755),
            .I(N__11748));
    InMux I__1776 (
            .O(N__11754),
            .I(N__11745));
    LocalMux I__1775 (
            .O(N__11751),
            .I(N__11742));
    LocalMux I__1774 (
            .O(N__11748),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__1773 (
            .O(N__11745),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv4 I__1772 (
            .O(N__11742),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__1771 (
            .O(N__11735),
            .I(bfn_5_17_0_));
    InMux I__1770 (
            .O(N__11732),
            .I(N__11727));
    InMux I__1769 (
            .O(N__11731),
            .I(N__11724));
    InMux I__1768 (
            .O(N__11730),
            .I(N__11721));
    LocalMux I__1767 (
            .O(N__11727),
            .I(N__11718));
    LocalMux I__1766 (
            .O(N__11724),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__1765 (
            .O(N__11721),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__1764 (
            .O(N__11718),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__1763 (
            .O(N__11711),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    CascadeMux I__1762 (
            .O(N__11708),
            .I(N__11703));
    CascadeMux I__1761 (
            .O(N__11707),
            .I(N__11700));
    InMux I__1760 (
            .O(N__11706),
            .I(N__11697));
    InMux I__1759 (
            .O(N__11703),
            .I(N__11692));
    InMux I__1758 (
            .O(N__11700),
            .I(N__11692));
    LocalMux I__1757 (
            .O(N__11697),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__1756 (
            .O(N__11692),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__1755 (
            .O(N__11687),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    CascadeMux I__1754 (
            .O(N__11684),
            .I(N__11679));
    CascadeMux I__1753 (
            .O(N__11683),
            .I(N__11676));
    InMux I__1752 (
            .O(N__11682),
            .I(N__11673));
    InMux I__1751 (
            .O(N__11679),
            .I(N__11668));
    InMux I__1750 (
            .O(N__11676),
            .I(N__11668));
    LocalMux I__1749 (
            .O(N__11673),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__1748 (
            .O(N__11668),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__1747 (
            .O(N__11663),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__1746 (
            .O(N__11660),
            .I(N__11655));
    InMux I__1745 (
            .O(N__11659),
            .I(N__11650));
    InMux I__1744 (
            .O(N__11658),
            .I(N__11650));
    LocalMux I__1743 (
            .O(N__11655),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__1742 (
            .O(N__11650),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__1741 (
            .O(N__11645),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__1740 (
            .O(N__11642),
            .I(N__11637));
    InMux I__1739 (
            .O(N__11641),
            .I(N__11632));
    InMux I__1738 (
            .O(N__11640),
            .I(N__11632));
    LocalMux I__1737 (
            .O(N__11637),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__1736 (
            .O(N__11632),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__1735 (
            .O(N__11627),
            .I(N__11622));
    InMux I__1734 (
            .O(N__11626),
            .I(N__11617));
    InMux I__1733 (
            .O(N__11625),
            .I(N__11617));
    LocalMux I__1732 (
            .O(N__11622),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__1731 (
            .O(N__11617),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__1730 (
            .O(N__11612),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    CascadeMux I__1729 (
            .O(N__11609),
            .I(N__11604));
    CascadeMux I__1728 (
            .O(N__11608),
            .I(N__11601));
    InMux I__1727 (
            .O(N__11607),
            .I(N__11598));
    InMux I__1726 (
            .O(N__11604),
            .I(N__11593));
    InMux I__1725 (
            .O(N__11601),
            .I(N__11593));
    LocalMux I__1724 (
            .O(N__11598),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__1723 (
            .O(N__11593),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__1722 (
            .O(N__11588),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    CascadeMux I__1721 (
            .O(N__11585),
            .I(N__11580));
    CascadeMux I__1720 (
            .O(N__11584),
            .I(N__11577));
    InMux I__1719 (
            .O(N__11583),
            .I(N__11574));
    InMux I__1718 (
            .O(N__11580),
            .I(N__11569));
    InMux I__1717 (
            .O(N__11577),
            .I(N__11569));
    LocalMux I__1716 (
            .O(N__11574),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__1715 (
            .O(N__11569),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__1714 (
            .O(N__11564),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__1713 (
            .O(N__11561),
            .I(N__11556));
    InMux I__1712 (
            .O(N__11560),
            .I(N__11553));
    InMux I__1711 (
            .O(N__11559),
            .I(N__11550));
    LocalMux I__1710 (
            .O(N__11556),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__1709 (
            .O(N__11553),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__1708 (
            .O(N__11550),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__1707 (
            .O(N__11543),
            .I(bfn_5_16_0_));
    InMux I__1706 (
            .O(N__11540),
            .I(N__11535));
    InMux I__1705 (
            .O(N__11539),
            .I(N__11532));
    InMux I__1704 (
            .O(N__11538),
            .I(N__11529));
    LocalMux I__1703 (
            .O(N__11535),
            .I(N__11526));
    LocalMux I__1702 (
            .O(N__11532),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__1701 (
            .O(N__11529),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    Odrv4 I__1700 (
            .O(N__11526),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__1699 (
            .O(N__11519),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    CascadeMux I__1698 (
            .O(N__11516),
            .I(N__11511));
    CascadeMux I__1697 (
            .O(N__11515),
            .I(N__11508));
    InMux I__1696 (
            .O(N__11514),
            .I(N__11505));
    InMux I__1695 (
            .O(N__11511),
            .I(N__11500));
    InMux I__1694 (
            .O(N__11508),
            .I(N__11500));
    LocalMux I__1693 (
            .O(N__11505),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__1692 (
            .O(N__11500),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__1691 (
            .O(N__11495),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    CascadeMux I__1690 (
            .O(N__11492),
            .I(N__11487));
    CascadeMux I__1689 (
            .O(N__11491),
            .I(N__11484));
    InMux I__1688 (
            .O(N__11490),
            .I(N__11481));
    InMux I__1687 (
            .O(N__11487),
            .I(N__11476));
    InMux I__1686 (
            .O(N__11484),
            .I(N__11476));
    LocalMux I__1685 (
            .O(N__11481),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__1684 (
            .O(N__11476),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__1683 (
            .O(N__11471),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__1682 (
            .O(N__11468),
            .I(N__11463));
    InMux I__1681 (
            .O(N__11467),
            .I(N__11458));
    InMux I__1680 (
            .O(N__11466),
            .I(N__11458));
    LocalMux I__1679 (
            .O(N__11463),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__1678 (
            .O(N__11458),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__1677 (
            .O(N__11453),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__1676 (
            .O(N__11450),
            .I(N__11445));
    InMux I__1675 (
            .O(N__11449),
            .I(N__11440));
    InMux I__1674 (
            .O(N__11448),
            .I(N__11440));
    LocalMux I__1673 (
            .O(N__11445),
            .I(N__11437));
    LocalMux I__1672 (
            .O(N__11440),
            .I(N__11434));
    Odrv4 I__1671 (
            .O(N__11437),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    Odrv4 I__1670 (
            .O(N__11434),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    CascadeMux I__1669 (
            .O(N__11429),
            .I(N__11424));
    InMux I__1668 (
            .O(N__11428),
            .I(N__11421));
    InMux I__1667 (
            .O(N__11427),
            .I(N__11416));
    InMux I__1666 (
            .O(N__11424),
            .I(N__11416));
    LocalMux I__1665 (
            .O(N__11421),
            .I(N__11413));
    LocalMux I__1664 (
            .O(N__11416),
            .I(N__11410));
    Odrv4 I__1663 (
            .O(N__11413),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    Odrv4 I__1662 (
            .O(N__11410),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    CascadeMux I__1661 (
            .O(N__11405),
            .I(N__11401));
    InMux I__1660 (
            .O(N__11404),
            .I(N__11397));
    InMux I__1659 (
            .O(N__11401),
            .I(N__11392));
    InMux I__1658 (
            .O(N__11400),
            .I(N__11392));
    LocalMux I__1657 (
            .O(N__11397),
            .I(N__11389));
    LocalMux I__1656 (
            .O(N__11392),
            .I(N__11386));
    Odrv4 I__1655 (
            .O(N__11389),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    Odrv4 I__1654 (
            .O(N__11386),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    InMux I__1653 (
            .O(N__11381),
            .I(N__11370));
    InMux I__1652 (
            .O(N__11380),
            .I(N__11370));
    InMux I__1651 (
            .O(N__11379),
            .I(N__11370));
    InMux I__1650 (
            .O(N__11378),
            .I(N__11365));
    InMux I__1649 (
            .O(N__11377),
            .I(N__11365));
    LocalMux I__1648 (
            .O(N__11370),
            .I(N__11357));
    LocalMux I__1647 (
            .O(N__11365),
            .I(N__11354));
    InMux I__1646 (
            .O(N__11364),
            .I(N__11347));
    InMux I__1645 (
            .O(N__11363),
            .I(N__11347));
    InMux I__1644 (
            .O(N__11362),
            .I(N__11347));
    InMux I__1643 (
            .O(N__11361),
            .I(N__11342));
    InMux I__1642 (
            .O(N__11360),
            .I(N__11342));
    Span4Mux_h I__1641 (
            .O(N__11357),
            .I(N__11339));
    Span4Mux_v I__1640 (
            .O(N__11354),
            .I(N__11336));
    LocalMux I__1639 (
            .O(N__11347),
            .I(N__11331));
    LocalMux I__1638 (
            .O(N__11342),
            .I(N__11331));
    Odrv4 I__1637 (
            .O(N__11339),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ));
    Odrv4 I__1636 (
            .O(N__11336),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ));
    Odrv12 I__1635 (
            .O(N__11331),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ));
    InMux I__1634 (
            .O(N__11324),
            .I(N__11315));
    InMux I__1633 (
            .O(N__11323),
            .I(N__11315));
    InMux I__1632 (
            .O(N__11322),
            .I(N__11308));
    InMux I__1631 (
            .O(N__11321),
            .I(N__11308));
    InMux I__1630 (
            .O(N__11320),
            .I(N__11308));
    LocalMux I__1629 (
            .O(N__11315),
            .I(\delay_measurement_inst.N_197_1 ));
    LocalMux I__1628 (
            .O(N__11308),
            .I(\delay_measurement_inst.N_197_1 ));
    CascadeMux I__1627 (
            .O(N__11303),
            .I(N__11299));
    InMux I__1626 (
            .O(N__11302),
            .I(N__11296));
    InMux I__1625 (
            .O(N__11299),
            .I(N__11293));
    LocalMux I__1624 (
            .O(N__11296),
            .I(N__11290));
    LocalMux I__1623 (
            .O(N__11293),
            .I(N__11287));
    Odrv4 I__1622 (
            .O(N__11290),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    Odrv4 I__1621 (
            .O(N__11287),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    CEMux I__1620 (
            .O(N__11282),
            .I(N__11278));
    CEMux I__1619 (
            .O(N__11281),
            .I(N__11275));
    LocalMux I__1618 (
            .O(N__11278),
            .I(N__11271));
    LocalMux I__1617 (
            .O(N__11275),
            .I(N__11268));
    CEMux I__1616 (
            .O(N__11274),
            .I(N__11265));
    Span4Mux_h I__1615 (
            .O(N__11271),
            .I(N__11262));
    Span4Mux_v I__1614 (
            .O(N__11268),
            .I(N__11259));
    LocalMux I__1613 (
            .O(N__11265),
            .I(N__11256));
    Odrv4 I__1612 (
            .O(N__11262),
            .I(\delay_measurement_inst.N_81_i_0 ));
    Odrv4 I__1611 (
            .O(N__11259),
            .I(\delay_measurement_inst.N_81_i_0 ));
    Odrv4 I__1610 (
            .O(N__11256),
            .I(\delay_measurement_inst.N_81_i_0 ));
    InMux I__1609 (
            .O(N__11249),
            .I(N__11246));
    LocalMux I__1608 (
            .O(N__11246),
            .I(N__11243));
    Span4Mux_v I__1607 (
            .O(N__11243),
            .I(N__11239));
    InMux I__1606 (
            .O(N__11242),
            .I(N__11236));
    Span4Mux_h I__1605 (
            .O(N__11239),
            .I(N__11232));
    LocalMux I__1604 (
            .O(N__11236),
            .I(N__11229));
    InMux I__1603 (
            .O(N__11235),
            .I(N__11226));
    Odrv4 I__1602 (
            .O(N__11232),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    Odrv4 I__1601 (
            .O(N__11229),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__1600 (
            .O(N__11226),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__1599 (
            .O(N__11219),
            .I(bfn_5_15_0_));
    InMux I__1598 (
            .O(N__11216),
            .I(N__11213));
    LocalMux I__1597 (
            .O(N__11213),
            .I(N__11210));
    Span4Mux_h I__1596 (
            .O(N__11210),
            .I(N__11205));
    InMux I__1595 (
            .O(N__11209),
            .I(N__11202));
    InMux I__1594 (
            .O(N__11208),
            .I(N__11199));
    Odrv4 I__1593 (
            .O(N__11205),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__1592 (
            .O(N__11202),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__1591 (
            .O(N__11199),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__1590 (
            .O(N__11192),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    CascadeMux I__1589 (
            .O(N__11189),
            .I(N__11184));
    CascadeMux I__1588 (
            .O(N__11188),
            .I(N__11181));
    InMux I__1587 (
            .O(N__11187),
            .I(N__11178));
    InMux I__1586 (
            .O(N__11184),
            .I(N__11173));
    InMux I__1585 (
            .O(N__11181),
            .I(N__11173));
    LocalMux I__1584 (
            .O(N__11178),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__1583 (
            .O(N__11173),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__1582 (
            .O(N__11168),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    CascadeMux I__1581 (
            .O(N__11165),
            .I(N__11160));
    CascadeMux I__1580 (
            .O(N__11164),
            .I(N__11157));
    InMux I__1579 (
            .O(N__11163),
            .I(N__11154));
    InMux I__1578 (
            .O(N__11160),
            .I(N__11149));
    InMux I__1577 (
            .O(N__11157),
            .I(N__11149));
    LocalMux I__1576 (
            .O(N__11154),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__1575 (
            .O(N__11149),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__1574 (
            .O(N__11144),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__1573 (
            .O(N__11141),
            .I(N__11136));
    InMux I__1572 (
            .O(N__11140),
            .I(N__11131));
    InMux I__1571 (
            .O(N__11139),
            .I(N__11131));
    LocalMux I__1570 (
            .O(N__11136),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__1569 (
            .O(N__11131),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__1568 (
            .O(N__11126),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    CascadeMux I__1567 (
            .O(N__11123),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_4Z0Z_3_cascade_ ));
    InMux I__1566 (
            .O(N__11120),
            .I(N__11117));
    LocalMux I__1565 (
            .O(N__11117),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3 ));
    CascadeMux I__1564 (
            .O(N__11114),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_6Z0Z_3_cascade_ ));
    InMux I__1563 (
            .O(N__11111),
            .I(N__11108));
    LocalMux I__1562 (
            .O(N__11108),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0Z0Z_6 ));
    CascadeMux I__1561 (
            .O(N__11105),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0Z0Z_6_cascade_ ));
    CascadeMux I__1560 (
            .O(N__11102),
            .I(\phase_controller_inst1.stoper_tr.N_92_cascade_ ));
    CascadeMux I__1559 (
            .O(N__11099),
            .I(N__11095));
    CascadeMux I__1558 (
            .O(N__11098),
            .I(N__11091));
    InMux I__1557 (
            .O(N__11095),
            .I(N__11087));
    InMux I__1556 (
            .O(N__11094),
            .I(N__11084));
    InMux I__1555 (
            .O(N__11091),
            .I(N__11079));
    InMux I__1554 (
            .O(N__11090),
            .I(N__11079));
    LocalMux I__1553 (
            .O(N__11087),
            .I(\delay_measurement_inst.elapsed_time_tr_9 ));
    LocalMux I__1552 (
            .O(N__11084),
            .I(\delay_measurement_inst.elapsed_time_tr_9 ));
    LocalMux I__1551 (
            .O(N__11079),
            .I(\delay_measurement_inst.elapsed_time_tr_9 ));
    InMux I__1550 (
            .O(N__11072),
            .I(N__11061));
    InMux I__1549 (
            .O(N__11071),
            .I(N__11061));
    InMux I__1548 (
            .O(N__11070),
            .I(N__11049));
    InMux I__1547 (
            .O(N__11069),
            .I(N__11049));
    InMux I__1546 (
            .O(N__11068),
            .I(N__11049));
    InMux I__1545 (
            .O(N__11067),
            .I(N__11049));
    InMux I__1544 (
            .O(N__11066),
            .I(N__11049));
    LocalMux I__1543 (
            .O(N__11061),
            .I(N__11046));
    InMux I__1542 (
            .O(N__11060),
            .I(N__11043));
    LocalMux I__1541 (
            .O(N__11049),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ));
    Odrv4 I__1540 (
            .O(N__11046),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ));
    LocalMux I__1539 (
            .O(N__11043),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ));
    CascadeMux I__1538 (
            .O(N__11036),
            .I(N__11026));
    InMux I__1537 (
            .O(N__11035),
            .I(N__11023));
    InMux I__1536 (
            .O(N__11034),
            .I(N__11018));
    InMux I__1535 (
            .O(N__11033),
            .I(N__11018));
    InMux I__1534 (
            .O(N__11032),
            .I(N__11007));
    InMux I__1533 (
            .O(N__11031),
            .I(N__11007));
    InMux I__1532 (
            .O(N__11030),
            .I(N__11007));
    InMux I__1531 (
            .O(N__11029),
            .I(N__11007));
    InMux I__1530 (
            .O(N__11026),
            .I(N__11007));
    LocalMux I__1529 (
            .O(N__11023),
            .I(\delay_measurement_inst.N_165 ));
    LocalMux I__1528 (
            .O(N__11018),
            .I(\delay_measurement_inst.N_165 ));
    LocalMux I__1527 (
            .O(N__11007),
            .I(\delay_measurement_inst.N_165 ));
    CascadeMux I__1526 (
            .O(N__11000),
            .I(N__10995));
    CascadeMux I__1525 (
            .O(N__10999),
            .I(N__10992));
    CascadeMux I__1524 (
            .O(N__10998),
            .I(N__10987));
    InMux I__1523 (
            .O(N__10995),
            .I(N__10983));
    InMux I__1522 (
            .O(N__10992),
            .I(N__10972));
    InMux I__1521 (
            .O(N__10991),
            .I(N__10972));
    InMux I__1520 (
            .O(N__10990),
            .I(N__10972));
    InMux I__1519 (
            .O(N__10987),
            .I(N__10972));
    InMux I__1518 (
            .O(N__10986),
            .I(N__10972));
    LocalMux I__1517 (
            .O(N__10983),
            .I(N__10969));
    LocalMux I__1516 (
            .O(N__10972),
            .I(N__10966));
    Odrv4 I__1515 (
            .O(N__10969),
            .I(\delay_measurement_inst.N_212 ));
    Odrv4 I__1514 (
            .O(N__10966),
            .I(\delay_measurement_inst.N_212 ));
    InMux I__1513 (
            .O(N__10961),
            .I(N__10957));
    InMux I__1512 (
            .O(N__10960),
            .I(N__10954));
    LocalMux I__1511 (
            .O(N__10957),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    LocalMux I__1510 (
            .O(N__10954),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    CascadeMux I__1509 (
            .O(N__10949),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10_cascade_ ));
    InMux I__1508 (
            .O(N__10946),
            .I(N__10943));
    LocalMux I__1507 (
            .O(N__10943),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ));
    InMux I__1506 (
            .O(N__10940),
            .I(N__10937));
    LocalMux I__1505 (
            .O(N__10937),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ));
    CascadeMux I__1504 (
            .O(N__10934),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_15_cascade_ ));
    InMux I__1503 (
            .O(N__10931),
            .I(N__10928));
    LocalMux I__1502 (
            .O(N__10928),
            .I(N__10925));
    Span12Mux_v I__1501 (
            .O(N__10925),
            .I(N__10922));
    Odrv12 I__1500 (
            .O(N__10922),
            .I(il_max_comp2_c));
    InMux I__1499 (
            .O(N__10919),
            .I(N__10916));
    LocalMux I__1498 (
            .O(N__10916),
            .I(il_max_comp2_D1));
    InMux I__1497 (
            .O(N__10913),
            .I(N__10910));
    LocalMux I__1496 (
            .O(N__10910),
            .I(N__10907));
    Odrv4 I__1495 (
            .O(N__10907),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ));
    InMux I__1494 (
            .O(N__10904),
            .I(N__10901));
    LocalMux I__1493 (
            .O(N__10901),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ));
    InMux I__1492 (
            .O(N__10898),
            .I(N__10895));
    LocalMux I__1491 (
            .O(N__10895),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ));
    InMux I__1490 (
            .O(N__10892),
            .I(N__10889));
    LocalMux I__1489 (
            .O(N__10889),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ));
    InMux I__1488 (
            .O(N__10886),
            .I(N__10883));
    LocalMux I__1487 (
            .O(N__10883),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ));
    InMux I__1486 (
            .O(N__10880),
            .I(N__10877));
    LocalMux I__1485 (
            .O(N__10877),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ));
    InMux I__1484 (
            .O(N__10874),
            .I(N__10871));
    LocalMux I__1483 (
            .O(N__10871),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ));
    InMux I__1482 (
            .O(N__10868),
            .I(N__10865));
    LocalMux I__1481 (
            .O(N__10865),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ));
    InMux I__1480 (
            .O(N__10862),
            .I(N__10859));
    LocalMux I__1479 (
            .O(N__10859),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ));
    InMux I__1478 (
            .O(N__10856),
            .I(N__10853));
    LocalMux I__1477 (
            .O(N__10853),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ));
    InMux I__1476 (
            .O(N__10850),
            .I(N__10847));
    LocalMux I__1475 (
            .O(N__10847),
            .I(N__10844));
    Odrv4 I__1474 (
            .O(N__10844),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ));
    InMux I__1473 (
            .O(N__10841),
            .I(N__10838));
    LocalMux I__1472 (
            .O(N__10838),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_0 ));
    InMux I__1471 (
            .O(N__10835),
            .I(N__10832));
    LocalMux I__1470 (
            .O(N__10832),
            .I(N__10829));
    Odrv4 I__1469 (
            .O(N__10829),
            .I(\phase_controller_slave.stoper_hc.target_timeZ1Z_6 ));
    InMux I__1468 (
            .O(N__10826),
            .I(N__10823));
    LocalMux I__1467 (
            .O(N__10823),
            .I(N__10820));
    Odrv4 I__1466 (
            .O(N__10820),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ));
    InMux I__1465 (
            .O(N__10817),
            .I(N__10814));
    LocalMux I__1464 (
            .O(N__10814),
            .I(N__10811));
    Odrv4 I__1463 (
            .O(N__10811),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ));
    InMux I__1462 (
            .O(N__10808),
            .I(N__10805));
    LocalMux I__1461 (
            .O(N__10805),
            .I(N__10802));
    Odrv4 I__1460 (
            .O(N__10802),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ));
    InMux I__1459 (
            .O(N__10799),
            .I(N__10796));
    LocalMux I__1458 (
            .O(N__10796),
            .I(N__10793));
    Odrv4 I__1457 (
            .O(N__10793),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ));
    InMux I__1456 (
            .O(N__10790),
            .I(N__10787));
    LocalMux I__1455 (
            .O(N__10787),
            .I(N__10784));
    Odrv4 I__1454 (
            .O(N__10784),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__1453 (
            .O(N__10781),
            .I(N__10778));
    InMux I__1452 (
            .O(N__10778),
            .I(N__10775));
    LocalMux I__1451 (
            .O(N__10775),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__1450 (
            .O(N__10772),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__1449 (
            .O(N__10769),
            .I(N__10766));
    LocalMux I__1448 (
            .O(N__10766),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__1447 (
            .O(N__10763),
            .I(bfn_4_18_0_));
    InMux I__1446 (
            .O(N__10760),
            .I(N__10757));
    LocalMux I__1445 (
            .O(N__10757),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__1444 (
            .O(N__10754),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__1443 (
            .O(N__10751),
            .I(N__10748));
    LocalMux I__1442 (
            .O(N__10748),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__1441 (
            .O(N__10745),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__1440 (
            .O(N__10742),
            .I(N__10739));
    InMux I__1439 (
            .O(N__10739),
            .I(N__10736));
    LocalMux I__1438 (
            .O(N__10736),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ));
    InMux I__1437 (
            .O(N__10733),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__1436 (
            .O(N__10730),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CEMux I__1435 (
            .O(N__10727),
            .I(N__10712));
    CEMux I__1434 (
            .O(N__10726),
            .I(N__10712));
    CEMux I__1433 (
            .O(N__10725),
            .I(N__10712));
    CEMux I__1432 (
            .O(N__10724),
            .I(N__10712));
    CEMux I__1431 (
            .O(N__10723),
            .I(N__10712));
    GlobalMux I__1430 (
            .O(N__10712),
            .I(N__10709));
    gio2CtrlBuf I__1429 (
            .O(N__10709),
            .I(\delay_measurement_inst.delay_tr_timer.N_138_i_g ));
    InMux I__1428 (
            .O(N__10706),
            .I(N__10703));
    LocalMux I__1427 (
            .O(N__10703),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ));
    InMux I__1426 (
            .O(N__10700),
            .I(N__10697));
    LocalMux I__1425 (
            .O(N__10697),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ));
    InMux I__1424 (
            .O(N__10694),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__1423 (
            .O(N__10691),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__1422 (
            .O(N__10688),
            .I(bfn_4_17_0_));
    InMux I__1421 (
            .O(N__10685),
            .I(N__10682));
    LocalMux I__1420 (
            .O(N__10682),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__1419 (
            .O(N__10679),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__1418 (
            .O(N__10676),
            .I(N__10673));
    LocalMux I__1417 (
            .O(N__10673),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__1416 (
            .O(N__10670),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__1415 (
            .O(N__10667),
            .I(N__10664));
    LocalMux I__1414 (
            .O(N__10664),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__1413 (
            .O(N__10661),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__1412 (
            .O(N__10658),
            .I(N__10655));
    LocalMux I__1411 (
            .O(N__10655),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__1410 (
            .O(N__10652),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__1409 (
            .O(N__10649),
            .I(N__10646));
    LocalMux I__1408 (
            .O(N__10646),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__1407 (
            .O(N__10643),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__1406 (
            .O(N__10640),
            .I(N__10637));
    LocalMux I__1405 (
            .O(N__10637),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__1404 (
            .O(N__10634),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__1403 (
            .O(N__10631),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__1402 (
            .O(N__10628),
            .I(N__10625));
    LocalMux I__1401 (
            .O(N__10625),
            .I(N__10621));
    InMux I__1400 (
            .O(N__10624),
            .I(N__10618));
    Odrv12 I__1399 (
            .O(N__10621),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    LocalMux I__1398 (
            .O(N__10618),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    InMux I__1397 (
            .O(N__10613),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__1396 (
            .O(N__10610),
            .I(N__10606));
    InMux I__1395 (
            .O(N__10609),
            .I(N__10603));
    LocalMux I__1394 (
            .O(N__10606),
            .I(N__10600));
    LocalMux I__1393 (
            .O(N__10603),
            .I(N__10597));
    Odrv12 I__1392 (
            .O(N__10600),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    Odrv4 I__1391 (
            .O(N__10597),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    InMux I__1390 (
            .O(N__10592),
            .I(bfn_4_16_0_));
    InMux I__1389 (
            .O(N__10589),
            .I(N__10585));
    InMux I__1388 (
            .O(N__10588),
            .I(N__10582));
    LocalMux I__1387 (
            .O(N__10585),
            .I(N__10579));
    LocalMux I__1386 (
            .O(N__10582),
            .I(N__10576));
    Odrv12 I__1385 (
            .O(N__10579),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    Odrv4 I__1384 (
            .O(N__10576),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    InMux I__1383 (
            .O(N__10571),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__1382 (
            .O(N__10568),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__1381 (
            .O(N__10565),
            .I(N__10556));
    InMux I__1380 (
            .O(N__10564),
            .I(N__10556));
    InMux I__1379 (
            .O(N__10563),
            .I(N__10553));
    InMux I__1378 (
            .O(N__10562),
            .I(N__10550));
    InMux I__1377 (
            .O(N__10561),
            .I(N__10547));
    LocalMux I__1376 (
            .O(N__10556),
            .I(N__10544));
    LocalMux I__1375 (
            .O(N__10553),
            .I(N__10537));
    LocalMux I__1374 (
            .O(N__10550),
            .I(N__10537));
    LocalMux I__1373 (
            .O(N__10547),
            .I(N__10537));
    Odrv4 I__1372 (
            .O(N__10544),
            .I(\delay_measurement_inst.elapsed_time_tr_14 ));
    Odrv4 I__1371 (
            .O(N__10537),
            .I(\delay_measurement_inst.elapsed_time_tr_14 ));
    InMux I__1370 (
            .O(N__10532),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__1369 (
            .O(N__10529),
            .I(N__10525));
    CascadeMux I__1368 (
            .O(N__10528),
            .I(N__10521));
    InMux I__1367 (
            .O(N__10525),
            .I(N__10513));
    InMux I__1366 (
            .O(N__10524),
            .I(N__10513));
    InMux I__1365 (
            .O(N__10521),
            .I(N__10510));
    InMux I__1364 (
            .O(N__10520),
            .I(N__10505));
    InMux I__1363 (
            .O(N__10519),
            .I(N__10505));
    InMux I__1362 (
            .O(N__10518),
            .I(N__10502));
    LocalMux I__1361 (
            .O(N__10513),
            .I(N__10499));
    LocalMux I__1360 (
            .O(N__10510),
            .I(N__10492));
    LocalMux I__1359 (
            .O(N__10505),
            .I(N__10492));
    LocalMux I__1358 (
            .O(N__10502),
            .I(N__10492));
    Span4Mux_h I__1357 (
            .O(N__10499),
            .I(N__10489));
    Odrv4 I__1356 (
            .O(N__10492),
            .I(\delay_measurement_inst.elapsed_time_tr_15 ));
    Odrv4 I__1355 (
            .O(N__10489),
            .I(\delay_measurement_inst.elapsed_time_tr_15 ));
    InMux I__1354 (
            .O(N__10484),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__1353 (
            .O(N__10481),
            .I(N__10478));
    InMux I__1352 (
            .O(N__10478),
            .I(N__10473));
    InMux I__1351 (
            .O(N__10477),
            .I(N__10468));
    InMux I__1350 (
            .O(N__10476),
            .I(N__10468));
    LocalMux I__1349 (
            .O(N__10473),
            .I(N__10463));
    LocalMux I__1348 (
            .O(N__10468),
            .I(N__10463));
    Odrv4 I__1347 (
            .O(N__10463),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    InMux I__1346 (
            .O(N__10460),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__1345 (
            .O(N__10457),
            .I(N__10452));
    CascadeMux I__1344 (
            .O(N__10456),
            .I(N__10449));
    InMux I__1343 (
            .O(N__10455),
            .I(N__10443));
    InMux I__1342 (
            .O(N__10452),
            .I(N__10443));
    InMux I__1341 (
            .O(N__10449),
            .I(N__10440));
    InMux I__1340 (
            .O(N__10448),
            .I(N__10437));
    LocalMux I__1339 (
            .O(N__10443),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ));
    LocalMux I__1338 (
            .O(N__10440),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ));
    LocalMux I__1337 (
            .O(N__10437),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ));
    InMux I__1336 (
            .O(N__10430),
            .I(N__10427));
    LocalMux I__1335 (
            .O(N__10427),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_3 ));
    InMux I__1334 (
            .O(N__10424),
            .I(N__10420));
    InMux I__1333 (
            .O(N__10423),
            .I(N__10417));
    LocalMux I__1332 (
            .O(N__10420),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_2 ));
    LocalMux I__1331 (
            .O(N__10417),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_2 ));
    InMux I__1330 (
            .O(N__10412),
            .I(N__10408));
    CascadeMux I__1329 (
            .O(N__10411),
            .I(N__10405));
    LocalMux I__1328 (
            .O(N__10408),
            .I(N__10401));
    InMux I__1327 (
            .O(N__10405),
            .I(N__10398));
    InMux I__1326 (
            .O(N__10404),
            .I(N__10395));
    Odrv4 I__1325 (
            .O(N__10401),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    LocalMux I__1324 (
            .O(N__10398),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    LocalMux I__1323 (
            .O(N__10395),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    InMux I__1322 (
            .O(N__10388),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__1321 (
            .O(N__10385),
            .I(N__10382));
    LocalMux I__1320 (
            .O(N__10382),
            .I(N__10378));
    InMux I__1319 (
            .O(N__10381),
            .I(N__10375));
    Odrv4 I__1318 (
            .O(N__10378),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    LocalMux I__1317 (
            .O(N__10375),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    InMux I__1316 (
            .O(N__10370),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__1315 (
            .O(N__10367),
            .I(N__10364));
    InMux I__1314 (
            .O(N__10364),
            .I(N__10361));
    LocalMux I__1313 (
            .O(N__10361),
            .I(N__10357));
    CascadeMux I__1312 (
            .O(N__10360),
            .I(N__10354));
    Span4Mux_v I__1311 (
            .O(N__10357),
            .I(N__10350));
    InMux I__1310 (
            .O(N__10354),
            .I(N__10347));
    InMux I__1309 (
            .O(N__10353),
            .I(N__10344));
    Odrv4 I__1308 (
            .O(N__10350),
            .I(\delay_measurement_inst.elapsed_time_tr_6 ));
    LocalMux I__1307 (
            .O(N__10347),
            .I(\delay_measurement_inst.elapsed_time_tr_6 ));
    LocalMux I__1306 (
            .O(N__10344),
            .I(\delay_measurement_inst.elapsed_time_tr_6 ));
    InMux I__1305 (
            .O(N__10337),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__1304 (
            .O(N__10334),
            .I(N__10331));
    LocalMux I__1303 (
            .O(N__10331),
            .I(N__10326));
    InMux I__1302 (
            .O(N__10330),
            .I(N__10323));
    InMux I__1301 (
            .O(N__10329),
            .I(N__10320));
    Odrv4 I__1300 (
            .O(N__10326),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    LocalMux I__1299 (
            .O(N__10323),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    LocalMux I__1298 (
            .O(N__10320),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    InMux I__1297 (
            .O(N__10313),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__1296 (
            .O(N__10310),
            .I(N__10307));
    LocalMux I__1295 (
            .O(N__10307),
            .I(N__10304));
    Span4Mux_v I__1294 (
            .O(N__10304),
            .I(N__10299));
    InMux I__1293 (
            .O(N__10303),
            .I(N__10296));
    InMux I__1292 (
            .O(N__10302),
            .I(N__10293));
    Odrv4 I__1291 (
            .O(N__10299),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    LocalMux I__1290 (
            .O(N__10296),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    LocalMux I__1289 (
            .O(N__10293),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    InMux I__1288 (
            .O(N__10286),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__1287 (
            .O(N__10283),
            .I(N__10279));
    InMux I__1286 (
            .O(N__10282),
            .I(N__10274));
    InMux I__1285 (
            .O(N__10279),
            .I(N__10274));
    LocalMux I__1284 (
            .O(N__10274),
            .I(\delay_measurement_inst.N_200 ));
    InMux I__1283 (
            .O(N__10271),
            .I(N__10268));
    LocalMux I__1282 (
            .O(N__10268),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_3 ));
    CascadeMux I__1281 (
            .O(N__10265),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_ ));
    InMux I__1280 (
            .O(N__10262),
            .I(N__10259));
    LocalMux I__1279 (
            .O(N__10259),
            .I(\delay_measurement_inst.un1_tr_state_1_i_0_a2_0_7 ));
    InMux I__1278 (
            .O(N__10256),
            .I(N__10250));
    InMux I__1277 (
            .O(N__10255),
            .I(N__10250));
    LocalMux I__1276 (
            .O(N__10250),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10 ));
    CascadeMux I__1275 (
            .O(N__10247),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_ ));
    InMux I__1274 (
            .O(N__10244),
            .I(N__10241));
    LocalMux I__1273 (
            .O(N__10241),
            .I(\delay_measurement_inst.delay_tr_timer.N_203 ));
    InMux I__1272 (
            .O(N__10238),
            .I(N__10235));
    LocalMux I__1271 (
            .O(N__10235),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ));
    InMux I__1270 (
            .O(N__10232),
            .I(N__10228));
    InMux I__1269 (
            .O(N__10231),
            .I(N__10225));
    LocalMux I__1268 (
            .O(N__10228),
            .I(N__10222));
    LocalMux I__1267 (
            .O(N__10225),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__1266 (
            .O(N__10222),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__1265 (
            .O(N__10217),
            .I(N__10214));
    LocalMux I__1264 (
            .O(N__10214),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ));
    InMux I__1263 (
            .O(N__10211),
            .I(N__10207));
    InMux I__1262 (
            .O(N__10210),
            .I(N__10204));
    LocalMux I__1261 (
            .O(N__10207),
            .I(N__10201));
    LocalMux I__1260 (
            .O(N__10204),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__1259 (
            .O(N__10201),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__1258 (
            .O(N__10196),
            .I(N__10193));
    LocalMux I__1257 (
            .O(N__10193),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ));
    InMux I__1256 (
            .O(N__10190),
            .I(N__10186));
    InMux I__1255 (
            .O(N__10189),
            .I(N__10183));
    LocalMux I__1254 (
            .O(N__10186),
            .I(N__10180));
    LocalMux I__1253 (
            .O(N__10183),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__1252 (
            .O(N__10180),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__1251 (
            .O(N__10175),
            .I(N__10172));
    LocalMux I__1250 (
            .O(N__10172),
            .I(\delay_measurement_inst.N_168 ));
    InMux I__1249 (
            .O(N__10169),
            .I(N__10163));
    InMux I__1248 (
            .O(N__10168),
            .I(N__10163));
    LocalMux I__1247 (
            .O(N__10163),
            .I(\delay_measurement_inst.N_81_i ));
    CascadeMux I__1246 (
            .O(N__10160),
            .I(\delay_measurement_inst.N_81_i_cascade_ ));
    InMux I__1245 (
            .O(N__10157),
            .I(N__10153));
    InMux I__1244 (
            .O(N__10156),
            .I(N__10149));
    LocalMux I__1243 (
            .O(N__10153),
            .I(N__10146));
    InMux I__1242 (
            .O(N__10152),
            .I(N__10143));
    LocalMux I__1241 (
            .O(N__10149),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__1240 (
            .O(N__10146),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__1239 (
            .O(N__10143),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__1238 (
            .O(N__10136),
            .I(N__10133));
    LocalMux I__1237 (
            .O(N__10133),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ));
    CascadeMux I__1236 (
            .O(N__10130),
            .I(N__10127));
    InMux I__1235 (
            .O(N__10127),
            .I(N__10124));
    LocalMux I__1234 (
            .O(N__10124),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ));
    InMux I__1233 (
            .O(N__10121),
            .I(N__10118));
    LocalMux I__1232 (
            .O(N__10118),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ));
    InMux I__1231 (
            .O(N__10115),
            .I(N__10111));
    InMux I__1230 (
            .O(N__10114),
            .I(N__10108));
    LocalMux I__1229 (
            .O(N__10111),
            .I(N__10105));
    LocalMux I__1228 (
            .O(N__10108),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__1227 (
            .O(N__10105),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__1226 (
            .O(N__10100),
            .I(N__10097));
    LocalMux I__1225 (
            .O(N__10097),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ));
    InMux I__1224 (
            .O(N__10094),
            .I(N__10090));
    InMux I__1223 (
            .O(N__10093),
            .I(N__10087));
    LocalMux I__1222 (
            .O(N__10090),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__1221 (
            .O(N__10087),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__1220 (
            .O(N__10082),
            .I(N__10079));
    LocalMux I__1219 (
            .O(N__10079),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ));
    InMux I__1218 (
            .O(N__10076),
            .I(N__10072));
    InMux I__1217 (
            .O(N__10075),
            .I(N__10069));
    LocalMux I__1216 (
            .O(N__10072),
            .I(N__10066));
    LocalMux I__1215 (
            .O(N__10069),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__1214 (
            .O(N__10066),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__1213 (
            .O(N__10061),
            .I(N__10058));
    LocalMux I__1212 (
            .O(N__10058),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ));
    InMux I__1211 (
            .O(N__10055),
            .I(N__10051));
    InMux I__1210 (
            .O(N__10054),
            .I(N__10048));
    LocalMux I__1209 (
            .O(N__10051),
            .I(N__10045));
    LocalMux I__1208 (
            .O(N__10048),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__1207 (
            .O(N__10045),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__1206 (
            .O(N__10040),
            .I(N__10037));
    LocalMux I__1205 (
            .O(N__10037),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ));
    InMux I__1204 (
            .O(N__10034),
            .I(N__10030));
    InMux I__1203 (
            .O(N__10033),
            .I(N__10027));
    LocalMux I__1202 (
            .O(N__10030),
            .I(N__10024));
    LocalMux I__1201 (
            .O(N__10027),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__1200 (
            .O(N__10024),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__1199 (
            .O(N__10019),
            .I(N__10016));
    LocalMux I__1198 (
            .O(N__10016),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ));
    InMux I__1197 (
            .O(N__10013),
            .I(N__10009));
    InMux I__1196 (
            .O(N__10012),
            .I(N__10006));
    LocalMux I__1195 (
            .O(N__10009),
            .I(N__10003));
    LocalMux I__1194 (
            .O(N__10006),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__1193 (
            .O(N__10003),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ));
    CascadeMux I__1192 (
            .O(N__9998),
            .I(N__9995));
    InMux I__1191 (
            .O(N__9995),
            .I(N__9992));
    LocalMux I__1190 (
            .O(N__9992),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__1189 (
            .O(N__9989),
            .I(N__9986));
    InMux I__1188 (
            .O(N__9986),
            .I(N__9983));
    LocalMux I__1187 (
            .O(N__9983),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__1186 (
            .O(N__9980),
            .I(N__9977));
    InMux I__1185 (
            .O(N__9977),
            .I(N__9974));
    LocalMux I__1184 (
            .O(N__9974),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ));
    CascadeMux I__1183 (
            .O(N__9971),
            .I(N__9968));
    InMux I__1182 (
            .O(N__9968),
            .I(N__9965));
    LocalMux I__1181 (
            .O(N__9965),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ));
    CascadeMux I__1180 (
            .O(N__9962),
            .I(N__9959));
    InMux I__1179 (
            .O(N__9959),
            .I(N__9956));
    LocalMux I__1178 (
            .O(N__9956),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ));
    CascadeMux I__1177 (
            .O(N__9953),
            .I(N__9950));
    InMux I__1176 (
            .O(N__9950),
            .I(N__9947));
    LocalMux I__1175 (
            .O(N__9947),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ));
    CascadeMux I__1174 (
            .O(N__9944),
            .I(N__9941));
    InMux I__1173 (
            .O(N__9941),
            .I(N__9938));
    LocalMux I__1172 (
            .O(N__9938),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ));
    InMux I__1171 (
            .O(N__9935),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__1170 (
            .O(N__9932),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ));
    CascadeMux I__1169 (
            .O(N__9929),
            .I(N__9926));
    InMux I__1168 (
            .O(N__9926),
            .I(N__9923));
    LocalMux I__1167 (
            .O(N__9923),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ));
    InMux I__1166 (
            .O(N__9920),
            .I(N__9917));
    LocalMux I__1165 (
            .O(N__9917),
            .I(N__9913));
    InMux I__1164 (
            .O(N__9916),
            .I(N__9910));
    Odrv4 I__1163 (
            .O(N__9913),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__1162 (
            .O(N__9910),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__1161 (
            .O(N__9905),
            .I(N__9902));
    InMux I__1160 (
            .O(N__9902),
            .I(N__9899));
    LocalMux I__1159 (
            .O(N__9899),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ));
    InMux I__1158 (
            .O(N__9896),
            .I(N__9892));
    InMux I__1157 (
            .O(N__9895),
            .I(N__9889));
    LocalMux I__1156 (
            .O(N__9892),
            .I(N__9886));
    LocalMux I__1155 (
            .O(N__9889),
            .I(N__9883));
    Odrv12 I__1154 (
            .O(N__9886),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv4 I__1153 (
            .O(N__9883),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__1152 (
            .O(N__9878),
            .I(N__9875));
    InMux I__1151 (
            .O(N__9875),
            .I(N__9872));
    LocalMux I__1150 (
            .O(N__9872),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ));
    InMux I__1149 (
            .O(N__9869),
            .I(N__9866));
    LocalMux I__1148 (
            .O(N__9866),
            .I(N__9862));
    InMux I__1147 (
            .O(N__9865),
            .I(N__9859));
    Odrv12 I__1146 (
            .O(N__9862),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__1145 (
            .O(N__9859),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__1144 (
            .O(N__9854),
            .I(N__9851));
    InMux I__1143 (
            .O(N__9851),
            .I(N__9848));
    LocalMux I__1142 (
            .O(N__9848),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ));
    CascadeMux I__1141 (
            .O(N__9845),
            .I(N__9842));
    InMux I__1140 (
            .O(N__9842),
            .I(N__9838));
    InMux I__1139 (
            .O(N__9841),
            .I(N__9835));
    LocalMux I__1138 (
            .O(N__9838),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__1137 (
            .O(N__9835),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__1136 (
            .O(N__9830),
            .I(N__9827));
    InMux I__1135 (
            .O(N__9827),
            .I(N__9824));
    LocalMux I__1134 (
            .O(N__9824),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ));
    InMux I__1133 (
            .O(N__9821),
            .I(N__9818));
    LocalMux I__1132 (
            .O(N__9818),
            .I(N__9814));
    InMux I__1131 (
            .O(N__9817),
            .I(N__9811));
    Odrv4 I__1130 (
            .O(N__9814),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__1129 (
            .O(N__9811),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__1128 (
            .O(N__9806),
            .I(N__9803));
    InMux I__1127 (
            .O(N__9803),
            .I(N__9800));
    LocalMux I__1126 (
            .O(N__9800),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ));
    InMux I__1125 (
            .O(N__9797),
            .I(N__9794));
    LocalMux I__1124 (
            .O(N__9794),
            .I(N__9790));
    InMux I__1123 (
            .O(N__9793),
            .I(N__9787));
    Odrv4 I__1122 (
            .O(N__9790),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__1121 (
            .O(N__9787),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__1120 (
            .O(N__9782),
            .I(N__9779));
    InMux I__1119 (
            .O(N__9779),
            .I(N__9776));
    LocalMux I__1118 (
            .O(N__9776),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__1117 (
            .O(N__9773),
            .I(N__9770));
    InMux I__1116 (
            .O(N__9770),
            .I(N__9767));
    LocalMux I__1115 (
            .O(N__9767),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__1114 (
            .O(N__9764),
            .I(N__9761));
    InMux I__1113 (
            .O(N__9761),
            .I(N__9758));
    LocalMux I__1112 (
            .O(N__9758),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__1111 (
            .O(N__9755),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19_cascade_ ));
    InMux I__1110 (
            .O(N__9752),
            .I(N__9749));
    LocalMux I__1109 (
            .O(N__9749),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19 ));
    InMux I__1108 (
            .O(N__9746),
            .I(N__9743));
    LocalMux I__1107 (
            .O(N__9743),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19 ));
    CascadeMux I__1106 (
            .O(N__9740),
            .I(N__9737));
    InMux I__1105 (
            .O(N__9737),
            .I(N__9734));
    LocalMux I__1104 (
            .O(N__9734),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ));
    InMux I__1103 (
            .O(N__9731),
            .I(N__9728));
    LocalMux I__1102 (
            .O(N__9728),
            .I(N__9724));
    InMux I__1101 (
            .O(N__9727),
            .I(N__9721));
    Odrv12 I__1100 (
            .O(N__9724),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__1099 (
            .O(N__9721),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__1098 (
            .O(N__9716),
            .I(N__9713));
    InMux I__1097 (
            .O(N__9713),
            .I(N__9710));
    LocalMux I__1096 (
            .O(N__9710),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ));
    InMux I__1095 (
            .O(N__9707),
            .I(N__9704));
    LocalMux I__1094 (
            .O(N__9704),
            .I(N__9700));
    InMux I__1093 (
            .O(N__9703),
            .I(N__9697));
    Odrv4 I__1092 (
            .O(N__9700),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__1091 (
            .O(N__9697),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__1090 (
            .O(N__9692),
            .I(N__9689));
    InMux I__1089 (
            .O(N__9689),
            .I(N__9686));
    LocalMux I__1088 (
            .O(N__9686),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ));
    InMux I__1087 (
            .O(N__9683),
            .I(N__9680));
    LocalMux I__1086 (
            .O(N__9680),
            .I(N__9676));
    InMux I__1085 (
            .O(N__9679),
            .I(N__9673));
    Odrv12 I__1084 (
            .O(N__9676),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__1083 (
            .O(N__9673),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__1082 (
            .O(N__9668),
            .I(N__9665));
    InMux I__1081 (
            .O(N__9665),
            .I(N__9662));
    LocalMux I__1080 (
            .O(N__9662),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ));
    InMux I__1079 (
            .O(N__9659),
            .I(N__9656));
    LocalMux I__1078 (
            .O(N__9656),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ));
    InMux I__1077 (
            .O(N__9653),
            .I(N__9650));
    LocalMux I__1076 (
            .O(N__9650),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ));
    InMux I__1075 (
            .O(N__9647),
            .I(N__9644));
    LocalMux I__1074 (
            .O(N__9644),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ));
    InMux I__1073 (
            .O(N__9641),
            .I(N__9638));
    LocalMux I__1072 (
            .O(N__9638),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ));
    InMux I__1071 (
            .O(N__9635),
            .I(N__9632));
    LocalMux I__1070 (
            .O(N__9632),
            .I(N__9629));
    Odrv4 I__1069 (
            .O(N__9629),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ));
    InMux I__1068 (
            .O(N__9626),
            .I(N__9623));
    LocalMux I__1067 (
            .O(N__9623),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ));
    InMux I__1066 (
            .O(N__9620),
            .I(N__9617));
    LocalMux I__1065 (
            .O(N__9617),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ));
    InMux I__1064 (
            .O(N__9614),
            .I(N__9611));
    LocalMux I__1063 (
            .O(N__9611),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__1062 (
            .O(N__9608),
            .I(N__9605));
    InMux I__1061 (
            .O(N__9605),
            .I(N__9601));
    InMux I__1060 (
            .O(N__9604),
            .I(N__9598));
    LocalMux I__1059 (
            .O(N__9601),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    LocalMux I__1058 (
            .O(N__9598),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    InMux I__1057 (
            .O(N__9593),
            .I(N__9586));
    InMux I__1056 (
            .O(N__9592),
            .I(N__9586));
    InMux I__1055 (
            .O(N__9591),
            .I(N__9583));
    LocalMux I__1054 (
            .O(N__9586),
            .I(N__9580));
    LocalMux I__1053 (
            .O(N__9583),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    Odrv4 I__1052 (
            .O(N__9580),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    InMux I__1051 (
            .O(N__9575),
            .I(N__9572));
    LocalMux I__1050 (
            .O(N__9572),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6 ));
    CascadeMux I__1049 (
            .O(N__9569),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5_cascade_ ));
    InMux I__1048 (
            .O(N__9566),
            .I(N__9563));
    LocalMux I__1047 (
            .O(N__9563),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ));
    InMux I__1046 (
            .O(N__9560),
            .I(N__9557));
    LocalMux I__1045 (
            .O(N__9557),
            .I(N__9554));
    Odrv4 I__1044 (
            .O(N__9554),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ));
    InMux I__1043 (
            .O(N__9551),
            .I(N__9548));
    LocalMux I__1042 (
            .O(N__9548),
            .I(N__9545));
    Odrv4 I__1041 (
            .O(N__9545),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ));
    InMux I__1040 (
            .O(N__9542),
            .I(N__9539));
    LocalMux I__1039 (
            .O(N__9539),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ));
    InMux I__1038 (
            .O(N__9536),
            .I(N__9533));
    LocalMux I__1037 (
            .O(N__9533),
            .I(N__9530));
    Odrv4 I__1036 (
            .O(N__9530),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__1035 (
            .O(N__9527),
            .I(\delay_measurement_inst.N_212_cascade_ ));
    InMux I__1034 (
            .O(N__9524),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__1033 (
            .O(N__9521),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__1032 (
            .O(N__9518),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__1031 (
            .O(N__9515),
            .I(bfn_2_24_0_));
    InMux I__1030 (
            .O(N__9512),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__1029 (
            .O(N__9509),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__1028 (
            .O(N__9506),
            .I(N__9503));
    LocalMux I__1027 (
            .O(N__9503),
            .I(N__9500));
    Odrv4 I__1026 (
            .O(N__9500),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ));
    InMux I__1025 (
            .O(N__9497),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__1024 (
            .O(N__9494),
            .I(N__9491));
    LocalMux I__1023 (
            .O(N__9491),
            .I(N__9488));
    Odrv4 I__1022 (
            .O(N__9488),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ));
    InMux I__1021 (
            .O(N__9485),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__1020 (
            .O(N__9482),
            .I(N__9479));
    LocalMux I__1019 (
            .O(N__9479),
            .I(N__9476));
    Odrv4 I__1018 (
            .O(N__9476),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ));
    InMux I__1017 (
            .O(N__9473),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ));
    CascadeMux I__1016 (
            .O(N__9470),
            .I(N__9467));
    InMux I__1015 (
            .O(N__9467),
            .I(N__9464));
    LocalMux I__1014 (
            .O(N__9464),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ));
    InMux I__1013 (
            .O(N__9461),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__1012 (
            .O(N__9458),
            .I(N__9455));
    LocalMux I__1011 (
            .O(N__9455),
            .I(N__9452));
    Odrv4 I__1010 (
            .O(N__9452),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ));
    InMux I__1009 (
            .O(N__9449),
            .I(bfn_2_23_0_));
    CascadeMux I__1008 (
            .O(N__9446),
            .I(N__9443));
    InMux I__1007 (
            .O(N__9443),
            .I(N__9440));
    LocalMux I__1006 (
            .O(N__9440),
            .I(N__9437));
    Odrv4 I__1005 (
            .O(N__9437),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ));
    InMux I__1004 (
            .O(N__9434),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__1003 (
            .O(N__9431),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__1002 (
            .O(N__9428),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__1001 (
            .O(N__9425),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__1000 (
            .O(N__9422),
            .I(N__9419));
    LocalMux I__999 (
            .O(N__9419),
            .I(N__9416));
    Odrv4 I__998 (
            .O(N__9416),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ));
    InMux I__997 (
            .O(N__9413),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__996 (
            .O(N__9410),
            .I(N__9407));
    LocalMux I__995 (
            .O(N__9407),
            .I(N__9404));
    Odrv4 I__994 (
            .O(N__9404),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ));
    InMux I__993 (
            .O(N__9401),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__992 (
            .O(N__9398),
            .I(N__9395));
    LocalMux I__991 (
            .O(N__9395),
            .I(N__9392));
    Odrv4 I__990 (
            .O(N__9392),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ));
    InMux I__989 (
            .O(N__9389),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__988 (
            .O(N__9386),
            .I(N__9383));
    LocalMux I__987 (
            .O(N__9383),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ));
    InMux I__986 (
            .O(N__9380),
            .I(N__9376));
    InMux I__985 (
            .O(N__9379),
            .I(N__9373));
    LocalMux I__984 (
            .O(N__9376),
            .I(N__9370));
    LocalMux I__983 (
            .O(N__9373),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__982 (
            .O(N__9370),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__981 (
            .O(N__9365),
            .I(N__9362));
    InMux I__980 (
            .O(N__9362),
            .I(N__9359));
    LocalMux I__979 (
            .O(N__9359),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ));
    InMux I__978 (
            .O(N__9356),
            .I(N__9352));
    InMux I__977 (
            .O(N__9355),
            .I(N__9349));
    LocalMux I__976 (
            .O(N__9352),
            .I(N__9346));
    LocalMux I__975 (
            .O(N__9349),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__974 (
            .O(N__9346),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__973 (
            .O(N__9341),
            .I(N__9338));
    LocalMux I__972 (
            .O(N__9338),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ));
    InMux I__971 (
            .O(N__9335),
            .I(N__9331));
    InMux I__970 (
            .O(N__9334),
            .I(N__9328));
    LocalMux I__969 (
            .O(N__9331),
            .I(N__9325));
    LocalMux I__968 (
            .O(N__9328),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__967 (
            .O(N__9325),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__966 (
            .O(N__9320),
            .I(N__9317));
    LocalMux I__965 (
            .O(N__9317),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ));
    InMux I__964 (
            .O(N__9314),
            .I(N__9310));
    InMux I__963 (
            .O(N__9313),
            .I(N__9307));
    LocalMux I__962 (
            .O(N__9310),
            .I(N__9304));
    LocalMux I__961 (
            .O(N__9307),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__960 (
            .O(N__9304),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    CascadeMux I__959 (
            .O(N__9299),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_ ));
    InMux I__958 (
            .O(N__9296),
            .I(N__9293));
    LocalMux I__957 (
            .O(N__9293),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ));
    InMux I__956 (
            .O(N__9290),
            .I(N__9287));
    LocalMux I__955 (
            .O(N__9287),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ));
    InMux I__954 (
            .O(N__9284),
            .I(N__9280));
    InMux I__953 (
            .O(N__9283),
            .I(N__9277));
    LocalMux I__952 (
            .O(N__9280),
            .I(N__9274));
    LocalMux I__951 (
            .O(N__9277),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__950 (
            .O(N__9274),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__949 (
            .O(N__9269),
            .I(N__9266));
    LocalMux I__948 (
            .O(N__9266),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ));
    InMux I__947 (
            .O(N__9263),
            .I(N__9259));
    InMux I__946 (
            .O(N__9262),
            .I(N__9256));
    LocalMux I__945 (
            .O(N__9259),
            .I(N__9253));
    LocalMux I__944 (
            .O(N__9256),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__943 (
            .O(N__9253),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    CascadeMux I__942 (
            .O(N__9248),
            .I(N__9245));
    InMux I__941 (
            .O(N__9245),
            .I(N__9242));
    LocalMux I__940 (
            .O(N__9242),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ));
    InMux I__939 (
            .O(N__9239),
            .I(N__9235));
    InMux I__938 (
            .O(N__9238),
            .I(N__9232));
    LocalMux I__937 (
            .O(N__9235),
            .I(N__9229));
    LocalMux I__936 (
            .O(N__9232),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__935 (
            .O(N__9229),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__934 (
            .O(N__9224),
            .I(N__9221));
    LocalMux I__933 (
            .O(N__9221),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ));
    InMux I__932 (
            .O(N__9218),
            .I(N__9214));
    InMux I__931 (
            .O(N__9217),
            .I(N__9211));
    LocalMux I__930 (
            .O(N__9214),
            .I(N__9208));
    LocalMux I__929 (
            .O(N__9211),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__928 (
            .O(N__9208),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    CascadeMux I__927 (
            .O(N__9203),
            .I(N__9200));
    InMux I__926 (
            .O(N__9200),
            .I(N__9197));
    LocalMux I__925 (
            .O(N__9197),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ));
    InMux I__924 (
            .O(N__9194),
            .I(N__9190));
    InMux I__923 (
            .O(N__9193),
            .I(N__9187));
    LocalMux I__922 (
            .O(N__9190),
            .I(N__9184));
    LocalMux I__921 (
            .O(N__9187),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__920 (
            .O(N__9184),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__919 (
            .O(N__9179),
            .I(N__9176));
    LocalMux I__918 (
            .O(N__9176),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ));
    InMux I__917 (
            .O(N__9173),
            .I(N__9169));
    InMux I__916 (
            .O(N__9172),
            .I(N__9166));
    LocalMux I__915 (
            .O(N__9169),
            .I(N__9163));
    LocalMux I__914 (
            .O(N__9166),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__913 (
            .O(N__9163),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ));
    CascadeMux I__912 (
            .O(N__9158),
            .I(N__9155));
    InMux I__911 (
            .O(N__9155),
            .I(N__9152));
    LocalMux I__910 (
            .O(N__9152),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ));
    InMux I__909 (
            .O(N__9149),
            .I(N__9145));
    InMux I__908 (
            .O(N__9148),
            .I(N__9142));
    LocalMux I__907 (
            .O(N__9145),
            .I(N__9139));
    LocalMux I__906 (
            .O(N__9142),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__905 (
            .O(N__9139),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    CascadeMux I__904 (
            .O(N__9134),
            .I(N__9131));
    InMux I__903 (
            .O(N__9131),
            .I(N__9128));
    LocalMux I__902 (
            .O(N__9128),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__901 (
            .O(N__9125),
            .I(N__9122));
    InMux I__900 (
            .O(N__9122),
            .I(N__9119));
    LocalMux I__899 (
            .O(N__9119),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__898 (
            .O(N__9116),
            .I(N__9113));
    InMux I__897 (
            .O(N__9113),
            .I(N__9110));
    LocalMux I__896 (
            .O(N__9110),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__895 (
            .O(N__9107),
            .I(N__9104));
    InMux I__894 (
            .O(N__9104),
            .I(N__9101));
    LocalMux I__893 (
            .O(N__9101),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ));
    CascadeMux I__892 (
            .O(N__9098),
            .I(N__9095));
    InMux I__891 (
            .O(N__9095),
            .I(N__9092));
    LocalMux I__890 (
            .O(N__9092),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ));
    CascadeMux I__889 (
            .O(N__9089),
            .I(N__9086));
    InMux I__888 (
            .O(N__9086),
            .I(N__9083));
    LocalMux I__887 (
            .O(N__9083),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ));
    CascadeMux I__886 (
            .O(N__9080),
            .I(N__9077));
    InMux I__885 (
            .O(N__9077),
            .I(N__9074));
    LocalMux I__884 (
            .O(N__9074),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ));
    InMux I__883 (
            .O(N__9071),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__882 (
            .O(N__9068),
            .I(N__9065));
    LocalMux I__881 (
            .O(N__9065),
            .I(N__9062));
    Odrv4 I__880 (
            .O(N__9062),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ));
    InMux I__879 (
            .O(N__9059),
            .I(N__9056));
    LocalMux I__878 (
            .O(N__9056),
            .I(N__9052));
    InMux I__877 (
            .O(N__9055),
            .I(N__9049));
    Odrv4 I__876 (
            .O(N__9052),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__875 (
            .O(N__9049),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    CascadeMux I__874 (
            .O(N__9044),
            .I(N__9041));
    InMux I__873 (
            .O(N__9041),
            .I(N__9038));
    LocalMux I__872 (
            .O(N__9038),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ));
    InMux I__871 (
            .O(N__9035),
            .I(N__9032));
    LocalMux I__870 (
            .O(N__9032),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_6 ));
    InMux I__869 (
            .O(N__9029),
            .I(N__9026));
    LocalMux I__868 (
            .O(N__9026),
            .I(N__9022));
    InMux I__867 (
            .O(N__9025),
            .I(N__9019));
    Odrv4 I__866 (
            .O(N__9022),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__865 (
            .O(N__9019),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ));
    CascadeMux I__864 (
            .O(N__9014),
            .I(N__9011));
    InMux I__863 (
            .O(N__9011),
            .I(N__9008));
    LocalMux I__862 (
            .O(N__9008),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ));
    InMux I__861 (
            .O(N__9005),
            .I(N__9002));
    LocalMux I__860 (
            .O(N__9002),
            .I(N__8998));
    InMux I__859 (
            .O(N__9001),
            .I(N__8995));
    Odrv4 I__858 (
            .O(N__8998),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__857 (
            .O(N__8995),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    CascadeMux I__856 (
            .O(N__8990),
            .I(N__8987));
    InMux I__855 (
            .O(N__8987),
            .I(N__8984));
    LocalMux I__854 (
            .O(N__8984),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ));
    InMux I__853 (
            .O(N__8981),
            .I(N__8978));
    LocalMux I__852 (
            .O(N__8978),
            .I(N__8974));
    InMux I__851 (
            .O(N__8977),
            .I(N__8971));
    Odrv12 I__850 (
            .O(N__8974),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__849 (
            .O(N__8971),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ));
    CascadeMux I__848 (
            .O(N__8966),
            .I(N__8963));
    InMux I__847 (
            .O(N__8963),
            .I(N__8960));
    LocalMux I__846 (
            .O(N__8960),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ));
    CascadeMux I__845 (
            .O(N__8957),
            .I(N__8954));
    InMux I__844 (
            .O(N__8954),
            .I(N__8951));
    LocalMux I__843 (
            .O(N__8951),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__842 (
            .O(N__8948),
            .I(N__8945));
    InMux I__841 (
            .O(N__8945),
            .I(N__8942));
    LocalMux I__840 (
            .O(N__8942),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__839 (
            .O(N__8939),
            .I(N__8936));
    InMux I__838 (
            .O(N__8936),
            .I(N__8933));
    LocalMux I__837 (
            .O(N__8933),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__836 (
            .O(N__8930),
            .I(N__8927));
    InMux I__835 (
            .O(N__8927),
            .I(N__8924));
    LocalMux I__834 (
            .O(N__8924),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ));
    InMux I__833 (
            .O(N__8921),
            .I(N__8918));
    LocalMux I__832 (
            .O(N__8918),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__831 (
            .O(N__8915),
            .I(N__8912));
    InMux I__830 (
            .O(N__8912),
            .I(N__8908));
    InMux I__829 (
            .O(N__8911),
            .I(N__8904));
    LocalMux I__828 (
            .O(N__8908),
            .I(N__8901));
    InMux I__827 (
            .O(N__8907),
            .I(N__8898));
    LocalMux I__826 (
            .O(N__8904),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv12 I__825 (
            .O(N__8901),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__824 (
            .O(N__8898),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__823 (
            .O(N__8891),
            .I(N__8888));
    InMux I__822 (
            .O(N__8888),
            .I(N__8885));
    LocalMux I__821 (
            .O(N__8885),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ));
    InMux I__820 (
            .O(N__8882),
            .I(N__8879));
    LocalMux I__819 (
            .O(N__8879),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ));
    InMux I__818 (
            .O(N__8876),
            .I(N__8873));
    LocalMux I__817 (
            .O(N__8873),
            .I(N__8869));
    InMux I__816 (
            .O(N__8872),
            .I(N__8866));
    Odrv4 I__815 (
            .O(N__8869),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__814 (
            .O(N__8866),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    CascadeMux I__813 (
            .O(N__8861),
            .I(N__8858));
    InMux I__812 (
            .O(N__8858),
            .I(N__8855));
    LocalMux I__811 (
            .O(N__8855),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ));
    InMux I__810 (
            .O(N__8852),
            .I(N__8849));
    LocalMux I__809 (
            .O(N__8849),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ));
    InMux I__808 (
            .O(N__8846),
            .I(N__8843));
    LocalMux I__807 (
            .O(N__8843),
            .I(N__8839));
    InMux I__806 (
            .O(N__8842),
            .I(N__8836));
    Odrv4 I__805 (
            .O(N__8839),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__804 (
            .O(N__8836),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__803 (
            .O(N__8831),
            .I(N__8828));
    InMux I__802 (
            .O(N__8828),
            .I(N__8825));
    LocalMux I__801 (
            .O(N__8825),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ));
    InMux I__800 (
            .O(N__8822),
            .I(N__8819));
    LocalMux I__799 (
            .O(N__8819),
            .I(N__8816));
    Odrv4 I__798 (
            .O(N__8816),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ));
    InMux I__797 (
            .O(N__8813),
            .I(N__8810));
    LocalMux I__796 (
            .O(N__8810),
            .I(N__8806));
    InMux I__795 (
            .O(N__8809),
            .I(N__8803));
    Odrv4 I__794 (
            .O(N__8806),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__793 (
            .O(N__8803),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    CascadeMux I__792 (
            .O(N__8798),
            .I(N__8795));
    InMux I__791 (
            .O(N__8795),
            .I(N__8792));
    LocalMux I__790 (
            .O(N__8792),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ));
    InMux I__789 (
            .O(N__8789),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__788 (
            .O(N__8786),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__787 (
            .O(N__8783),
            .I(N__8780));
    LocalMux I__786 (
            .O(N__8780),
            .I(N_27_i_i));
    InMux I__785 (
            .O(N__8777),
            .I(N__8774));
    LocalMux I__784 (
            .O(N__8774),
            .I(un7_start_stop));
    InMux I__783 (
            .O(N__8771),
            .I(N__8768));
    LocalMux I__782 (
            .O(N__8768),
            .I(N__8765));
    Span12Mux_s5_v I__781 (
            .O(N__8765),
            .I(N__8762));
    Span12Mux_h I__780 (
            .O(N__8762),
            .I(N__8759));
    Span12Mux_h I__779 (
            .O(N__8759),
            .I(N__8753));
    InMux I__778 (
            .O(N__8758),
            .I(N__8750));
    InMux I__777 (
            .O(N__8757),
            .I(N__8747));
    InMux I__776 (
            .O(N__8756),
            .I(N__8744));
    Odrv12 I__775 (
            .O(N__8753),
            .I(CONSTANT_ONE_NET));
    LocalMux I__774 (
            .O(N__8750),
            .I(CONSTANT_ONE_NET));
    LocalMux I__773 (
            .O(N__8747),
            .I(CONSTANT_ONE_NET));
    LocalMux I__772 (
            .O(N__8744),
            .I(CONSTANT_ONE_NET));
    InMux I__771 (
            .O(N__8735),
            .I(bfn_1_19_0_));
    InMux I__770 (
            .O(N__8732),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__769 (
            .O(N__8729),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__768 (
            .O(N__8726),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__767 (
            .O(N__8723),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__766 (
            .O(N__8720),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__765 (
            .O(N__8717),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__764 (
            .O(N__8714),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__763 (
            .O(N__8711),
            .I(bfn_1_20_0_));
    InMux I__762 (
            .O(N__8708),
            .I(N__8705));
    LocalMux I__761 (
            .O(N__8705),
            .I(N__8702));
    Odrv4 I__760 (
            .O(N__8702),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ));
    InMux I__759 (
            .O(N__8699),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ));
    CascadeMux I__758 (
            .O(N__8696),
            .I(N__8693));
    InMux I__757 (
            .O(N__8693),
            .I(N__8690));
    LocalMux I__756 (
            .O(N__8690),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ));
    InMux I__755 (
            .O(N__8687),
            .I(N__8684));
    LocalMux I__754 (
            .O(N__8684),
            .I(N__8681));
    Odrv4 I__753 (
            .O(N__8681),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ));
    InMux I__752 (
            .O(N__8678),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__751 (
            .O(N__8675),
            .I(N__8672));
    LocalMux I__750 (
            .O(N__8672),
            .I(N__8669));
    Odrv4 I__749 (
            .O(N__8669),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ));
    InMux I__748 (
            .O(N__8666),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__747 (
            .O(N__8663),
            .I(N__8660));
    LocalMux I__746 (
            .O(N__8660),
            .I(N__8657));
    Odrv4 I__745 (
            .O(N__8657),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ));
    InMux I__744 (
            .O(N__8654),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__743 (
            .O(N__8651),
            .I(N__8648));
    LocalMux I__742 (
            .O(N__8648),
            .I(N__8645));
    Odrv4 I__741 (
            .O(N__8645),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ));
    InMux I__740 (
            .O(N__8642),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__739 (
            .O(N__8639),
            .I(N__8636));
    LocalMux I__738 (
            .O(N__8636),
            .I(N__8633));
    Odrv4 I__737 (
            .O(N__8633),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ));
    InMux I__736 (
            .O(N__8630),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__735 (
            .O(N__8627),
            .I(N__8624));
    LocalMux I__734 (
            .O(N__8624),
            .I(N__8621));
    Odrv4 I__733 (
            .O(N__8621),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ));
    InMux I__732 (
            .O(N__8618),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__731 (
            .O(N__8615),
            .I(N__8612));
    LocalMux I__730 (
            .O(N__8612),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0 ));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_1_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_20_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_1_20_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_3_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_20_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_3_20_0_));
    defparam IN_MUX_bfv_3_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_21_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_3_21_0_));
    defparam IN_MUX_bfv_2_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_22_0_));
    defparam IN_MUX_bfv_2_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_23_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_2_23_0_));
    defparam IN_MUX_bfv_2_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_24_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_2_24_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_7_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_21_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_7_21_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_4_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_15_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_4_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_17_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_4_17_0_));
    defparam IN_MUX_bfv_4_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_18_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_4_18_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_5_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_5_16_0_));
    defparam IN_MUX_bfv_5_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_17_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_5_17_0_));
    defparam IN_MUX_bfv_5_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_18_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_5_18_0_));
    defparam IN_MUX_bfv_8_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_26_0_));
    defparam IN_MUX_bfv_8_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_27_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_8_27_0_));
    defparam IN_MUX_bfv_8_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_28_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_8_28_0_));
    defparam IN_MUX_bfv_8_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_29_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_8_29_0_));
    defparam IN_MUX_bfv_9_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_26_0_));
    defparam IN_MUX_bfv_9_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_27_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_9_27_0_));
    defparam IN_MUX_bfv_9_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_28_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_9_28_0_));
    defparam IN_MUX_bfv_9_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_29_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_9_29_0_));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0  (
            .USERSIGNALTOGLOBALBUFFER(N__19511),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_138_i_g ));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__21734),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_136_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__8756),
            .CLKHFEN(N__8758),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__8757),
            .RGB2PWM(N__8783),
            .RGB1(rgb_g),
            .CURREN(N__8771),
            .RGB2(rgb_b),
            .RGB1PWM(N__8777),
            .RGB0PWM(N__22342),
            .RGB0(rgb_r));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_0  (
            .USERSIGNALTOGLOBALBUFFER(N__21458),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_139_i_g ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_1_14_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_1_14_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_1_14_2 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_0_LC_1_14_2  (
            .in0(N__15111),
            .in1(N__15069),
            .in2(N__19907),
            .in3(N__15170),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22041),
            .ce(N__21315),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_1_16_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_1_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_1_16_0 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_8_LC_1_16_0  (
            .in0(N__15064),
            .in1(N__19860),
            .in2(N__15262),
            .in3(N__8627),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22036),
            .ce(),
            .sr(N__22278));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_1_16_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_1_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_1_16_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_1_LC_1_16_1  (
            .in0(N__15254),
            .in1(N__15065),
            .in2(N__19898),
            .in3(N__8615),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22036),
            .ce(),
            .sr(N__22278));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_1_16_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_1_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_1_16_2 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_5_LC_1_16_2  (
            .in0(N__15062),
            .in1(N__19858),
            .in2(N__15260),
            .in3(N__8663),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22036),
            .ce(),
            .sr(N__22278));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_1_16_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_1_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_1_16_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_7_LC_1_16_3  (
            .in0(N__15257),
            .in1(N__15068),
            .in2(N__19901),
            .in3(N__8639),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22036),
            .ce(),
            .sr(N__22278));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_1_16_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_1_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_1_16_4 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_3_LC_1_16_4  (
            .in0(N__15061),
            .in1(N__19857),
            .in2(N__15259),
            .in3(N__8687),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22036),
            .ce(),
            .sr(N__22278));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_1_16_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_1_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_1_16_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_2_LC_1_16_5  (
            .in0(N__15255),
            .in1(N__15066),
            .in2(N__19899),
            .in3(N__8708),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22036),
            .ce(),
            .sr(N__22278));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_1_16_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_1_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_1_16_6 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_6_LC_1_16_6  (
            .in0(N__15063),
            .in1(N__19859),
            .in2(N__15261),
            .in3(N__8651),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22036),
            .ce(),
            .sr(N__22278));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_1_16_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_1_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_1_16_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_4_LC_1_16_7  (
            .in0(N__15256),
            .in1(N__15067),
            .in2(N__19900),
            .in3(N__8675),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22036),
            .ce(),
            .sr(N__22278));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_1_17_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_1_17_1 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_1_17_1  (
            .in0(N__15102),
            .in1(_gnd_net_),
            .in2(N__14953),
            .in3(N__8911),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_1_17_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_1_17_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(N__14946),
            .in2(_gnd_net_),
            .in3(N__15101),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_18_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(N__9296),
            .in2(N__8915),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_1_18_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_1_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_1_18_1  (
            .in0(_gnd_net_),
            .in1(N__8876),
            .in2(_gnd_net_),
            .in3(N__8699),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_1_18_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_1_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(N__8846),
            .in2(N__8696),
            .in3(N__8678),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_1_18_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_1_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(N__8813),
            .in2(_gnd_net_),
            .in3(N__8666),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_1_18_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_1_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_1_18_4  (
            .in0(_gnd_net_),
            .in1(N__9059),
            .in2(_gnd_net_),
            .in3(N__8654),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_1_18_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_1_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_1_18_5  (
            .in0(_gnd_net_),
            .in1(N__9029),
            .in2(_gnd_net_),
            .in3(N__8642),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_1_18_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_1_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_1_18_6  (
            .in0(_gnd_net_),
            .in1(N__9005),
            .in2(_gnd_net_),
            .in3(N__8630),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_1_18_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_1_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_1_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_1_18_7  (
            .in0(_gnd_net_),
            .in1(N__8981),
            .in2(_gnd_net_),
            .in3(N__8618),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_1_19_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_1_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(N__9148),
            .in2(_gnd_net_),
            .in3(N__8735),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_1_19_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_1_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(N__9193),
            .in2(_gnd_net_),
            .in3(N__8732),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_1_19_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_1_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(N__9172),
            .in2(_gnd_net_),
            .in3(N__8729),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_1_19_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_1_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_1_19_3  (
            .in0(_gnd_net_),
            .in1(N__9262),
            .in2(_gnd_net_),
            .in3(N__8726),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_1_19_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_1_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_1_19_4  (
            .in0(_gnd_net_),
            .in1(N__9217),
            .in2(_gnd_net_),
            .in3(N__8723),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_1_19_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_1_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_1_19_5  (
            .in0(_gnd_net_),
            .in1(N__9379),
            .in2(_gnd_net_),
            .in3(N__8720),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_1_19_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_1_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_1_19_6  (
            .in0(_gnd_net_),
            .in1(N__9283),
            .in2(_gnd_net_),
            .in3(N__8717),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_1_19_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_1_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_1_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_1_19_7  (
            .in0(_gnd_net_),
            .in1(N__9238),
            .in2(_gnd_net_),
            .in3(N__8714),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_1_20_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_1_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_1_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_1_20_0  (
            .in0(_gnd_net_),
            .in1(N__9313),
            .in2(_gnd_net_),
            .in3(N__8711),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ),
            .ltout(),
            .carryin(bfn_1_20_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_1_20_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_1_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_1_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_1_20_1  (
            .in0(_gnd_net_),
            .in1(N__9355),
            .in2(_gnd_net_),
            .in3(N__8789),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_1_20_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_1_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_1_20_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_1_20_2  (
            .in0(_gnd_net_),
            .in1(N__9334),
            .in2(_gnd_net_),
            .in3(N__8786),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_ibuf_gb_io_RNI79U7_LC_1_25_4.C_ON=1'b0;
    defparam reset_ibuf_gb_io_RNI79U7_LC_1_25_4.SEQ_MODE=4'b0000;
    defparam reset_ibuf_gb_io_RNI79U7_LC_1_25_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 reset_ibuf_gb_io_RNI79U7_LC_1_25_4 (
            .in0(N__22339),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(red_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.N_27_i_i_LC_1_29_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.N_27_i_i_LC_1_29_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.N_27_i_i_LC_1_29_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \phase_controller_slave.stoper_tr.N_27_i_i_LC_1_29_1  (
            .in0(_gnd_net_),
            .in1(N__21721),
            .in2(_gnd_net_),
            .in3(N__22340),
            .lcout(N_27_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un7_start_stop_LC_1_30_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un7_start_stop_LC_1_30_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un7_start_stop_LC_1_30_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un7_start_stop_LC_1_30_6  (
            .in0(N__22341),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21725),
            .lcout(un7_start_stop),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_1_30_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_30_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_30_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_30_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_2_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_2_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_2_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11249),
            .lcout(\delay_measurement_inst.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22042),
            .ce(N__10727),
            .sr(N__22254));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_2_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_2_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11216),
            .lcout(\delay_measurement_inst.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22042),
            .ce(N__10727),
            .sr(N__22254));
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_2_14_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_2_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_2_14_1 .LUT_INIT=16'b1000101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_2_LC_2_14_1  (
            .in0(N__13266),
            .in1(N__13327),
            .in2(N__13307),
            .in3(N__13354),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22038),
            .ce(N__13823),
            .sr(N__22260));
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_2_14_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_2_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_2_14_2 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_4_LC_2_14_2  (
            .in0(N__20135),
            .in1(N__13231),
            .in2(N__12857),
            .in3(N__13155),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22038),
            .ce(N__13823),
            .sr(N__22260));
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_2_14_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_2_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_2_14_3 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_5_LC_2_14_3  (
            .in0(N__13156),
            .in1(N__12738),
            .in2(N__13235),
            .in3(N__20136),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22038),
            .ce(N__13823),
            .sr(N__22260));
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_2_14_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_2_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_2_14_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_1_LC_2_14_4  (
            .in0(N__12712),
            .in1(N__13302),
            .in2(N__12700),
            .in3(N__13267),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22038),
            .ce(N__13823),
            .sr(N__22260));
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_2_14_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_2_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_2_14_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_3_LC_2_14_6  (
            .in0(N__13326),
            .in1(N__13306),
            .in2(_gnd_net_),
            .in3(N__13268),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22038),
            .ce(N__13823),
            .sr(N__22260));
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_2_14_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_2_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_2_14_7 .LUT_INIT=16'b0000000011110001;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_6_LC_2_14_7  (
            .in0(N__13157),
            .in1(N__20137),
            .in2(N__13183),
            .in3(N__13232),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22038),
            .ce(N__13823),
            .sr(N__22260));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_2_15_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_2_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__8921),
            .in2(N__8891),
            .in3(N__8907),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_2_15_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_2_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__8882),
            .in2(N__8861),
            .in3(N__8872),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_2_15_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_2_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__8852),
            .in2(N__8831),
            .in3(N__8842),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_2_15_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_2_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__8822),
            .in2(N__8798),
            .in3(N__8809),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_2_15_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_2_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__9068),
            .in2(N__9044),
            .in3(N__9055),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_2_15_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_2_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(N__9035),
            .in2(N__9014),
            .in3(N__9025),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_2_15_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_2_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__9659),
            .in2(N__8990),
            .in3(N__9001),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_2_15_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_2_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(N__9536),
            .in2(N__8966),
            .in3(N__8977),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_2_16_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_2_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__9566),
            .in2(N__8957),
            .in3(N__9149),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_2_16_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_2_16_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_2_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(N__9542),
            .in2(N__8948),
            .in3(N__9194),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_2_16_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_2_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__9653),
            .in2(N__8939),
            .in3(N__9173),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_2_16_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_2_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(N__9560),
            .in2(N__8930),
            .in3(N__9263),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_2_16_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_2_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_2_16_4  (
            .in0(_gnd_net_),
            .in1(N__9551),
            .in2(N__9134),
            .in3(N__9218),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_2_16_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_2_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_2_16_5  (
            .in0(_gnd_net_),
            .in1(N__9614),
            .in2(N__9125),
            .in3(N__9380),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_2_16_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_2_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_2_16_6  (
            .in0(_gnd_net_),
            .in1(N__9626),
            .in2(N__9116),
            .in3(N__9284),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_2_16_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_2_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(N__9635),
            .in2(N__9107),
            .in3(N__9239),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_2_17_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_2_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(N__9620),
            .in2(N__9098),
            .in3(N__9314),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_2_17_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_2_17_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_2_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(N__9641),
            .in2(N__9089),
            .in3(N__9356),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_2_17_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_2_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_2_17_2  (
            .in0(_gnd_net_),
            .in1(N__9647),
            .in2(N__9080),
            .in3(N__9335),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_2_17_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_2_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9071),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_2_17_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_2_17_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_2_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9299),
            .in3(N__14945),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_2_17_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_2_17_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_2_17_5  (
            .in0(N__15171),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15002),
            .lcout(\phase_controller_slave.stoper_tr.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_2_18_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_2_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_2_18_0 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_15_LC_2_18_0  (
            .in0(N__15071),
            .in1(N__19892),
            .in2(N__15263),
            .in3(N__9290),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22026),
            .ce(),
            .sr(N__22284));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_2_18_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_2_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_2_18_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_12_LC_2_18_1  (
            .in0(N__15228),
            .in1(N__15075),
            .in2(N__19904),
            .in3(N__9269),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22026),
            .ce(),
            .sr(N__22284));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_2_18_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_2_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_2_18_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_16_LC_2_18_2  (
            .in0(N__15072),
            .in1(N__19893),
            .in2(N__9248),
            .in3(N__15232),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22026),
            .ce(),
            .sr(N__22284));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_2_18_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_2_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_2_18_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_13_LC_2_18_3  (
            .in0(N__15229),
            .in1(N__15076),
            .in2(N__19905),
            .in3(N__9224),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22026),
            .ce(),
            .sr(N__22284));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_2_18_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_2_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_2_18_4 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_10_LC_2_18_4  (
            .in0(N__15070),
            .in1(N__19891),
            .in2(N__9203),
            .in3(N__15231),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22026),
            .ce(),
            .sr(N__22284));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_2_18_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_2_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_2_18_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_11_LC_2_18_5  (
            .in0(N__15227),
            .in1(N__15074),
            .in2(N__19903),
            .in3(N__9179),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22026),
            .ce(),
            .sr(N__22284));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_2_18_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_2_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_2_18_6 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_9_LC_2_18_6  (
            .in0(N__15073),
            .in1(N__19894),
            .in2(N__9158),
            .in3(N__15233),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22026),
            .ce(),
            .sr(N__22284));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_2_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_2_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_2_18_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_14_LC_2_18_7  (
            .in0(N__15230),
            .in1(N__15077),
            .in2(N__19906),
            .in3(N__9386),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22026),
            .ce(),
            .sr(N__22284));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_2_19_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_2_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_2_19_5 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_18_LC_2_19_5  (
            .in0(N__15235),
            .in1(N__19878),
            .in2(N__9365),
            .in3(N__15079),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22022),
            .ce(),
            .sr(N__22289));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_2_19_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_2_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_2_19_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_19_LC_2_19_6  (
            .in0(N__15078),
            .in1(N__15236),
            .in2(N__19902),
            .in3(N__9341),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22022),
            .ce(),
            .sr(N__22289));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_2_19_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_2_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_2_19_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_17_LC_2_19_7  (
            .in0(N__15234),
            .in1(N__19877),
            .in2(N__15083),
            .in3(N__9320),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22022),
            .ce(),
            .sr(N__22289));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_2_20_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_2_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_2_20_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_4_LC_2_20_0  (
            .in0(N__12354),
            .in1(N__15651),
            .in2(N__12499),
            .in3(N__9398),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22018),
            .ce(),
            .sr(N__22293));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_2_20_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_2_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_2_20_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_6_LC_2_20_1  (
            .in0(N__12484),
            .in1(N__12358),
            .in2(N__15701),
            .in3(N__9494),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22018),
            .ce(),
            .sr(N__22293));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_2_20_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_2_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_2_20_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_2_LC_2_20_2  (
            .in0(N__12353),
            .in1(N__15650),
            .in2(N__12498),
            .in3(N__9422),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22018),
            .ce(),
            .sr(N__22293));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_2_20_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_2_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_2_20_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_1_LC_2_20_3  (
            .in0(N__12482),
            .in1(N__12356),
            .in2(N__15699),
            .in3(N__10136),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22018),
            .ce(),
            .sr(N__22293));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_2_20_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_2_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_2_20_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_5_LC_2_20_4  (
            .in0(N__12355),
            .in1(N__15652),
            .in2(N__12500),
            .in3(N__9506),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22018),
            .ce(),
            .sr(N__22293));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_2_20_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_2_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_2_20_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_3_LC_2_20_5  (
            .in0(N__12483),
            .in1(N__12357),
            .in2(N__15700),
            .in3(N__9410),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22018),
            .ce(),
            .sr(N__22293));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_2_20_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_2_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_2_20_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_7_LC_2_20_7  (
            .in0(N__12485),
            .in1(N__12359),
            .in2(N__15702),
            .in3(N__9482),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22018),
            .ce(),
            .sr(N__22293));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_2_21_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_2_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_2_21_0 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_10_LC_2_21_0  (
            .in0(N__12479),
            .in1(N__15729),
            .in2(N__9446),
            .in3(N__12351),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22013),
            .ce(),
            .sr(N__22297));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_2_21_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_2_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_2_21_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_9_LC_2_21_3  (
            .in0(N__12350),
            .in1(N__12481),
            .in2(N__15737),
            .in3(N__9458),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22013),
            .ce(),
            .sr(N__22297));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_2_21_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_2_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_2_21_4 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_8_LC_2_21_4  (
            .in0(N__12480),
            .in1(N__15730),
            .in2(N__9470),
            .in3(N__12352),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22013),
            .ce(),
            .sr(N__22297));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_2_22_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_2_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_2_22_0  (
            .in0(_gnd_net_),
            .in1(N__10157),
            .in2(N__9929),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_22_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_2_22_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_2_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_2_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_2_22_1  (
            .in0(_gnd_net_),
            .in1(N__9731),
            .in2(_gnd_net_),
            .in3(N__9413),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_2_22_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_2_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_2_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_2_22_2  (
            .in0(_gnd_net_),
            .in1(N__9707),
            .in2(N__10130),
            .in3(N__9401),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_2_22_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_2_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_2_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_2_22_3  (
            .in0(_gnd_net_),
            .in1(N__9683),
            .in2(_gnd_net_),
            .in3(N__9389),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_2_22_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_2_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_2_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_2_22_4  (
            .in0(_gnd_net_),
            .in1(N__9920),
            .in2(_gnd_net_),
            .in3(N__9497),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_2_22_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_2_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_2_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_2_22_5  (
            .in0(_gnd_net_),
            .in1(N__9896),
            .in2(_gnd_net_),
            .in3(N__9485),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_2_22_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_2_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_2_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_2_22_6  (
            .in0(_gnd_net_),
            .in1(N__9869),
            .in2(_gnd_net_),
            .in3(N__9473),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_2_22_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_2_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_2_22_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_2_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9845),
            .in3(N__9461),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_2_23_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_2_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_2_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_2_23_0  (
            .in0(_gnd_net_),
            .in1(N__9821),
            .in2(_gnd_net_),
            .in3(N__9449),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ),
            .ltout(),
            .carryin(bfn_2_23_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_2_23_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_2_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_2_23_1  (
            .in0(_gnd_net_),
            .in1(N__9797),
            .in2(_gnd_net_),
            .in3(N__9434),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_2_23_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_2_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_2_23_2  (
            .in0(_gnd_net_),
            .in1(N__10114),
            .in2(_gnd_net_),
            .in3(N__9431),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_2_23_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_2_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_2_23_3  (
            .in0(_gnd_net_),
            .in1(N__10012),
            .in2(_gnd_net_),
            .in3(N__9428),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_2_23_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_2_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_2_23_4  (
            .in0(_gnd_net_),
            .in1(N__10075),
            .in2(_gnd_net_),
            .in3(N__9425),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_2_23_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_2_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_2_23_5  (
            .in0(_gnd_net_),
            .in1(N__10033),
            .in2(_gnd_net_),
            .in3(N__9524),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_2_23_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_2_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_2_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_2_23_6  (
            .in0(_gnd_net_),
            .in1(N__10054),
            .in2(_gnd_net_),
            .in3(N__9521),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_2_23_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_2_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_2_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_2_23_7  (
            .in0(_gnd_net_),
            .in1(N__10094),
            .in2(_gnd_net_),
            .in3(N__9518),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_2_24_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_2_24_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_2_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_2_24_0  (
            .in0(_gnd_net_),
            .in1(N__10210),
            .in2(_gnd_net_),
            .in3(N__9515),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ),
            .ltout(),
            .carryin(bfn_2_24_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_2_24_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_2_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_2_24_1  (
            .in0(_gnd_net_),
            .in1(N__10189),
            .in2(_gnd_net_),
            .in3(N__9512),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_2_24_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_2_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_2_24_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_2_24_2  (
            .in0(_gnd_net_),
            .in1(N__10231),
            .in2(_gnd_net_),
            .in3(N__9509),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_3_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_3_12_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_3_12_1 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_8_LC_3_12_1  (
            .in0(N__11034),
            .in1(N__10169),
            .in2(N__12776),
            .in3(N__10310),
            .lcout(measured_delay_tr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22043),
            .ce(),
            .sr(N__22242));
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_3_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_3_12_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_3_12_5 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_7_LC_3_12_5  (
            .in0(N__11033),
            .in1(N__10168),
            .in2(N__12817),
            .in3(N__10334),
            .lcout(measured_delay_tr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22043),
            .ce(),
            .sr(N__22242));
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_3_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_3_13_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_3_13_0 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_5_LC_3_13_0  (
            .in0(N__11067),
            .in1(N__11029),
            .in2(N__10998),
            .in3(N__10385),
            .lcout(measured_delay_tr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22039),
            .ce(N__11274),
            .sr(N__22248));
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_3_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_3_13_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_3_13_1 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_2_LC_3_13_1  (
            .in0(N__9591),
            .in1(N__10986),
            .in2(N__11036),
            .in3(N__11066),
            .lcout(measured_delay_tr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22039),
            .ce(N__11274),
            .sr(N__22248));
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_3_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_3_13_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_3_13_2 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_16_LC_3_13_2  (
            .in0(N__11364),
            .in1(_gnd_net_),
            .in2(N__10481),
            .in3(N__20940),
            .lcout(measured_delay_tr_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22039),
            .ce(N__11274),
            .sr(N__22248));
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_3_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_3_13_3 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_3_13_3 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_1_LC_3_13_3  (
            .in0(N__11031),
            .in1(N__10991),
            .in2(N__9608),
            .in3(N__11069),
            .lcout(measured_delay_tr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22039),
            .ce(N__11274),
            .sr(N__22248));
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_3_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_3_13_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_3_13_4 .LUT_INIT=16'b0011000000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_15_LC_3_13_4  (
            .in0(N__11363),
            .in1(N__10282),
            .in2(N__10528),
            .in3(N__20942),
            .lcout(measured_delay_tr_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22039),
            .ce(N__11274),
            .sr(N__22248));
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_3_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_3_13_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_3_13_5 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_14_LC_3_13_5  (
            .in0(N__20941),
            .in1(N__10563),
            .in2(N__10283),
            .in3(N__11362),
            .lcout(measured_delay_tr_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22039),
            .ce(N__11274),
            .sr(N__22248));
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_3_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_3_13_6 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_3_13_6 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_3_LC_3_13_6  (
            .in0(N__11070),
            .in1(N__11032),
            .in2(N__10999),
            .in3(N__10412),
            .lcout(measured_delay_tr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22039),
            .ce(N__11274),
            .sr(N__22248));
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_3_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_3_13_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_3_13_7 .LUT_INIT=16'b0011000111110101;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_6_LC_3_13_7  (
            .in0(N__11030),
            .in1(N__10990),
            .in2(N__10367),
            .in3(N__11068),
            .lcout(measured_delay_tr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22039),
            .ce(N__11274),
            .sr(N__22248));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_3_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_3_14_0 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_3_14_0  (
            .in0(N__20070),
            .in1(N__19996),
            .in2(_gnd_net_),
            .in3(N__12952),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_3_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_3_14_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_3_14_1  (
            .in0(N__10302),
            .in1(N__10329),
            .in2(_gnd_net_),
            .in3(N__10353),
            .lcout(\delay_measurement_inst.N_212 ),
            .ltout(\delay_measurement_inst.N_212_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIC9OF1_14_LC_3_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIC9OF1_14_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIC9OF1_14_LC_3_14_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIC9OF1_14_LC_3_14_2  (
            .in0(N__10524),
            .in1(N__10561),
            .in2(N__9527),
            .in3(N__10423),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_3_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_3_14_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_3_14_3  (
            .in0(_gnd_net_),
            .in1(N__13325),
            .in2(_gnd_net_),
            .in3(N__13353),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_3_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_3_14_4 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_3_14_4  (
            .in0(N__11361),
            .in1(_gnd_net_),
            .in2(N__10529),
            .in3(N__10256),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6FAF_1_LC_3_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6FAF_1_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6FAF_1_LC_3_14_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6FAF_1_LC_3_14_5  (
            .in0(N__9592),
            .in1(N__9604),
            .in2(N__10360),
            .in3(N__11090),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_3_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_3_14_6 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_3_14_6  (
            .in0(N__10404),
            .in1(N__9593),
            .in2(N__11098),
            .in3(N__10430),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_3_14_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_3_14_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_3_14_7  (
            .in0(N__10255),
            .in1(N__9575),
            .in2(N__9569),
            .in3(N__11360),
            .lcout(\delay_measurement_inst.N_168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_3_15_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_3_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_3_15_0 .LUT_INIT=16'b1111010011110101;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_9_LC_3_15_0  (
            .in0(N__12906),
            .in1(N__20020),
            .in2(N__12586),
            .in3(N__12544),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22035),
            .ce(N__13822),
            .sr(N__22261));
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_3_15_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_3_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_3_15_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_12_LC_3_15_2  (
            .in0(N__12904),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13019),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22035),
            .ce(N__13822),
            .sr(N__22261));
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_3_15_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_3_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_3_15_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_13_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__12905),
            .in2(_gnd_net_),
            .in3(N__12994),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22035),
            .ce(N__13822),
            .sr(N__22261));
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_3_15_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_3_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_3_15_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_10_LC_3_15_4  (
            .in0(N__12881),
            .in1(_gnd_net_),
            .in2(N__12910),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22035),
            .ce(N__13822),
            .sr(N__22261));
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_3_15_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_3_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_3_15_5 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_8_LC_3_15_5  (
            .in0(N__13154),
            .in1(_gnd_net_),
            .in2(N__20131),
            .in3(N__12777),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22035),
            .ce(N__13822),
            .sr(N__22261));
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_3_15_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_3_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_3_15_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_7_LC_3_15_6  (
            .in0(N__12818),
            .in1(N__20109),
            .in2(_gnd_net_),
            .in3(N__13153),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22035),
            .ce(N__13822),
            .sr(N__22261));
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_3_15_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_3_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_3_15_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_11_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(N__12903),
            .in2(_gnd_net_),
            .in3(N__12611),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22035),
            .ce(N__13822),
            .sr(N__22261));
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_3_16_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_3_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_3_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_19_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13783),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22031),
            .ce(N__13812),
            .sr(N__22270));
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_3_16_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_3_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_3_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_18_LC_3_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13690),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22031),
            .ce(N__13812),
            .sr(N__22270));
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_3_16_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_3_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_3_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_16_LC_3_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13648),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22031),
            .ce(N__13812),
            .sr(N__22270));
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_3_16_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_3_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_3_16_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_15_LC_3_16_5  (
            .in0(N__20018),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20130),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22031),
            .ce(N__13812),
            .sr(N__22270));
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_3_16_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_3_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_3_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_17_LC_3_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13732),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22031),
            .ce(N__13812),
            .sr(N__22270));
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_3_16_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_3_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_3_16_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_14_LC_3_16_7  (
            .in0(N__20019),
            .in1(N__20129),
            .in2(_gnd_net_),
            .in3(N__12961),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22031),
            .ce(N__13812),
            .sr(N__22270));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIE5AP1_23_LC_3_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIE5AP1_23_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIE5AP1_23_LC_3_17_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIE5AP1_23_LC_3_17_4  (
            .in0(N__10640),
            .in1(N__10649),
            .in2(N__10781),
            .in3(N__10658),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_3_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_3_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_3_17_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_3_17_6  (
            .in0(_gnd_net_),
            .in1(N__10667),
            .in2(_gnd_net_),
            .in3(N__10676),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_3_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_3_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_3_17_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_3_17_7  (
            .in0(N__10685),
            .in1(N__9746),
            .in2(N__9755),
            .in3(N__9752),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_3_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_3_18_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_3_18_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_3_18_7  (
            .in0(N__10751),
            .in1(N__10760),
            .in2(N__10742),
            .in3(N__10769),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_3_19_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_3_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(N__10841),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_19_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__10850),
            .in2(N__9740),
            .in3(N__10152),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_19_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__10856),
            .in2(N__9716),
            .in3(N__9727),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_19_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(N__10700),
            .in2(N__9692),
            .in3(N__9703),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_19_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_19_4  (
            .in0(_gnd_net_),
            .in1(N__10826),
            .in2(N__9668),
            .in3(N__9679),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_19_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_19_5  (
            .in0(_gnd_net_),
            .in1(N__10706),
            .in2(N__9905),
            .in3(N__9916),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_19_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__10835),
            .in2(N__9878),
            .in3(N__9895),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_19_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(N__10862),
            .in2(N__9854),
            .in3(N__9865),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_20_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_20_0  (
            .in0(_gnd_net_),
            .in1(N__10913),
            .in2(N__9830),
            .in3(N__9841),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_3_20_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_20_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_20_1  (
            .in0(_gnd_net_),
            .in1(N__10892),
            .in2(N__9806),
            .in3(N__9817),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_20_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_20_2  (
            .in0(_gnd_net_),
            .in1(N__10808),
            .in2(N__9782),
            .in3(N__9793),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_20_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_20_3  (
            .in0(_gnd_net_),
            .in1(N__10790),
            .in2(N__9773),
            .in3(N__10115),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_20_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_20_4  (
            .in0(_gnd_net_),
            .in1(N__10817),
            .in2(N__9764),
            .in3(N__10013),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_20_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_20_5  (
            .in0(_gnd_net_),
            .in1(N__10799),
            .in2(N__9998),
            .in3(N__10076),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_20_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_20_6  (
            .in0(_gnd_net_),
            .in1(N__10898),
            .in2(N__9989),
            .in3(N__10034),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_20_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_20_7  (
            .in0(_gnd_net_),
            .in1(N__10904),
            .in2(N__9980),
            .in3(N__10055),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_21_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_21_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_21_0  (
            .in0(N__10093),
            .in1(N__10874),
            .in2(N__9971),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_3_21_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_21_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_21_1  (
            .in0(_gnd_net_),
            .in1(N__10868),
            .in2(N__9962),
            .in3(N__10211),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_21_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_21_2  (
            .in0(_gnd_net_),
            .in1(N__10880),
            .in2(N__9953),
            .in3(N__10190),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_21_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_21_3  (
            .in0(_gnd_net_),
            .in1(N__10886),
            .in2(N__9944),
            .in3(N__10232),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_21_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9935),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_21_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_21_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9932),
            .in3(N__18101),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_3_21_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_3_21_6 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_3_21_6  (
            .in0(N__18051),
            .in1(_gnd_net_),
            .in2(N__18109),
            .in3(N__10156),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_3_21_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_3_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_3_21_7  (
            .in0(_gnd_net_),
            .in1(N__18102),
            .in2(_gnd_net_),
            .in3(N__18050),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_3_22_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_3_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_3_22_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_11_LC_3_22_0  (
            .in0(N__12467),
            .in1(N__12347),
            .in2(N__15734),
            .in3(N__10121),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22000),
            .ce(),
            .sr(N__22298));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_3_22_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_3_22_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_3_22_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_16_LC_3_22_1  (
            .in0(N__12346),
            .in1(N__15716),
            .in2(N__12497),
            .in3(N__10100),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22000),
            .ce(),
            .sr(N__22298));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_3_22_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_3_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_3_22_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_13_LC_3_22_2  (
            .in0(N__12468),
            .in1(N__12348),
            .in2(N__15735),
            .in3(N__10082),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22000),
            .ce(),
            .sr(N__22298));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_3_22_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_3_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_3_22_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_15_LC_3_22_4  (
            .in0(N__12469),
            .in1(N__12349),
            .in2(N__15736),
            .in3(N__10061),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22000),
            .ce(),
            .sr(N__22298));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_3_22_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_3_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_3_22_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_14_LC_3_22_5  (
            .in0(N__12345),
            .in1(N__15715),
            .in2(N__12496),
            .in3(N__10040),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22000),
            .ce(),
            .sr(N__22298));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_3_22_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_3_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_3_22_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_12_LC_3_22_7  (
            .in0(N__12344),
            .in1(N__15714),
            .in2(N__12495),
            .in3(N__10019),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22000),
            .ce(),
            .sr(N__22298));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_3_23_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_3_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_3_23_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_19_LC_3_23_2  (
            .in0(N__12293),
            .in1(N__15703),
            .in2(N__12464),
            .in3(N__10238),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21995),
            .ce(),
            .sr(N__22301));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_3_23_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_3_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_3_23_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_17_LC_3_23_3  (
            .in0(N__12414),
            .in1(N__12294),
            .in2(N__15731),
            .in3(N__10217),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21995),
            .ce(),
            .sr(N__22301));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_3_23_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_3_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_3_23_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_18_LC_3_23_5  (
            .in0(N__12415),
            .in1(N__12295),
            .in2(N__15732),
            .in3(N__10196),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21995),
            .ce(),
            .sr(N__22301));
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_3_24_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_3_24_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_3_24_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_0_LC_3_24_6  (
            .in0(N__12416),
            .in1(N__12296),
            .in2(N__15733),
            .in3(N__18060),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21992),
            .ce(N__21289),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_3_24_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_3_24_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_3_24_7 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_1_LC_3_24_7  (
            .in0(N__18061),
            .in1(N__15710),
            .in2(N__12341),
            .in3(N__12417),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21992),
            .ce(N__21289),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_4_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_4_12_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_4_12_1 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_12_LC_4_12_1  (
            .in0(N__11321),
            .in1(N__20939),
            .in2(_gnd_net_),
            .in3(N__10589),
            .lcout(measured_delay_tr_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22040),
            .ce(N__11281),
            .sr(N__22241));
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_4_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_4_12_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_4_12_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_10_LC_4_12_2  (
            .in0(N__20937),
            .in1(N__11322),
            .in2(_gnd_net_),
            .in3(N__10628),
            .lcout(measured_delay_tr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22040),
            .ce(N__11281),
            .sr(N__22241));
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_4_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_4_12_3 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_11_LC_4_12_3  (
            .in0(N__11320),
            .in1(N__20938),
            .in2(_gnd_net_),
            .in3(N__10610),
            .lcout(measured_delay_tr_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22040),
            .ce(N__11281),
            .sr(N__22241));
    defparam \delay_measurement_inst.tr_state_RNI5KUTL_0_LC_4_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_RNI5KUTL_0_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.tr_state_RNI5KUTL_0_LC_4_13_0 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \delay_measurement_inst.tr_state_RNI5KUTL_0_LC_4_13_0  (
            .in0(N__11060),
            .in1(N__10262),
            .in2(N__20873),
            .in3(N__10175),
            .lcout(\delay_measurement_inst.N_81_i ),
            .ltout(\delay_measurement_inst.N_81_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_state_RNICTS5M_0_LC_4_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_RNICTS5M_0_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.tr_state_RNICTS5M_0_LC_4_13_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \delay_measurement_inst.tr_state_RNICTS5M_0_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10160),
            .in3(N__22335),
            .lcout(\delay_measurement_inst.N_81_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA9RL2_15_LC_4_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA9RL2_15_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA9RL2_15_LC_4_13_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA9RL2_15_LC_4_13_2  (
            .in0(N__20935),
            .in1(N__10519),
            .in2(_gnd_net_),
            .in3(N__10455),
            .lcout(\delay_measurement_inst.N_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_4_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_4_13_4 .LUT_INIT=16'b0000000011110001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_4_13_4  (
            .in0(N__10562),
            .in1(N__10520),
            .in2(N__10456),
            .in3(N__11377),
            .lcout(\delay_measurement_inst.N_197_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_4_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_4_13_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_4_13_5  (
            .in0(N__13677),
            .in1(N__13719),
            .in2(N__13784),
            .in3(N__13640),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_4_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_4_13_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_4_13_6  (
            .in0(N__13008),
            .in1(N__12603),
            .in2(N__12987),
            .in3(N__12873),
            .lcout(\phase_controller_inst1.stoper_tr.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_4_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_4_13_7 .LUT_INIT=16'b1101110111011100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_4_13_7  (
            .in0(N__11378),
            .in1(N__20936),
            .in2(N__10457),
            .in3(N__10244),
            .lcout(\delay_measurement_inst.N_165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBIVI2_3_LC_4_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBIVI2_3_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBIVI2_3_LC_4_14_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBIVI2_3_LC_4_14_0  (
            .in0(N__10564),
            .in1(N__10448),
            .in2(N__10411),
            .in3(N__10424),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAFV93_7_LC_4_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAFV93_7_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAFV93_7_LC_4_14_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAFV93_7_LC_4_14_1  (
            .in0(N__10271),
            .in1(N__10303),
            .in2(N__10265),
            .in3(N__10330),
            .lcout(\delay_measurement_inst.un1_tr_state_1_i_0_a2_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_4_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_4_14_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_4_14_2  (
            .in0(N__10588),
            .in1(N__10609),
            .in2(N__11303),
            .in3(N__10624),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_4_14_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_4_14_3 .LUT_INIT=16'b0001000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_4_14_3  (
            .in0(N__11094),
            .in1(N__10518),
            .in2(N__10247),
            .in3(N__10565),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_4_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_4_14_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_4_14_5  (
            .in0(N__10477),
            .in1(N__11427),
            .in2(N__11405),
            .in3(N__11449),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_4_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_4_14_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_4_14_6  (
            .in0(N__11448),
            .in1(N__11400),
            .in2(N__11429),
            .in3(N__10476),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_4_14_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_4_14_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(N__10381),
            .in2(_gnd_net_),
            .in3(N__10960),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_4_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_4_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_4_15_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__11242),
            .in2(N__11188),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_4_15_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__22032),
            .ce(N__10726),
            .sr(N__22255));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_4_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_4_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_4_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__11209),
            .in2(N__11164),
            .in3(N__10388),
            .lcout(\delay_measurement_inst.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__22032),
            .ce(N__10726),
            .sr(N__22255));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_4_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_4_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_4_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(N__11139),
            .in2(N__11189),
            .in3(N__10370),
            .lcout(\delay_measurement_inst.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__22032),
            .ce(N__10726),
            .sr(N__22255));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_4_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_4_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_4_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(N__11625),
            .in2(N__11165),
            .in3(N__10337),
            .lcout(\delay_measurement_inst.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__22032),
            .ce(N__10726),
            .sr(N__22255));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_4_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_4_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_4_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__11140),
            .in2(N__11608),
            .in3(N__10313),
            .lcout(\delay_measurement_inst.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__22032),
            .ce(N__10726),
            .sr(N__22255));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_4_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_4_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_4_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__11626),
            .in2(N__11584),
            .in3(N__10286),
            .lcout(\delay_measurement_inst.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__22032),
            .ce(N__10726),
            .sr(N__22255));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_4_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_4_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_4_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(N__11559),
            .in2(N__11609),
            .in3(N__10631),
            .lcout(\delay_measurement_inst.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__22032),
            .ce(N__10726),
            .sr(N__22255));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_4_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_4_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_4_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(N__11540),
            .in2(N__11585),
            .in3(N__10613),
            .lcout(\delay_measurement_inst.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__22032),
            .ce(N__10726),
            .sr(N__22255));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_4_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_4_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_4_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__11561),
            .in2(N__11515),
            .in3(N__10592),
            .lcout(\delay_measurement_inst.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_4_16_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__22027),
            .ce(N__10725),
            .sr(N__22262));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_4_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_4_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_4_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__11539),
            .in2(N__11491),
            .in3(N__10571),
            .lcout(\delay_measurement_inst.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__22027),
            .ce(N__10725),
            .sr(N__22262));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_4_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_4_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_4_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(N__11466),
            .in2(N__11516),
            .in3(N__10568),
            .lcout(\delay_measurement_inst.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__22027),
            .ce(N__10725),
            .sr(N__22262));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_4_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_4_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_4_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(N__11820),
            .in2(N__11492),
            .in3(N__10532),
            .lcout(\delay_measurement_inst.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__22027),
            .ce(N__10725),
            .sr(N__22262));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_4_16_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_4_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_4_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(N__11467),
            .in2(N__11803),
            .in3(N__10484),
            .lcout(\delay_measurement_inst.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__22027),
            .ce(N__10725),
            .sr(N__22262));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_4_16_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_4_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_4_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(N__11821),
            .in2(N__11779),
            .in3(N__10460),
            .lcout(\delay_measurement_inst.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__22027),
            .ce(N__10725),
            .sr(N__22262));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_4_16_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_4_16_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_4_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(N__11756),
            .in2(N__11804),
            .in3(N__10694),
            .lcout(\delay_measurement_inst.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__22027),
            .ce(N__10725),
            .sr(N__22262));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_4_16_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_4_16_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_4_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_4_16_7  (
            .in0(_gnd_net_),
            .in1(N__11732),
            .in2(N__11780),
            .in3(N__10691),
            .lcout(\delay_measurement_inst.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__22027),
            .ce(N__10725),
            .sr(N__22262));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_4_17_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_4_17_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_4_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_4_17_0  (
            .in0(_gnd_net_),
            .in1(N__11755),
            .in2(N__11707),
            .in3(N__10688),
            .lcout(\delay_measurement_inst.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_4_17_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__22023),
            .ce(N__10724),
            .sr(N__22271));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_4_17_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_4_17_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_4_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_4_17_1  (
            .in0(_gnd_net_),
            .in1(N__11731),
            .in2(N__11683),
            .in3(N__10679),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__22023),
            .ce(N__10724),
            .sr(N__22271));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_4_17_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_4_17_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_4_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_4_17_2  (
            .in0(_gnd_net_),
            .in1(N__11658),
            .in2(N__11708),
            .in3(N__10670),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__22023),
            .ce(N__10724),
            .sr(N__22271));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_4_17_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_4_17_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_4_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_4_17_3  (
            .in0(_gnd_net_),
            .in1(N__11640),
            .in2(N__11684),
            .in3(N__10661),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__22023),
            .ce(N__10724),
            .sr(N__22271));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_4_17_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_4_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_4_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_4_17_4  (
            .in0(_gnd_net_),
            .in1(N__11659),
            .in2(N__12133),
            .in3(N__10652),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__22023),
            .ce(N__10724),
            .sr(N__22271));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_4_17_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_4_17_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_4_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_4_17_5  (
            .in0(_gnd_net_),
            .in1(N__11641),
            .in2(N__12109),
            .in3(N__10643),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__22023),
            .ce(N__10724),
            .sr(N__22271));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_4_17_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_4_17_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_4_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_4_17_6  (
            .in0(_gnd_net_),
            .in1(N__12086),
            .in2(N__12134),
            .in3(N__10634),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__22023),
            .ce(N__10724),
            .sr(N__22271));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_4_17_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_4_17_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_4_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_4_17_7  (
            .in0(_gnd_net_),
            .in1(N__12062),
            .in2(N__12110),
            .in3(N__10772),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__22023),
            .ce(N__10724),
            .sr(N__22271));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_4_18_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_4_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_4_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(N__12085),
            .in2(N__12037),
            .in3(N__10763),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_4_18_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__22019),
            .ce(N__10723),
            .sr(N__22275));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_4_18_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_4_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_4_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_4_18_1  (
            .in0(_gnd_net_),
            .in1(N__12061),
            .in2(N__12013),
            .in3(N__10754),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__22019),
            .ce(N__10723),
            .sr(N__22275));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_4_18_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_4_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_4_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_4_18_2  (
            .in0(_gnd_net_),
            .in1(N__11989),
            .in2(N__12038),
            .in3(N__10745),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__22019),
            .ce(N__10723),
            .sr(N__22275));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_4_18_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_4_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_4_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_4_18_3  (
            .in0(_gnd_net_),
            .in1(N__11851),
            .in2(N__12014),
            .in3(N__10733),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__22019),
            .ce(N__10723),
            .sr(N__22275));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_4_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_4_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_4_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_4_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10730),
            .lcout(\delay_measurement_inst.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22019),
            .ce(N__10723),
            .sr(N__22275));
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_4_19_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_4_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_4_19_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_5_LC_4_19_0  (
            .in0(N__15353),
            .in1(N__14731),
            .in2(_gnd_net_),
            .in3(N__15455),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22014),
            .ce(N__12245),
            .sr(N__22279));
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_4_19_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_4_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_4_19_1 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_3_LC_4_19_1  (
            .in0(N__15580),
            .in1(N__13591),
            .in2(N__15920),
            .in3(N__14665),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22014),
            .ce(N__12245),
            .sr(N__22279));
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_4_19_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_4_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_4_19_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_7_LC_4_19_2  (
            .in0(N__15354),
            .in1(N__16148),
            .in2(_gnd_net_),
            .in3(N__15456),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22014),
            .ce(N__12245),
            .sr(N__22279));
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_4_19_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_4_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_4_19_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_2_LC_4_19_3  (
            .in0(N__15453),
            .in1(N__13589),
            .in2(N__16106),
            .in3(N__15356),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22014),
            .ce(N__12245),
            .sr(N__22279));
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_4_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_4_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_4_19_4 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_1_LC_4_19_4  (
            .in0(N__13590),
            .in1(N__15916),
            .in2(N__14222),
            .in3(N__15579),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22014),
            .ce(N__12245),
            .sr(N__22279));
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_4_19_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_4_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_4_19_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_0_LC_4_19_5  (
            .in0(N__15452),
            .in1(N__13588),
            .in2(N__14129),
            .in3(N__15355),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22014),
            .ce(N__12245),
            .sr(N__22279));
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_4_19_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_4_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_4_19_6 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_4_19_6  (
            .in0(N__14569),
            .in1(N__15915),
            .in2(_gnd_net_),
            .in3(N__15578),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22014),
            .ce(N__12245),
            .sr(N__22279));
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_4_19_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_4_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_4_19_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_4_LC_4_19_7  (
            .in0(N__15454),
            .in1(N__15352),
            .in2(_gnd_net_),
            .in3(N__14264),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22014),
            .ce(N__12245),
            .sr(N__22279));
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_4_20_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_4_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_4_20_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_12_LC_4_20_0  (
            .in0(N__15331),
            .in1(N__16013),
            .in2(_gnd_net_),
            .in3(N__15436),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22008),
            .ce(N__12241),
            .sr(N__22285));
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_4_20_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_4_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_4_20_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_10_LC_4_20_2  (
            .in0(N__15329),
            .in1(N__15965),
            .in2(_gnd_net_),
            .in3(N__15434),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22008),
            .ce(N__12241),
            .sr(N__22285));
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_4_20_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_4_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_4_20_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_13_LC_4_20_3  (
            .in0(N__15437),
            .in1(N__15332),
            .in2(_gnd_net_),
            .in3(N__14510),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22008),
            .ce(N__12241),
            .sr(N__22285));
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_4_20_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_4_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_4_20_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_11_LC_4_20_5  (
            .in0(N__15435),
            .in1(N__15330),
            .in2(_gnd_net_),
            .in3(N__15785),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22008),
            .ce(N__12241),
            .sr(N__22285));
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_4_20_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_4_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_4_20_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_8_LC_4_20_6  (
            .in0(N__16059),
            .in1(_gnd_net_),
            .in2(N__15357),
            .in3(N__15439),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22008),
            .ce(N__12241),
            .sr(N__22285));
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_4_20_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_4_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_4_20_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_15_LC_4_20_7  (
            .in0(N__15438),
            .in1(N__15333),
            .in2(_gnd_net_),
            .in3(N__14398),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22008),
            .ce(N__12241),
            .sr(N__22285));
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_4_21_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_4_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_4_21_3 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_14_LC_4_21_3  (
            .in0(N__15895),
            .in1(N__14830),
            .in2(_gnd_net_),
            .in3(N__15553),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22001),
            .ce(N__12240),
            .sr(N__22290));
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_4_21_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_4_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_4_21_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_9_LC_4_21_4  (
            .in0(N__15554),
            .in1(N__15896),
            .in2(_gnd_net_),
            .in3(N__16195),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22001),
            .ce(N__12240),
            .sr(N__22290));
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_4_22_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_4_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_4_22_2 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_19_LC_4_22_2  (
            .in0(N__14457),
            .in1(N__15892),
            .in2(_gnd_net_),
            .in3(N__15533),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21996),
            .ce(N__12239),
            .sr(N__22294));
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_4_22_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_4_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_4_22_5 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_18_LC_4_22_5  (
            .in0(N__15532),
            .in1(_gnd_net_),
            .in2(N__15906),
            .in3(N__14338),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21996),
            .ce(N__12239),
            .sr(N__22294));
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_4_22_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_4_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_4_22_6 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_16_LC_4_22_6  (
            .in0(N__14875),
            .in1(N__15885),
            .in2(_gnd_net_),
            .in3(N__15530),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21996),
            .ce(N__12239),
            .sr(N__22294));
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_4_22_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_4_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_4_22_7 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_17_LC_4_22_7  (
            .in0(N__15531),
            .in1(_gnd_net_),
            .in2(N__15905),
            .in3(N__14616),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21996),
            .ce(N__12239),
            .sr(N__22294));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_4_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_4_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_4_23_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_4_23_0  (
            .in0(N__14876),
            .in1(N__14507),
            .in2(N__14570),
            .in3(N__15959),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_4_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_4_23_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_4_23_2  (
            .in0(N__14339),
            .in1(N__14722),
            .in2(N__14459),
            .in3(N__14262),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_4_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_4_23_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_4_23_4  (
            .in0(N__16139),
            .in1(N__16006),
            .in2(N__16061),
            .in3(N__15778),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_15_LC_4_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_15_LC_4_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_15_LC_4_23_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_15_LC_4_23_5  (
            .in0(N__12644),
            .in1(N__18735),
            .in2(N__10949),
            .in3(N__18691),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_4_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_4_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_4_23_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_LC_4_23_6  (
            .in0(N__10946),
            .in1(N__10940),
            .in2(N__10934),
            .in3(N__12668),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlt31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_4_23_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_4_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_4_23_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_4_23_7  (
            .in0(_gnd_net_),
            .in1(N__12396),
            .in2(_gnd_net_),
            .in3(N__12279),
            .lcout(\phase_controller_slave.stoper_hc.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_12_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_12_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_12_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_5_12_2 (
            .in0(N__10931),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22037),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_12_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_12_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_5_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10919),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22037),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_5_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_5_12_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__21485),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_5_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_5_13_0 .LUT_INIT=16'b0000011100000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_5_13_0  (
            .in0(N__12957),
            .in1(N__12566),
            .in2(N__20027),
            .in3(N__12535),
            .lcout(\phase_controller_inst1.stoper_tr.N_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_5_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_5_13_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_5_13_1  (
            .in0(N__13676),
            .in1(N__13718),
            .in2(N__13769),
            .in3(N__13644),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_4_3_LC_5_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_4_3_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_4_3_LC_5_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_4_3_LC_5_13_2  (
            .in0(N__12956),
            .in1(N__12739),
            .in2(N__20026),
            .in3(N__12843),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_4Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_6_3_LC_5_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_6_3_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_6_3_LC_5_13_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_6_3_LC_5_13_3  (
            .in0(N__12822),
            .in1(N__11111),
            .in2(N__11123),
            .in3(N__11120),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_6Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_5_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_5_13_4 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__12567),
            .in2(N__11114),
            .in3(N__12537),
            .lcout(\phase_controller_inst1.stoper_tr.N_109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0_6_LC_5_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0_6_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0_6_LC_5_13_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0_6_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(N__12778),
            .in2(_gnd_net_),
            .in3(N__13179),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_5_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_5_13_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_5_13_6  (
            .in0(N__20014),
            .in1(N__12823),
            .in2(N__11105),
            .in3(N__12536),
            .lcout(\phase_controller_inst1.stoper_tr.N_92 ),
            .ltout(\phase_controller_inst1.stoper_tr.N_92_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_5_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_5_13_7 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_5_13_7  (
            .in0(N__20071),
            .in1(_gnd_net_),
            .in2(N__11102),
            .in3(N__13118),
            .lcout(\phase_controller_inst1.stoper_tr.N_110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_5_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_5_14_1 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_9_LC_5_14_1  (
            .in0(N__20947),
            .in1(N__11324),
            .in2(N__11099),
            .in3(N__11071),
            .lcout(measured_delay_tr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22033),
            .ce(N__11282),
            .sr(N__22243));
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_5_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_5_14_2 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_4_LC_5_14_2  (
            .in0(N__11072),
            .in1(N__11035),
            .in2(N__11000),
            .in3(N__10961),
            .lcout(measured_delay_tr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22033),
            .ce(N__11282),
            .sr(N__22243));
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_5_14_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_5_14_3 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_18_LC_5_14_3  (
            .in0(N__20945),
            .in1(N__11450),
            .in2(_gnd_net_),
            .in3(N__11380),
            .lcout(measured_delay_tr_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22033),
            .ce(N__11282),
            .sr(N__22243));
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_5_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_5_14_4 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_19_LC_5_14_4  (
            .in0(N__11381),
            .in1(N__20946),
            .in2(_gnd_net_),
            .in3(N__11428),
            .lcout(measured_delay_tr_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22033),
            .ce(N__11282),
            .sr(N__22243));
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_5_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_5_14_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_5_14_5 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_17_LC_5_14_5  (
            .in0(N__20944),
            .in1(N__11404),
            .in2(_gnd_net_),
            .in3(N__11379),
            .lcout(measured_delay_tr_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22033),
            .ce(N__11282),
            .sr(N__22243));
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_5_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_5_14_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_5_14_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_13_LC_5_14_6  (
            .in0(N__11323),
            .in1(N__20943),
            .in2(_gnd_net_),
            .in3(N__11302),
            .lcout(measured_delay_tr_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22033),
            .ce(N__11282),
            .sr(N__22243));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_5_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_5_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_5_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_5_15_0  (
            .in0(N__11972),
            .in1(N__11235),
            .in2(_gnd_net_),
            .in3(N__11219),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__22028),
            .ce(N__11837),
            .sr(N__22249));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_5_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_5_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_5_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_5_15_1  (
            .in0(N__11968),
            .in1(N__11208),
            .in2(_gnd_net_),
            .in3(N__11192),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__22028),
            .ce(N__11837),
            .sr(N__22249));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_5_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_5_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_5_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_5_15_2  (
            .in0(N__11973),
            .in1(N__11187),
            .in2(_gnd_net_),
            .in3(N__11168),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__22028),
            .ce(N__11837),
            .sr(N__22249));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_5_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_5_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_5_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_5_15_3  (
            .in0(N__11969),
            .in1(N__11163),
            .in2(_gnd_net_),
            .in3(N__11144),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__22028),
            .ce(N__11837),
            .sr(N__22249));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_5_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_5_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_5_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_5_15_4  (
            .in0(N__11974),
            .in1(N__11141),
            .in2(_gnd_net_),
            .in3(N__11126),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__22028),
            .ce(N__11837),
            .sr(N__22249));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_5_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_5_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_5_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_5_15_5  (
            .in0(N__11970),
            .in1(N__11627),
            .in2(_gnd_net_),
            .in3(N__11612),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__22028),
            .ce(N__11837),
            .sr(N__22249));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_5_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_5_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_5_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_5_15_6  (
            .in0(N__11975),
            .in1(N__11607),
            .in2(_gnd_net_),
            .in3(N__11588),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__22028),
            .ce(N__11837),
            .sr(N__22249));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_5_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_5_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_5_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_5_15_7  (
            .in0(N__11971),
            .in1(N__11583),
            .in2(_gnd_net_),
            .in3(N__11564),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__22028),
            .ce(N__11837),
            .sr(N__22249));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_5_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_5_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_5_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_5_16_0  (
            .in0(N__11949),
            .in1(N__11560),
            .in2(_gnd_net_),
            .in3(N__11543),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_5_16_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__22024),
            .ce(N__11838),
            .sr(N__22256));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_5_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_5_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_5_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_5_16_1  (
            .in0(N__11953),
            .in1(N__11538),
            .in2(_gnd_net_),
            .in3(N__11519),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__22024),
            .ce(N__11838),
            .sr(N__22256));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_5_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_5_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_5_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_5_16_2  (
            .in0(N__11946),
            .in1(N__11514),
            .in2(_gnd_net_),
            .in3(N__11495),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__22024),
            .ce(N__11838),
            .sr(N__22256));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_5_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_5_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_5_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_5_16_3  (
            .in0(N__11950),
            .in1(N__11490),
            .in2(_gnd_net_),
            .in3(N__11471),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__22024),
            .ce(N__11838),
            .sr(N__22256));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_5_16_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_5_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_5_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_5_16_4  (
            .in0(N__11947),
            .in1(N__11468),
            .in2(_gnd_net_),
            .in3(N__11453),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__22024),
            .ce(N__11838),
            .sr(N__22256));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_5_16_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_5_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_5_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_5_16_5  (
            .in0(N__11951),
            .in1(N__11822),
            .in2(_gnd_net_),
            .in3(N__11807),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__22024),
            .ce(N__11838),
            .sr(N__22256));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_5_16_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_5_16_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_5_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_5_16_6  (
            .in0(N__11948),
            .in1(N__11802),
            .in2(_gnd_net_),
            .in3(N__11783),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__22024),
            .ce(N__11838),
            .sr(N__22256));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_5_16_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_5_16_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_5_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_5_16_7  (
            .in0(N__11952),
            .in1(N__11778),
            .in2(_gnd_net_),
            .in3(N__11759),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__22024),
            .ce(N__11838),
            .sr(N__22256));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_5_17_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_5_17_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_5_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_5_17_0  (
            .in0(N__11954),
            .in1(N__11754),
            .in2(_gnd_net_),
            .in3(N__11735),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_5_17_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__22020),
            .ce(N__11839),
            .sr(N__22263));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_5_17_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_5_17_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_5_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_5_17_1  (
            .in0(N__11958),
            .in1(N__11730),
            .in2(_gnd_net_),
            .in3(N__11711),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__22020),
            .ce(N__11839),
            .sr(N__22263));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_5_17_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_5_17_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_5_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_5_17_2  (
            .in0(N__11955),
            .in1(N__11706),
            .in2(_gnd_net_),
            .in3(N__11687),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__22020),
            .ce(N__11839),
            .sr(N__22263));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_5_17_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_5_17_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_5_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_5_17_3  (
            .in0(N__11959),
            .in1(N__11682),
            .in2(_gnd_net_),
            .in3(N__11663),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__22020),
            .ce(N__11839),
            .sr(N__22263));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_5_17_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_5_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_5_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_5_17_4  (
            .in0(N__11956),
            .in1(N__11660),
            .in2(_gnd_net_),
            .in3(N__11645),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__22020),
            .ce(N__11839),
            .sr(N__22263));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_5_17_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_5_17_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_5_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_5_17_5  (
            .in0(N__11960),
            .in1(N__11642),
            .in2(_gnd_net_),
            .in3(N__12137),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__22020),
            .ce(N__11839),
            .sr(N__22263));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_5_17_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_5_17_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_5_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_5_17_6  (
            .in0(N__11957),
            .in1(N__12132),
            .in2(_gnd_net_),
            .in3(N__12113),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__22020),
            .ce(N__11839),
            .sr(N__22263));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_5_17_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_5_17_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_5_17_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_5_17_7  (
            .in0(N__11961),
            .in1(N__12108),
            .in2(_gnd_net_),
            .in3(N__12089),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__22020),
            .ce(N__11839),
            .sr(N__22263));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_5_18_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_5_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_5_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_5_18_0  (
            .in0(N__11962),
            .in1(N__12084),
            .in2(_gnd_net_),
            .in3(N__12065),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_5_18_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__22015),
            .ce(N__11840),
            .sr(N__22272));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_5_18_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_5_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_5_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_5_18_1  (
            .in0(N__11966),
            .in1(N__12060),
            .in2(_gnd_net_),
            .in3(N__12041),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__22015),
            .ce(N__11840),
            .sr(N__22272));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_5_18_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_5_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_5_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_5_18_2  (
            .in0(N__11963),
            .in1(N__12036),
            .in2(_gnd_net_),
            .in3(N__12017),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__22015),
            .ce(N__11840),
            .sr(N__22272));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_5_18_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_5_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_5_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_5_18_3  (
            .in0(N__11967),
            .in1(N__12012),
            .in2(_gnd_net_),
            .in3(N__11993),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__22015),
            .ce(N__11840),
            .sr(N__22272));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_5_18_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_5_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_5_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_5_18_4  (
            .in0(N__11964),
            .in1(N__11990),
            .in2(_gnd_net_),
            .in3(N__11978),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__22015),
            .ce(N__11840),
            .sr(N__22272));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_5_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_5_18_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_5_18_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_5_18_5  (
            .in0(N__11852),
            .in1(N__11965),
            .in2(_gnd_net_),
            .in3(N__11855),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22015),
            .ce(N__11840),
            .sr(N__22272));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_5_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_5_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_5_19_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_5_19_0  (
            .in0(N__15450),
            .in1(N__15350),
            .in2(_gnd_net_),
            .in3(N__14732),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22009),
            .ce(N__18499),
            .sr(N__22276));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_5_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_5_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_5_19_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_5_19_1  (
            .in0(N__15351),
            .in1(N__16147),
            .in2(_gnd_net_),
            .in3(N__15451),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22009),
            .ce(N__18499),
            .sr(N__22276));
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_5_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_5_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_5_19_5 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_5_19_5  (
            .in0(N__14565),
            .in1(N__15907),
            .in2(_gnd_net_),
            .in3(N__15576),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22009),
            .ce(N__18499),
            .sr(N__22276));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_5_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_5_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_5_19_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_5_19_7  (
            .in0(N__15349),
            .in1(N__14263),
            .in2(_gnd_net_),
            .in3(N__15449),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22009),
            .ce(N__18499),
            .sr(N__22276));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_5_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_5_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_5_20_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_5_20_0  (
            .in0(N__15412),
            .in1(N__15310),
            .in2(_gnd_net_),
            .in3(N__14399),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22002),
            .ce(N__18500),
            .sr(N__22280));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_5_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_5_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_5_20_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_5_20_5  (
            .in0(N__15309),
            .in1(N__15411),
            .in2(_gnd_net_),
            .in3(N__14509),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22002),
            .ce(N__18500),
            .sr(N__22280));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_d_0_LC_5_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_d_0_LC_5_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_d_0_LC_5_21_0 .LUT_INIT=16'b0001001110110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto31_d_0_LC_5_21_0  (
            .in0(N__12515),
            .in1(N__12184),
            .in2(N__12146),
            .in3(N__12161),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto31_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_5_21_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_5_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_5_21_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_5_21_1  (
            .in0(N__15665),
            .in1(N__12465),
            .in2(_gnd_net_),
            .in3(N__12342),
            .lcout(\phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_start_0_a0_0_LC_5_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_start_0_a0_0_LC_5_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_start_0_a0_0_LC_5_21_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_start_0_a0_0_LC_5_21_4  (
            .in0(N__18740),
            .in1(N__18710),
            .in2(N__12662),
            .in3(N__15894),
            .lcout(\phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m3_e_1_LC_5_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m3_e_1_LC_5_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m3_e_1_LC_5_21_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m3_e_1_LC_5_21_7  (
            .in0(N__15893),
            .in1(N__14393),
            .in2(_gnd_net_),
            .in3(N__14829),
            .lcout(\phase_controller_inst1.stoper_hc.un1_m3_eZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_1_LC_5_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_1_LC_5_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_1_LC_5_22_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m3_0_1_LC_5_22_0  (
            .in0(N__16009),
            .in1(N__15784),
            .in2(N__14508),
            .in3(N__15961),
            .lcout(\phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_a0_1_LC_5_22_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_a0_1_LC_5_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_a0_1_LC_5_22_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto31_a0_1_LC_5_22_1  (
            .in0(N__15884),
            .in1(N__14831),
            .in2(_gnd_net_),
            .in3(N__12514),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto31_a0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_5_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_5_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_5_22_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_5_22_2  (
            .in0(N__14333),
            .in1(N__14615),
            .in2(N__14458),
            .in3(N__14874),
            .lcout(phase_controller_inst1_stoper_hc_un1_startlto19_2),
            .ltout(phase_controller_inst1_stoper_hc_un1_startlto19_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_1_RNIQA9D_15_LC_5_22_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_1_RNIQA9D_15_LC_5_22_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_1_RNIQA9D_15_LC_5_22_3 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_1_RNIQA9D_15_LC_5_22_3  (
            .in0(_gnd_net_),
            .in1(N__15882),
            .in2(N__12503),
            .in3(N__14392),
            .lcout(d_N_5_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_5_22_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_5_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_5_22_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_5_22_4  (
            .in0(N__15698),
            .in1(N__12466),
            .in2(_gnd_net_),
            .in3(N__12343),
            .lcout(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_a2_LC_5_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_a2_LC_5_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_a2_LC_5_22_5 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto31_a2_LC_5_22_5  (
            .in0(N__12655),
            .in1(N__18736),
            .in2(N__18709),
            .in3(N__15883),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto31_aZ0Z2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_1_LC_5_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_1_LC_5_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto31_1_LC_5_22_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto31_1_LC_5_22_6  (
            .in0(N__12194),
            .in1(N__12160),
            .in2(N__12188),
            .in3(N__12185),
            .lcout(\phase_controller_inst1.stoper_hc.un1_start ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_2_LC_5_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_2_LC_5_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_2_LC_5_23_0 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m3_0_2_LC_5_23_0  (
            .in0(N__16138),
            .in1(N__16045),
            .in2(N__16196),
            .in3(N__12173),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_LC_5_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_LC_5_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m3_0_LC_5_23_1 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m3_0_LC_5_23_1  (
            .in0(N__14554),
            .in1(N__16194),
            .in2(N__12164),
            .in3(N__12677),
            .lcout(\phase_controller_inst1.stoper_hc.un1_N_6_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_3_LC_5_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_3_LC_5_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_3_LC_5_23_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m2_e_3_LC_5_23_2  (
            .in0(N__14252),
            .in1(N__14651),
            .in2(N__14730),
            .in3(N__14121),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_LC_5_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_LC_5_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_m2_e_LC_5_23_3 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_m2_e_LC_5_23_3  (
            .in0(N__14206),
            .in1(_gnd_net_),
            .in2(N__12680),
            .in3(N__16094),
            .lcout(\phase_controller_inst1.stoper_hc.un1_m2_eZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_5_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_5_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_5_23_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_5_23_4  (
            .in0(N__16190),
            .in1(N__14684),
            .in2(_gnd_net_),
            .in3(N__14617),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_5_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_5_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_5_23_5 .LUT_INIT=16'b0011000001110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_5_23_5  (
            .in0(N__14207),
            .in1(N__14652),
            .in2(N__12671),
            .in3(N__16095),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_0_LC_5_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_0_LC_5_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_0_LC_5_23_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_0_LC_5_23_6  (
            .in0(N__14149),
            .in1(N__14170),
            .in2(_gnd_net_),
            .in3(N__14683),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto30_2_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_5_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_5_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_5_23_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_5_23_7  (
            .in0(N__14171),
            .in1(N__14828),
            .in2(N__14397),
            .in3(N__14150),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_4.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_4 (
            .in0(N__12638),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_7_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_7_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_7_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_7_12_2  (
            .in0(N__12923),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12610),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22034),
            .ce(N__19944),
            .sr(N__22233));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_7_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_7_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_7_12_3 .LUT_INIT=16'b1111001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_7_12_3  (
            .in0(N__20032),
            .in1(N__12926),
            .in2(N__12587),
            .in3(N__12548),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22034),
            .ce(N__19944),
            .sr(N__22233));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_7_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_7_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_7_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_7_12_4  (
            .in0(N__12924),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13015),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22034),
            .ce(N__19944),
            .sr(N__22233));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_7_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_7_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_7_12_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__12925),
            .in2(_gnd_net_),
            .in3(N__12995),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22034),
            .ce(N__19944),
            .sr(N__22233));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_7_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_7_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_7_12_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_7_12_6  (
            .in0(N__20128),
            .in1(N__20031),
            .in2(_gnd_net_),
            .in3(N__12962),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22034),
            .ce(N__19944),
            .sr(N__22233));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_7_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_7_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_7_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(N__12922),
            .in2(_gnd_net_),
            .in3(N__12880),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22034),
            .ce(N__19944),
            .sr(N__22233));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_7_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_7_13_0 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_7_13_0  (
            .in0(N__13138),
            .in1(N__20118),
            .in2(N__13234),
            .in3(N__12856),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22029),
            .ce(N__19949),
            .sr(N__22237));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_7_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_7_13_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_7_13_1  (
            .in0(N__12827),
            .in1(N__20116),
            .in2(_gnd_net_),
            .in3(N__13136),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22029),
            .ce(N__19949),
            .sr(N__22237));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_7_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_7_13_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_7_13_2  (
            .in0(N__13137),
            .in1(N__20117),
            .in2(_gnd_net_),
            .in3(N__12782),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22029),
            .ce(N__19949),
            .sr(N__22237));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_7_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_7_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_7_13_3 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_7_13_3  (
            .in0(N__20119),
            .in1(N__12743),
            .in2(N__13233),
            .in3(N__13139),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22029),
            .ce(N__19949),
            .sr(N__22237));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_7_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_7_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_7_13_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_7_13_4  (
            .in0(N__12719),
            .in1(N__13289),
            .in2(N__12701),
            .in3(N__13264),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22029),
            .ce(N__19949),
            .sr(N__22237));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_7_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_7_13_5 .LUT_INIT=16'b1000101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_7_13_5  (
            .in0(N__13263),
            .in1(N__13337),
            .in2(N__13301),
            .in3(N__13358),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22029),
            .ce(N__19949),
            .sr(N__22237));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_7_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_7_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_7_13_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_7_13_6  (
            .in0(N__13336),
            .in1(N__13293),
            .in2(_gnd_net_),
            .in3(N__13265),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22029),
            .ce(N__19949),
            .sr(N__22237));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_7_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_7_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_7_13_7 .LUT_INIT=16'b0011000000110001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_7_13_7  (
            .in0(N__20120),
            .in1(N__13224),
            .in2(N__13187),
            .in3(N__13140),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22029),
            .ce(N__19949),
            .sr(N__22237));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_7_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_7_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__13100),
            .in2(N__13094),
            .in3(N__17067),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_7_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_7_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__13085),
            .in2(N__13076),
            .in3(N__17035),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_7_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_7_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__13067),
            .in2(N__13061),
            .in3(N__17014),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_7_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_7_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__13052),
            .in2(N__13046),
            .in3(N__16981),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_7_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_7_14_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_7_14_4  (
            .in0(N__16960),
            .in1(N__13037),
            .in2(N__13028),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_7_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_7_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__13487),
            .in2(N__13481),
            .in3(N__16939),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_7_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_7_14_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_7_14_6  (
            .in0(N__17290),
            .in1(N__13472),
            .in2(N__13466),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_7_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_7_14_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_7_14_7  (
            .in0(N__17269),
            .in1(N__13457),
            .in2(N__13448),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_7_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_7_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__13439),
            .in2(N__13430),
            .in3(N__17248),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_7_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_7_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__13421),
            .in2(N__13412),
            .in3(N__17227),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_7_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_7_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__13403),
            .in2(N__13394),
            .in3(N__17203),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_7_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_7_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__13385),
            .in2(N__13376),
            .in3(N__17183),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_7_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_7_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__13367),
            .in2(N__13565),
            .in3(N__17155),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_7_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_7_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(N__13556),
            .in2(N__13547),
            .in3(N__17131),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_7_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_7_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(N__19961),
            .in2(N__13538),
            .in3(N__17668),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_7_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_7_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(N__13616),
            .in2(N__13529),
            .in3(N__17644),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_7_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_7_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__13697),
            .in2(N__13520),
            .in3(N__17623),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_7_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_7_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__13658),
            .in2(N__13511),
            .in3(N__17602),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_7_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_7_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(N__13739),
            .in2(N__13502),
            .in3(N__17581),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13493),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_16_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13490),
            .in3(N__19734),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_7_16_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_7_16_6 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_7_16_6  (
            .in0(N__15237),
            .in1(_gnd_net_),
            .in2(N__15008),
            .in3(N__19789),
            .lcout(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_7_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_7_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_7_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13782),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22010),
            .ce(N__19929),
            .sr(N__22250));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_7_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_7_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_7_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13733),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22010),
            .ce(N__19929),
            .sr(N__22250));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_7_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_7_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_7_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13691),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22010),
            .ce(N__19929),
            .sr(N__22250));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_7_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_7_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_7_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13652),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22010),
            .ce(N__19929),
            .sr(N__22250));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_7_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_7_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_7_18_0 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_7_18_0  (
            .in0(N__15903),
            .in1(N__13606),
            .in2(N__14221),
            .in3(N__15586),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22003),
            .ce(N__18487),
            .sr(N__22257));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_7_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_7_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_7_18_4 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_7_18_4  (
            .in0(N__15904),
            .in1(N__15587),
            .in2(N__14666),
            .in3(N__13607),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22003),
            .ce(N__18487),
            .sr(N__22257));
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_7_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_7_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_7_18_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_0_LC_7_18_5  (
            .in0(N__13604),
            .in1(N__14122),
            .in2(N__15373),
            .in3(N__15466),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22003),
            .ce(N__18487),
            .sr(N__22257));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_7_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_7_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_7_18_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_7_18_7  (
            .in0(N__13605),
            .in1(N__16102),
            .in2(N__15374),
            .in3(N__15467),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22003),
            .ce(N__18487),
            .sr(N__22257));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_7_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_7_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13949),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_7_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_7_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__13940),
            .in2(N__13934),
            .in3(N__18414),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_7_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_7_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__13925),
            .in2(N__13919),
            .in3(N__17311),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_7_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_7_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__13910),
            .in2(N__13904),
            .in3(N__17866),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_7_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_7_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__13895),
            .in2(N__13886),
            .in3(N__17827),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_7_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_7_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__13877),
            .in2(N__13868),
            .in3(N__17806),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_7_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_7_19_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_7_19_6  (
            .in0(N__17785),
            .in1(N__13859),
            .in2(N__13850),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_7_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_7_19_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_7_19_7  (
            .in0(N__17764),
            .in1(N__13841),
            .in2(N__13832),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_7_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_7_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_7_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__15473),
            .in2(N__14042),
            .in3(N__17737),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_7_20_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_7_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_7_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(N__15497),
            .in2(N__14033),
            .in3(N__17710),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_7_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_7_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(N__15491),
            .in2(N__14024),
            .in3(N__17689),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_7_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_7_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(N__15482),
            .in2(N__14015),
            .in3(N__18031),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_7_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_7_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_7_20_4  (
            .in0(_gnd_net_),
            .in1(N__15269),
            .in2(N__14006),
            .in3(N__18010),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_7_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_7_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_7_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(N__13997),
            .in2(N__13988),
            .in3(N__17989),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_7_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_7_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_7_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(N__14279),
            .in2(N__13979),
            .in3(N__17968),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_7_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_7_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_7_20_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_7_20_7  (
            .in0(N__17947),
            .in1(N__13970),
            .in2(N__13958),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_7_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_7_21_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_7_21_0  (
            .in0(N__17927),
            .in1(N__14048),
            .in2(N__14090),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_7_21_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_7_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_7_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__14288),
            .in2(N__14081),
            .in3(N__17902),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_7_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_7_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(N__14297),
            .in2(N__14072),
            .in3(N__17878),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_7_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_7_21_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_7_21_3  (
            .in0(N__18520),
            .in1(N__14270),
            .in2(N__14063),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14054),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(N__18438),
            .in2(_gnd_net_),
            .in3(N__18387),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_7_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_7_21_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(N__18267),
            .in2(_gnd_net_),
            .in3(N__18163),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed11 ),
            .ltout(\phase_controller_inst1.stoper_hc.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_7_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_7_21_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_7_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14051),
            .in3(N__18388),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_7_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_7_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_7_22_2 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_7_22_2  (
            .in0(N__15873),
            .in1(N__14873),
            .in2(_gnd_net_),
            .in3(N__15559),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21985),
            .ce(N__18491),
            .sr(N__22281));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_7_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_7_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_7_22_3 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_7_22_3  (
            .in0(N__15561),
            .in1(N__15875),
            .in2(_gnd_net_),
            .in3(N__14337),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21985),
            .ce(N__18491),
            .sr(N__22281));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_7_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_7_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_7_22_4 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_7_22_4  (
            .in0(N__15874),
            .in1(N__14614),
            .in2(_gnd_net_),
            .in3(N__15560),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21985),
            .ce(N__18491),
            .sr(N__22281));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_7_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_7_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_7_22_6 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_7_22_6  (
            .in0(N__15872),
            .in1(N__14824),
            .in2(_gnd_net_),
            .in3(N__15558),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21985),
            .ce(N__18491),
            .sr(N__22281));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_7_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_7_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_7_22_7 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_7_22_7  (
            .in0(N__15562),
            .in1(N__15876),
            .in2(_gnd_net_),
            .in3(N__14449),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21985),
            .ce(N__18491),
            .sr(N__22281));
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_7_23_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_7_23_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_7_23_0 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_4_LC_7_23_0  (
            .in0(N__14251),
            .in1(N__19104),
            .in2(N__16277),
            .in3(N__18611),
            .lcout(measured_delay_hc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21982),
            .ce(),
            .sr(N__22286));
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_7_23_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_7_23_1 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_7_23_1 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_1_LC_7_23_1  (
            .in0(N__19102),
            .in1(N__18914),
            .in2(N__14214),
            .in3(N__18990),
            .lcout(measured_delay_hc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21982),
            .ce(),
            .sr(N__22286));
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_7_23_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_7_23_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_7_23_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_22_LC_7_23_2  (
            .in0(N__18993),
            .in1(N__14169),
            .in2(_gnd_net_),
            .in3(N__19101),
            .lcout(measured_delay_hc_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21982),
            .ce(),
            .sr(N__22286));
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_7_23_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_7_23_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_7_23_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_21_LC_7_23_3  (
            .in0(N__19100),
            .in1(N__14148),
            .in2(_gnd_net_),
            .in3(N__18992),
            .lcout(measured_delay_hc_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21982),
            .ce(),
            .sr(N__22286));
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_7_23_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_7_23_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_7_23_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_0_LC_7_23_4  (
            .in0(N__14120),
            .in1(N__19098),
            .in2(_gnd_net_),
            .in3(N__18610),
            .lcout(measured_delay_hc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21982),
            .ce(),
            .sr(N__22286));
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_7_23_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_7_23_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_7_23_5 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_5_LC_7_23_5  (
            .in0(N__19105),
            .in1(N__16606),
            .in2(N__14729),
            .in3(N__18995),
            .lcout(measured_delay_hc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21982),
            .ce(),
            .sr(N__22286));
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_7_23_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_7_23_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_7_23_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_20_LC_7_23_6  (
            .in0(N__18991),
            .in1(N__14682),
            .in2(_gnd_net_),
            .in3(N__19099),
            .lcout(measured_delay_hc_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21982),
            .ce(),
            .sr(N__22286));
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_7_23_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_7_23_7 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_7_23_7 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_3_LC_7_23_7  (
            .in0(N__19103),
            .in1(N__14650),
            .in2(N__16304),
            .in3(N__18994),
            .lcout(measured_delay_hc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21982),
            .ce(),
            .sr(N__22286));
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_7_24_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_7_24_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_7_24_0 .LUT_INIT=16'b1110111011111010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_17_LC_7_24_0  (
            .in0(N__18603),
            .in1(N__16721),
            .in2(N__14618),
            .in3(N__19110),
            .lcout(measured_delay_hc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21979),
            .ce(),
            .sr(N__22291));
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_7_24_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_7_24_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_7_24_1 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_6_LC_7_24_1  (
            .in0(N__19113),
            .in1(N__16577),
            .in2(N__14558),
            .in3(N__18606),
            .lcout(measured_delay_hc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21979),
            .ce(),
            .sr(N__22291));
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_7_24_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_7_24_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_7_24_2 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_13_LC_7_24_2  (
            .in0(N__16400),
            .in1(N__19106),
            .in2(N__14497),
            .in3(N__18983),
            .lcout(measured_delay_hc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21979),
            .ce(),
            .sr(N__22291));
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_7_24_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_7_24_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_7_24_3 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_19_LC_7_24_3  (
            .in0(N__19112),
            .in1(N__16667),
            .in2(N__14450),
            .in3(N__18605),
            .lcout(measured_delay_hc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21979),
            .ce(),
            .sr(N__22291));
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_7_24_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_7_24_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_7_24_4 .LUT_INIT=16'b1011100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_15_LC_7_24_4  (
            .in0(N__16798),
            .in1(N__19108),
            .in2(N__14385),
            .in3(N__18984),
            .lcout(measured_delay_hc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21979),
            .ce(),
            .sr(N__22291));
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_7_24_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_7_24_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_7_24_5 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_18_LC_7_24_5  (
            .in0(N__19111),
            .in1(N__16694),
            .in2(N__14332),
            .in3(N__18604),
            .lcout(measured_delay_hc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21979),
            .ce(),
            .sr(N__22291));
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_7_24_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_7_24_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_7_24_6 .LUT_INIT=16'b1111101011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_16_LC_7_24_6  (
            .in0(N__18602),
            .in1(N__14863),
            .in2(N__16751),
            .in3(N__19109),
            .lcout(measured_delay_hc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21979),
            .ce(),
            .sr(N__22291));
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_7_24_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_7_24_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_7_24_7 .LUT_INIT=16'b1111111111100100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_14_LC_7_24_7  (
            .in0(N__19107),
            .in1(N__14814),
            .in2(N__16838),
            .in3(N__18601),
            .lcout(measured_delay_hc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21979),
            .ce(),
            .sr(N__22291));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_14_LC_7_25_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_14_LC_7_25_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_14_LC_7_25_3 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_14_LC_7_25_3  (
            .in0(N__16322),
            .in1(N__14774),
            .in2(N__14762),
            .in3(N__14741),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_13_LC_7_26_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_13_LC_7_26_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_13_LC_7_26_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_13_LC_7_26_3  (
            .in0(N__16596),
            .in1(N__16263),
            .in2(N__16746),
            .in3(N__16392),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU0I2_19_LC_7_26_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU0I2_19_LC_7_26_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU0I2_19_LC_7_26_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU0I2_19_LC_7_26_4  (
            .in0(N__16662),
            .in1(N__16573),
            .in2(N__14777),
            .in3(N__14768),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_7_26_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_7_26_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_7_26_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_7_26_6  (
            .in0(_gnd_net_),
            .in1(N__16683),
            .in2(_gnd_net_),
            .in3(N__16710),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_7_28_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_7_28_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_7_28_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_7_28_1  (
            .in0(N__16619),
            .in1(N__17083),
            .in2(N__16919),
            .in3(N__16633),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_7_28_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_7_28_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_7_28_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_7_28_3  (
            .in0(N__14909),
            .in1(N__14750),
            .in2(N__16637),
            .in3(N__14903),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_7_28_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_7_28_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_7_28_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_7_28_4  (
            .in0(N__16886),
            .in1(N__16895),
            .in2(N__16877),
            .in3(N__16904),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_23_LC_7_28_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_23_LC_7_28_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_23_LC_7_28_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_23_LC_7_28_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14744),
            .in3(N__14902),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_7_28_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_7_28_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_7_28_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_7_28_6  (
            .in0(_gnd_net_),
            .in1(N__16915),
            .in2(_gnd_net_),
            .in3(N__16618),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_7_29_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_7_29_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_7_29_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_7_29_6  (
            .in0(N__16847),
            .in1(N__16856),
            .in2(N__17111),
            .in3(N__16865),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_12_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_12_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_8_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14894),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22030),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_8_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_8_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_8_13_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_8_13_0  (
            .in0(N__17543),
            .in1(N__17431),
            .in2(N__20846),
            .in3(N__17258),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22025),
            .ce(),
            .sr(N__22234));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_8_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_8_13_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_8_13_1  (
            .in0(N__17426),
            .in1(N__20825),
            .in2(N__17559),
            .in3(N__16949),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22025),
            .ce(),
            .sr(N__22234));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_8_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_8_13_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_8_13_2  (
            .in0(N__17542),
            .in1(N__17430),
            .in2(N__20845),
            .in3(N__16970),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22025),
            .ce(),
            .sr(N__22234));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_8_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_8_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_8_13_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_8_13_3  (
            .in0(N__17428),
            .in1(N__20827),
            .in2(N__17561),
            .in3(N__17279),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22025),
            .ce(),
            .sr(N__22234));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_8_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_8_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_8_13_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_8_13_4  (
            .in0(N__17541),
            .in1(N__17429),
            .in2(N__20844),
            .in3(N__17024),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22025),
            .ce(),
            .sr(N__22234));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_8_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_8_13_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_8_13_5  (
            .in0(N__17427),
            .in1(N__20826),
            .in2(N__17560),
            .in3(N__16928),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22025),
            .ce(),
            .sr(N__22234));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_8_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_8_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_8_13_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_8_13_7  (
            .in0(N__17425),
            .in1(N__20824),
            .in2(N__17558),
            .in3(N__16991),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22025),
            .ce(),
            .sr(N__22234));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_8_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_8_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_8_14_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_8_14_0  (
            .in0(N__17403),
            .in1(N__17532),
            .in2(N__20840),
            .in3(N__17237),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22021),
            .ce(),
            .sr(N__22238));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_8_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_8_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_8_14_1 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_8_14_1  (
            .in0(N__17525),
            .in1(N__20808),
            .in2(N__17216),
            .in3(N__17404),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22021),
            .ce(),
            .sr(N__22238));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_8_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_8_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_8_14_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_8_14_2  (
            .in0(N__17401),
            .in1(N__17530),
            .in2(N__20838),
            .in3(N__17165),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22021),
            .ce(),
            .sr(N__22238));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_8_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_8_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_8_14_3 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_8_14_3  (
            .in0(N__17527),
            .in1(N__20810),
            .in2(N__17657),
            .in3(N__17406),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22021),
            .ce(),
            .sr(N__22238));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_8_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_8_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_8_14_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_8_14_4  (
            .in0(N__17400),
            .in1(N__17529),
            .in2(N__20837),
            .in3(N__17192),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22021),
            .ce(),
            .sr(N__22238));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_8_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_8_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_8_14_5 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_8_14_5  (
            .in0(N__17528),
            .in1(N__20811),
            .in2(N__17435),
            .in3(N__17633),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22021),
            .ce(),
            .sr(N__22238));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_8_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_8_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_8_14_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_8_14_6  (
            .in0(N__17402),
            .in1(N__17531),
            .in2(N__20839),
            .in3(N__17120),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22021),
            .ce(),
            .sr(N__22238));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_8_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_8_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_8_14_7 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_8_14_7  (
            .in0(N__17526),
            .in1(N__20809),
            .in2(N__17144),
            .in3(N__17405),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22021),
            .ce(),
            .sr(N__22238));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_8_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_8_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_8_15_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_8_15_1  (
            .in0(N__17394),
            .in1(N__20813),
            .in2(N__17556),
            .in3(N__17591),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22016),
            .ce(),
            .sr(N__22239));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_8_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_8_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_8_15_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_8_15_2  (
            .in0(N__17540),
            .in1(N__17397),
            .in2(N__20842),
            .in3(N__14927),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22016),
            .ce(),
            .sr(N__22239));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_8_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_8_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_8_15_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_8_15_3  (
            .in0(N__17395),
            .in1(N__20814),
            .in2(N__17557),
            .in3(N__17567),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22016),
            .ce(),
            .sr(N__22239));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_8_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_8_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_8_15_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_8_15_4  (
            .in0(N__17539),
            .in1(N__17396),
            .in2(N__20841),
            .in3(N__17612),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22016),
            .ce(),
            .sr(N__22239));
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_8_15_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_8_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_8_15_7 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_LC_8_15_7  (
            .in0(N__20487),
            .in1(N__14960),
            .in2(N__14918),
            .in3(N__15122),
            .lcout(\phase_controller_slave.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22016),
            .ce(),
            .sr(N__22239));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_8_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_8_16_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_8_16_2  (
            .in0(N__20779),
            .in1(N__17470),
            .in2(_gnd_net_),
            .in3(N__17371),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_8_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_8_16_3 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_8_16_3  (
            .in0(N__19735),
            .in1(N__19706),
            .in2(_gnd_net_),
            .in3(N__17071),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_8_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_8_16_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(N__17469),
            .in2(_gnd_net_),
            .in3(N__17370),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed11 ),
            .ltout(\phase_controller_inst1.stoper_tr.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_8_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_8_16_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14921),
            .in3(N__19705),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_8_16_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_8_16_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_8_16_6  (
            .in0(N__19790),
            .in1(N__14997),
            .in2(_gnd_net_),
            .in3(N__15238),
            .lcout(\phase_controller_slave.stoper_tr.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_8_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_8_16_7 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_8_16_7  (
            .in0(N__17372),
            .in1(_gnd_net_),
            .in2(N__17508),
            .in3(N__20780),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_8_17_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_8_17_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_8_17_4 .LUT_INIT=16'b0010000001100100;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_1_LC_8_17_4  (
            .in0(N__15001),
            .in1(N__15258),
            .in2(N__19873),
            .in3(N__15118),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22004),
            .ce(N__21331),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_8_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_8_17_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_8_17_5 .LUT_INIT=16'b0010000001100100;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_1_LC_8_17_5  (
            .in0(N__17506),
            .in1(N__17399),
            .in2(N__20843),
            .in3(N__19713),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22004),
            .ce(N__21331),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_18_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_18_0  (
            .in0(N__18232),
            .in1(N__20634),
            .in2(N__18350),
            .in3(N__17753),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21997),
            .ce(),
            .sr(N__22251));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_18_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_18_1  (
            .in0(N__18337),
            .in1(N__18235),
            .in2(N__20657),
            .in3(N__17774),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21997),
            .ce(),
            .sr(N__22251));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_18_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_18_3  (
            .in0(N__18336),
            .in1(N__18234),
            .in2(N__20656),
            .in3(N__17795),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21997),
            .ce(),
            .sr(N__22251));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_18_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_18_4  (
            .in0(N__18231),
            .in1(N__20633),
            .in2(N__18349),
            .in3(N__17816),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21997),
            .ce(),
            .sr(N__22251));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_18_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_18_5  (
            .in0(N__18335),
            .in1(N__18233),
            .in2(N__20655),
            .in3(N__17300),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21997),
            .ce(),
            .sr(N__22251));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_18_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_18_6  (
            .in0(N__18230),
            .in1(N__20632),
            .in2(N__18348),
            .in3(N__17837),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21997),
            .ce(),
            .sr(N__22251));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_19_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_19_0  (
            .in0(N__18328),
            .in1(N__18227),
            .in2(N__20646),
            .in3(N__17957),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21993),
            .ce(),
            .sr(N__22258));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_19_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_19_1  (
            .in0(N__18223),
            .in1(N__18332),
            .in2(N__20652),
            .in3(N__18020),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21993),
            .ce(),
            .sr(N__22258));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_19_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_19_2  (
            .in0(N__18329),
            .in1(N__18228),
            .in2(N__20647),
            .in3(N__17936),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21993),
            .ce(),
            .sr(N__22258));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_19_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_19_3  (
            .in0(N__18225),
            .in1(N__18334),
            .in2(N__20654),
            .in3(N__17912),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21993),
            .ce(),
            .sr(N__22258));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_19_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_19_4  (
            .in0(N__18330),
            .in1(N__18229),
            .in2(N__20648),
            .in3(N__17699),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21993),
            .ce(),
            .sr(N__22258));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_19_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_19_5  (
            .in0(N__18222),
            .in1(N__18331),
            .in2(N__20651),
            .in3(N__17678),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21993),
            .ce(),
            .sr(N__22258));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_19_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_19_6  (
            .in0(N__18327),
            .in1(N__18226),
            .in2(N__20645),
            .in3(N__17999),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21993),
            .ce(),
            .sr(N__22258));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_19_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_19_7  (
            .in0(N__18224),
            .in1(N__18333),
            .in2(N__20653),
            .in3(N__17978),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21993),
            .ce(),
            .sr(N__22258));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_20_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_20_0  (
            .in0(N__18218),
            .in1(N__18325),
            .in2(N__20650),
            .in3(N__18506),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21990),
            .ce(),
            .sr(N__22264));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_20_1 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_20_1  (
            .in0(N__18324),
            .in1(N__20616),
            .in2(N__17726),
            .in3(N__18221),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21990),
            .ce(),
            .sr(N__22264));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_8_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_8_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_8_20_3 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_8_20_3  (
            .in0(N__20403),
            .in1(N__18442),
            .in2(N__18134),
            .in3(N__18394),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21990),
            .ce(),
            .sr(N__22264));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_20_4 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_20_4  (
            .in0(N__18217),
            .in1(N__20611),
            .in2(N__18533),
            .in3(N__18326),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21990),
            .ce(),
            .sr(N__22264));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_20_5 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_20_5  (
            .in0(N__18322),
            .in1(N__20615),
            .in2(N__17891),
            .in3(N__18220),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21990),
            .ce(),
            .sr(N__22264));
    defparam \phase_controller_slave.start_timer_hc_LC_8_20_6 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_LC_8_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_hc_LC_8_20_6 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \phase_controller_slave.start_timer_hc_LC_8_20_6  (
            .in0(N__15633),
            .in1(N__18356),
            .in2(N__20348),
            .in3(N__18125),
            .lcout(\phase_controller_slave.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21990),
            .ce(),
            .sr(N__22264));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_20_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_20_7  (
            .in0(N__18323),
            .in1(N__18219),
            .in2(N__20649),
            .in3(N__18362),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21990),
            .ce(),
            .sr(N__22264));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_8_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_8_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_8_21_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_8_21_0  (
            .in0(N__15871),
            .in1(N__16186),
            .in2(_gnd_net_),
            .in3(N__15577),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21986),
            .ce(N__18492),
            .sr(N__22273));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_8_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_8_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_8_21_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_8_21_1  (
            .in0(N__15358),
            .in1(N__15960),
            .in2(_gnd_net_),
            .in3(N__15462),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21986),
            .ce(N__18492),
            .sr(N__22273));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_8_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_8_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_8_21_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_8_21_2  (
            .in0(N__15463),
            .in1(N__15359),
            .in2(_gnd_net_),
            .in3(N__15779),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21986),
            .ce(N__18492),
            .sr(N__22273));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_8_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_8_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_8_21_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_8_21_3  (
            .in0(N__15361),
            .in1(N__16055),
            .in2(_gnd_net_),
            .in3(N__15465),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21986),
            .ce(N__18492),
            .sr(N__22273));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_8_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_8_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_8_21_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_8_21_6  (
            .in0(N__15464),
            .in1(N__15360),
            .in2(_gnd_net_),
            .in3(N__16007),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21986),
            .ce(N__18492),
            .sr(N__22273));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_8_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_8_22_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_8_22_4 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_0_LC_8_22_4  (
            .in0(N__18316),
            .in1(N__18211),
            .in2(N__20644),
            .in3(N__18392),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21983),
            .ce(N__21324),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_8_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_8_22_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_8_22_7 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_1_LC_8_22_7  (
            .in0(N__18393),
            .in1(N__20595),
            .in2(N__18236),
            .in3(N__18317),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21983),
            .ce(N__21324),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_8_23_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_8_23_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_8_23_0 .LUT_INIT=16'b1111010111011101;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_9_LC_8_23_0  (
            .in0(N__18982),
            .in1(N__16185),
            .in2(N__16508),
            .in3(N__19097),
            .lcout(measured_delay_hc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21980),
            .ce(),
            .sr(N__22282));
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_8_23_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_8_23_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_8_23_1 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_7_LC_8_23_1  (
            .in0(N__19095),
            .in1(N__18980),
            .in2(N__16146),
            .in3(N__16553),
            .lcout(measured_delay_hc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21980),
            .ce(),
            .sr(N__22282));
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_8_23_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_8_23_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_8_23_2 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_2_LC_8_23_2  (
            .in0(N__18979),
            .in1(N__16093),
            .in2(N__18896),
            .in3(N__19094),
            .lcout(measured_delay_hc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21980),
            .ce(),
            .sr(N__22282));
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_8_23_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_8_23_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_8_23_3 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_8_LC_8_23_3  (
            .in0(N__19096),
            .in1(N__16532),
            .in2(N__16060),
            .in3(N__18981),
            .lcout(measured_delay_hc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21980),
            .ce(),
            .sr(N__22282));
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_8_23_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_8_23_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_8_23_4 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_12_LC_8_23_4  (
            .in0(N__18599),
            .in1(N__19093),
            .in2(N__16008),
            .in3(N__16427),
            .lcout(measured_delay_hc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21980),
            .ce(),
            .sr(N__22282));
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_8_23_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_8_23_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_8_23_5 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_10_LC_8_23_5  (
            .in0(N__16472),
            .in1(N__15952),
            .in2(N__19118),
            .in3(N__18978),
            .lcout(measured_delay_hc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21980),
            .ce(),
            .sr(N__22282));
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_8_23_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_8_23_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_8_23_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_31_LC_8_23_6  (
            .in0(N__18600),
            .in1(N__15838),
            .in2(_gnd_net_),
            .in3(N__19088),
            .lcout(measured_delay_hc_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21980),
            .ce(),
            .sr(N__22282));
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_8_23_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_8_23_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_8_23_7 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_11_LC_8_23_7  (
            .in0(N__19092),
            .in1(N__18598),
            .in2(N__15783),
            .in3(N__16451),
            .lcout(measured_delay_hc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21980),
            .ce(),
            .sr(N__22282));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINHL3C_0_31_LC_8_24_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINHL3C_0_31_LC_8_24_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINHL3C_0_31_LC_8_24_0 .LUT_INIT=16'b0000110100000101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINHL3C_0_31_LC_8_24_0  (
            .in0(N__16216),
            .in1(N__16366),
            .in2(N__17096),
            .in3(N__16226),
            .lcout(\delay_measurement_inst.delay_hc_reg3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5FBM1_9_LC_8_24_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5FBM1_9_LC_8_24_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5FBM1_9_LC_8_24_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5FBM1_9_LC_8_24_1  (
            .in0(N__16346),
            .in1(N__16503),
            .in2(_gnd_net_),
            .in3(N__16795),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5FBM1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_8_24_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_8_24_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_8_24_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_8_24_2  (
            .in0(N__16796),
            .in1(N__16832),
            .in2(_gnd_net_),
            .in3(N__16316),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIABFQE_14_LC_8_24_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIABFQE_14_LC_8_24_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIABFQE_14_LC_8_24_3 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIABFQE_14_LC_8_24_3  (
            .in0(N__16247),
            .in1(N__16202),
            .in2(N__16241),
            .in3(N__16238),
            .lcout(\delay_measurement_inst.un1_elapsed_time_hc ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_8_24_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_8_24_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_8_24_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_8_24_4  (
            .in0(N__18907),
            .in1(N__16300),
            .in2(N__16607),
            .in3(N__18888),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FS83_4_LC_8_24_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FS83_4_LC_8_24_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FS83_4_LC_8_24_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FS83_4_LC_8_24_5  (
            .in0(N__16270),
            .in1(N__16793),
            .in2(N__16232),
            .in3(N__16358),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9U7V4_9_LC_8_24_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9U7V4_9_LC_8_24_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9U7V4_9_LC_8_24_6 .LUT_INIT=16'b0000111011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9U7V4_9_LC_8_24_6  (
            .in0(N__16794),
            .in1(N__16507),
            .in2(N__16229),
            .in3(N__16345),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINHL3C_31_LC_8_24_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINHL3C_31_LC_8_24_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINHL3C_31_LC_8_24_7 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINHL3C_31_LC_8_24_7  (
            .in0(N__16367),
            .in1(N__17095),
            .in2(N__16220),
            .in3(N__16217),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2_6_LC_8_25_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2_6_LC_8_25_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2_6_LC_8_25_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2_6_LC_8_25_0  (
            .in0(N__16572),
            .in1(N__16344),
            .in2(N__16799),
            .in3(N__16357),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2Z0Z_6 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIEHL24_14_LC_8_25_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIEHL24_14_LC_8_25_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIEHL24_14_LC_8_25_1 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIEHL24_14_LC_8_25_1  (
            .in0(N__16315),
            .in1(N__16834),
            .in2(N__16370),
            .in3(N__16792),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_25_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_25_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_25_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_25_2  (
            .in0(_gnd_net_),
            .in1(N__16524),
            .in2(_gnd_net_),
            .in3(N__16548),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_25_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_25_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_25_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_25_3  (
            .in0(N__16425),
            .in1(N__16449),
            .in2(N__16399),
            .in3(N__16467),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7KIH1_10_LC_8_25_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7KIH1_10_LC_8_25_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7KIH1_10_LC_8_25_4 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7KIH1_10_LC_8_25_4  (
            .in0(N__16468),
            .in1(N__16293),
            .in2(N__18892),
            .in3(N__16493),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_11_LC_8_25_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_11_LC_8_25_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_11_LC_8_25_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_11_LC_8_25_5  (
            .in0(N__16549),
            .in1(N__16426),
            .in2(N__16531),
            .in3(N__16450),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2ALD3_14_LC_8_25_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2ALD3_14_LC_8_25_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2ALD3_14_LC_8_25_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2ALD3_14_LC_8_25_6  (
            .in0(N__16331),
            .in1(N__16833),
            .in2(N__16325),
            .in3(N__16797),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_25_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_25_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_25_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_25_7  (
            .in0(N__16690),
            .in1(N__16747),
            .in2(N__16666),
            .in3(N__16717),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_26_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_26_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_26_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_26_0  (
            .in0(_gnd_net_),
            .in1(N__18847),
            .in2(N__18805),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_8_26_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__21973),
            .ce(N__18868),
            .sr(N__22295));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_26_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_26_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_26_1  (
            .in0(_gnd_net_),
            .in1(N__18826),
            .in2(N__18781),
            .in3(N__16250),
            .lcout(\delay_measurement_inst.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__21973),
            .ce(N__18868),
            .sr(N__22295));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_26_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_26_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_26_2  (
            .in0(_gnd_net_),
            .in1(N__18756),
            .in2(N__18806),
            .in3(N__16580),
            .lcout(\delay_measurement_inst.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__21973),
            .ce(N__18868),
            .sr(N__22295));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_26_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_26_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_26_3  (
            .in0(_gnd_net_),
            .in1(N__19314),
            .in2(N__18782),
            .in3(N__16556),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__21973),
            .ce(N__18868),
            .sr(N__22295));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_26_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_26_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_26_4  (
            .in0(_gnd_net_),
            .in1(N__18757),
            .in2(N__19297),
            .in3(N__16535),
            .lcout(\delay_measurement_inst.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__21973),
            .ce(N__18868),
            .sr(N__22295));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_26_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_26_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_26_5  (
            .in0(_gnd_net_),
            .in1(N__19315),
            .in2(N__19273),
            .in3(N__16511),
            .lcout(\delay_measurement_inst.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__21973),
            .ce(N__18868),
            .sr(N__22295));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_26_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_26_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_26_6  (
            .in0(_gnd_net_),
            .in1(N__19250),
            .in2(N__19298),
            .in3(N__16475),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__21973),
            .ce(N__18868),
            .sr(N__22295));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_26_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_26_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_26_7  (
            .in0(_gnd_net_),
            .in1(N__19226),
            .in2(N__19274),
            .in3(N__16454),
            .lcout(\delay_measurement_inst.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__21973),
            .ce(N__18868),
            .sr(N__22295));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_27_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_27_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_27_0  (
            .in0(_gnd_net_),
            .in1(N__19249),
            .in2(N__19201),
            .in3(N__16430),
            .lcout(\delay_measurement_inst.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_8_27_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__21971),
            .ce(N__18867),
            .sr(N__22299));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_27_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_27_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_27_1  (
            .in0(_gnd_net_),
            .in1(N__19225),
            .in2(N__19177),
            .in3(N__16403),
            .lcout(\delay_measurement_inst.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__21971),
            .ce(N__18867),
            .sr(N__22299));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_27_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_27_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_27_2  (
            .in0(_gnd_net_),
            .in1(N__19152),
            .in2(N__19202),
            .in3(N__16373),
            .lcout(\delay_measurement_inst.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__21971),
            .ce(N__18867),
            .sr(N__22299));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_27_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_27_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_27_3  (
            .in0(_gnd_net_),
            .in1(N__19134),
            .in2(N__19178),
            .in3(N__16802),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__21971),
            .ce(N__18867),
            .sr(N__22299));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_27_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_27_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_27_4  (
            .in0(_gnd_net_),
            .in1(N__19153),
            .in2(N__19495),
            .in3(N__16754),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__21971),
            .ce(N__18867),
            .sr(N__22299));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_27_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_27_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_27_5  (
            .in0(_gnd_net_),
            .in1(N__19135),
            .in2(N__19471),
            .in3(N__16724),
            .lcout(\delay_measurement_inst.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__21971),
            .ce(N__18867),
            .sr(N__22299));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_27_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_27_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_27_6  (
            .in0(_gnd_net_),
            .in1(N__19448),
            .in2(N__19496),
            .in3(N__16697),
            .lcout(\delay_measurement_inst.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__21971),
            .ce(N__18867),
            .sr(N__22299));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_27_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_27_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_27_7  (
            .in0(_gnd_net_),
            .in1(N__19424),
            .in2(N__19472),
            .in3(N__16670),
            .lcout(\delay_measurement_inst.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__21971),
            .ce(N__18867),
            .sr(N__22299));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_28_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_28_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_28_0  (
            .in0(_gnd_net_),
            .in1(N__19447),
            .in2(N__19399),
            .in3(N__16640),
            .lcout(\delay_measurement_inst.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_8_28_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__21967),
            .ce(N__18866),
            .sr(N__22302));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_28_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_28_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_28_1  (
            .in0(_gnd_net_),
            .in1(N__19423),
            .in2(N__19375),
            .in3(N__16622),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__21967),
            .ce(N__18866),
            .sr(N__22302));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_28_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_28_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_28_2  (
            .in0(_gnd_net_),
            .in1(N__19350),
            .in2(N__19400),
            .in3(N__16610),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__21967),
            .ce(N__18866),
            .sr(N__22302));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_28_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_28_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_28_3  (
            .in0(_gnd_net_),
            .in1(N__19332),
            .in2(N__19376),
            .in3(N__16907),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__21967),
            .ce(N__18866),
            .sr(N__22302));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_28_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_28_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_28_4  (
            .in0(_gnd_net_),
            .in1(N__19351),
            .in2(N__19684),
            .in3(N__16898),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__21967),
            .ce(N__18866),
            .sr(N__22302));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_28_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_28_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_28_5  (
            .in0(_gnd_net_),
            .in1(N__19333),
            .in2(N__19660),
            .in3(N__16889),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__21967),
            .ce(N__18866),
            .sr(N__22302));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_28_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_28_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_28_6  (
            .in0(_gnd_net_),
            .in1(N__19637),
            .in2(N__19685),
            .in3(N__16880),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__21967),
            .ce(N__18866),
            .sr(N__22302));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_28_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_28_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_28_7  (
            .in0(_gnd_net_),
            .in1(N__19613),
            .in2(N__19661),
            .in3(N__16868),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__21967),
            .ce(N__18866),
            .sr(N__22302));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_29_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_29_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_29_0  (
            .in0(_gnd_net_),
            .in1(N__19636),
            .in2(N__19588),
            .in3(N__16859),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_8_29_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__21963),
            .ce(N__18865),
            .sr(N__22304));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_29_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_29_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_29_1  (
            .in0(_gnd_net_),
            .in1(N__19612),
            .in2(N__19564),
            .in3(N__16850),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__21963),
            .ce(N__18865),
            .sr(N__22304));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_29_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_29_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_29_2  (
            .in0(_gnd_net_),
            .in1(N__19540),
            .in2(N__19589),
            .in3(N__16841),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__21963),
            .ce(N__18865),
            .sr(N__22304));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_29_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_29_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_29_3  (
            .in0(_gnd_net_),
            .in1(N__19522),
            .in2(N__19565),
            .in3(N__17102),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__21963),
            .ce(N__18865),
            .sr(N__22304));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_29_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_29_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_29_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_29_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17099),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21963),
            .ce(N__18865),
            .sr(N__22304));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_9_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_9_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__17072),
            .in2(N__17051),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_9_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_9_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__17036),
            .in2(_gnd_net_),
            .in3(N__17018),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_9_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_9_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__17015),
            .in2(N__17003),
            .in3(N__16985),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_9_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_9_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__16982),
            .in2(_gnd_net_),
            .in3(N__16964),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_9_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_9_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__16961),
            .in2(_gnd_net_),
            .in3(N__16943),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_9_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_9_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__16940),
            .in2(_gnd_net_),
            .in3(N__16922),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_9_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_9_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__17291),
            .in2(_gnd_net_),
            .in3(N__17273),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_9_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_9_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__17270),
            .in2(_gnd_net_),
            .in3(N__17252),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_9_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_9_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__17249),
            .in2(_gnd_net_),
            .in3(N__17231),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_9_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_9_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__17228),
            .in2(_gnd_net_),
            .in3(N__17207),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_9_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_9_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__17204),
            .in2(_gnd_net_),
            .in3(N__17186),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_9_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_9_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__17179),
            .in2(_gnd_net_),
            .in3(N__17159),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_9_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_9_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__17156),
            .in2(_gnd_net_),
            .in3(N__17135),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_9_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_9_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__17132),
            .in2(_gnd_net_),
            .in3(N__17114),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_9_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_9_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__17669),
            .in2(_gnd_net_),
            .in3(N__17648),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_9_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_9_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__17645),
            .in2(_gnd_net_),
            .in3(N__17627),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_9_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_9_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__17624),
            .in2(_gnd_net_),
            .in3(N__17606),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_9_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_9_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__17603),
            .in2(_gnd_net_),
            .in3(N__17585),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_9_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_9_15_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__17582),
            .in2(_gnd_net_),
            .in3(N__17570),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_9_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_9_16_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_0_LC_9_16_6  (
            .in0(N__17507),
            .in1(N__17398),
            .in2(N__20812),
            .in3(N__19714),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22005),
            .ce(N__21342),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__18422),
            .in2(N__17327),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_9_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_9_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(N__17312),
            .in2(_gnd_net_),
            .in3(N__17294),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_9_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_9_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(N__17867),
            .in2(N__17855),
            .in3(N__17831),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_9_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_9_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__17828),
            .in2(_gnd_net_),
            .in3(N__17810),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_9_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_9_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(N__17807),
            .in2(_gnd_net_),
            .in3(N__17789),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_9_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_9_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__17786),
            .in2(_gnd_net_),
            .in3(N__17768),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_9_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_9_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(N__17765),
            .in2(_gnd_net_),
            .in3(N__17747),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_9_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_9_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(N__17744),
            .in2(_gnd_net_),
            .in3(N__17714),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_9_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_9_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__17711),
            .in2(_gnd_net_),
            .in3(N__17693),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_9_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_9_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__17690),
            .in2(_gnd_net_),
            .in3(N__17672),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_9_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_9_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__18032),
            .in2(_gnd_net_),
            .in3(N__18014),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_9_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_9_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__18011),
            .in2(_gnd_net_),
            .in3(N__17993),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_9_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_9_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__17990),
            .in2(_gnd_net_),
            .in3(N__17972),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_9_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_9_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__17969),
            .in2(_gnd_net_),
            .in3(N__17951),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_9_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_9_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__17948),
            .in2(_gnd_net_),
            .in3(N__17930),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_9_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_9_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__17926),
            .in2(_gnd_net_),
            .in3(N__17906),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_9_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_9_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__17903),
            .in2(_gnd_net_),
            .in3(N__17882),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_9_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_9_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__17879),
            .in2(_gnd_net_),
            .in3(N__18524),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_9_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_9_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__18521),
            .in2(_gnd_net_),
            .in3(N__18509),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_9_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_9_19_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_9_19_5  (
            .in0(N__18215),
            .in1(N__20523),
            .in2(_gnd_net_),
            .in3(N__18347),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_20_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_20_2  (
            .in0(N__18446),
            .in1(N__18418),
            .in2(_gnd_net_),
            .in3(N__18398),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_9_20_4 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_9_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_1_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__20285),
            .in2(_gnd_net_),
            .in3(N__20365),
            .lcout(\phase_controller_slave.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_9_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_9_20_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_9_20_5  (
            .in0(N__20545),
            .in1(N__18321),
            .in2(_gnd_net_),
            .in3(N__18216),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_9_20_6 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_9_20_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_0_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__21222),
            .in2(_gnd_net_),
            .in3(N__21203),
            .lcout(\phase_controller_slave.N_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.S1_LC_9_21_3 .C_ON=1'b0;
    defparam \phase_controller_slave.S1_LC_9_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S1_LC_9_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.S1_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20288),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21984),
            .ce(),
            .sr(N__22265));
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_9_21_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_9_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_9_21_6 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_LC_9_21_6  (
            .in0(N__21205),
            .in1(N__18110),
            .in2(N__18077),
            .in3(N__18062),
            .lcout(\phase_controller_slave.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21984),
            .ce(),
            .sr(N__22265));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_5_LC_9_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_5_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_5_LC_9_23_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_14_5_LC_9_23_2  (
            .in0(N__18622),
            .in1(N__18634),
            .in2(N__18674),
            .in3(N__18544),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_4_LC_9_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_4_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_14_4_LC_9_23_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_14_4_LC_9_23_4  (
            .in0(N__18646),
            .in1(N__18658),
            .in2(N__18929),
            .in3(N__18556),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_9_24_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_9_24_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_9_24_0 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_30_LC_9_24_0  (
            .in0(N__18609),
            .in1(_gnd_net_),
            .in2(N__19117),
            .in3(N__18673),
            .lcout(measured_delay_hc_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21976),
            .ce(),
            .sr(N__22283));
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_9_24_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_9_24_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_9_24_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_24_LC_9_24_1  (
            .in0(N__18659),
            .in1(N__19073),
            .in2(_gnd_net_),
            .in3(N__18985),
            .lcout(measured_delay_hc_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21976),
            .ce(),
            .sr(N__22283));
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_9_24_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_9_24_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_9_24_2 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_25_LC_9_24_2  (
            .in0(N__18986),
            .in1(_gnd_net_),
            .in2(N__19114),
            .in3(N__18647),
            .lcout(measured_delay_hc_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21976),
            .ce(),
            .sr(N__22283));
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_9_24_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_9_24_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_9_24_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_28_LC_9_24_3  (
            .in0(N__18635),
            .in1(N__19081),
            .in2(_gnd_net_),
            .in3(N__18989),
            .lcout(measured_delay_hc_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21976),
            .ce(),
            .sr(N__22283));
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_9_24_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_9_24_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_9_24_4 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_29_LC_9_24_4  (
            .in0(N__18608),
            .in1(_gnd_net_),
            .in2(N__19116),
            .in3(N__18623),
            .lcout(measured_delay_hc_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21976),
            .ce(),
            .sr(N__22283));
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_9_24_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_9_24_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_9_24_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_23_LC_9_24_5  (
            .in0(N__18557),
            .in1(N__18607),
            .in2(_gnd_net_),
            .in3(N__19072),
            .lcout(measured_delay_hc_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21976),
            .ce(),
            .sr(N__22283));
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_9_24_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_9_24_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_9_24_6 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_27_LC_9_24_6  (
            .in0(N__18988),
            .in1(_gnd_net_),
            .in2(N__19115),
            .in3(N__18545),
            .lcout(measured_delay_hc_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21976),
            .ce(),
            .sr(N__22283));
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_9_24_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_9_24_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_9_24_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_26_LC_9_24_7  (
            .in0(N__18928),
            .in1(N__19077),
            .in2(_gnd_net_),
            .in3(N__18987),
            .lcout(measured_delay_hc_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21976),
            .ce(),
            .sr(N__22283));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_25_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_25_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18848),
            .lcout(\delay_measurement_inst.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21974),
            .ce(N__18869),
            .sr(N__22287));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_25_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_25_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_25_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_25_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18827),
            .lcout(\delay_measurement_inst.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21974),
            .ce(N__18869),
            .sr(N__22287));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_26_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_26_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_26_0  (
            .in0(N__21034),
            .in1(N__18846),
            .in2(_gnd_net_),
            .in3(N__18830),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_26_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__21972),
            .ce(N__21596),
            .sr(N__22292));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_26_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_26_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_26_1  (
            .in0(N__21059),
            .in1(N__18825),
            .in2(_gnd_net_),
            .in3(N__18809),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__21972),
            .ce(N__21596),
            .sr(N__22292));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_26_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_26_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_26_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_26_2  (
            .in0(N__21035),
            .in1(N__18804),
            .in2(_gnd_net_),
            .in3(N__18785),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__21972),
            .ce(N__21596),
            .sr(N__22292));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_26_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_26_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_26_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_26_3  (
            .in0(N__21060),
            .in1(N__18780),
            .in2(_gnd_net_),
            .in3(N__18761),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__21972),
            .ce(N__21596),
            .sr(N__22292));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_26_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_26_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_26_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_26_4  (
            .in0(N__21036),
            .in1(N__18758),
            .in2(_gnd_net_),
            .in3(N__18743),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__21972),
            .ce(N__21596),
            .sr(N__22292));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_26_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_26_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_26_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_26_5  (
            .in0(N__21061),
            .in1(N__19316),
            .in2(_gnd_net_),
            .in3(N__19301),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__21972),
            .ce(N__21596),
            .sr(N__22292));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_26_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_26_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_26_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_26_6  (
            .in0(N__21037),
            .in1(N__19296),
            .in2(_gnd_net_),
            .in3(N__19277),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__21972),
            .ce(N__21596),
            .sr(N__22292));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_26_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_26_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_26_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_26_7  (
            .in0(N__21062),
            .in1(N__19272),
            .in2(_gnd_net_),
            .in3(N__19253),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__21972),
            .ce(N__21596),
            .sr(N__22292));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_27_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_27_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_27_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_27_0  (
            .in0(N__21041),
            .in1(N__19248),
            .in2(_gnd_net_),
            .in3(N__19229),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_27_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__21968),
            .ce(N__21606),
            .sr(N__22296));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_27_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_27_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_27_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_27_1  (
            .in0(N__21045),
            .in1(N__19224),
            .in2(_gnd_net_),
            .in3(N__19205),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__21968),
            .ce(N__21606),
            .sr(N__22296));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_27_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_27_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_27_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_27_2  (
            .in0(N__21038),
            .in1(N__19200),
            .in2(_gnd_net_),
            .in3(N__19181),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__21968),
            .ce(N__21606),
            .sr(N__22296));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_27_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_27_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_27_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_27_3  (
            .in0(N__21042),
            .in1(N__19176),
            .in2(_gnd_net_),
            .in3(N__19157),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__21968),
            .ce(N__21606),
            .sr(N__22296));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_27_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_27_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_27_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_27_4  (
            .in0(N__21039),
            .in1(N__19154),
            .in2(_gnd_net_),
            .in3(N__19139),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__21968),
            .ce(N__21606),
            .sr(N__22296));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_27_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_27_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_27_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_27_5  (
            .in0(N__21043),
            .in1(N__19136),
            .in2(_gnd_net_),
            .in3(N__19121),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__21968),
            .ce(N__21606),
            .sr(N__22296));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_27_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_27_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_27_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_27_6  (
            .in0(N__21040),
            .in1(N__19494),
            .in2(_gnd_net_),
            .in3(N__19475),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__21968),
            .ce(N__21606),
            .sr(N__22296));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_27_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_27_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_27_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_27_7  (
            .in0(N__21044),
            .in1(N__19470),
            .in2(_gnd_net_),
            .in3(N__19451),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__21968),
            .ce(N__21606),
            .sr(N__22296));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_28_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_28_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_28_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_28_0  (
            .in0(N__21072),
            .in1(N__19446),
            .in2(_gnd_net_),
            .in3(N__19427),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_9_28_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__21964),
            .ce(N__21607),
            .sr(N__22300));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_28_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_28_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_28_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_28_1  (
            .in0(N__21055),
            .in1(N__19422),
            .in2(_gnd_net_),
            .in3(N__19403),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__21964),
            .ce(N__21607),
            .sr(N__22300));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_28_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_28_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_28_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_28_2  (
            .in0(N__21073),
            .in1(N__19398),
            .in2(_gnd_net_),
            .in3(N__19379),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__21964),
            .ce(N__21607),
            .sr(N__22300));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_28_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_28_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_28_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_28_3  (
            .in0(N__21056),
            .in1(N__19374),
            .in2(_gnd_net_),
            .in3(N__19355),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__21964),
            .ce(N__21607),
            .sr(N__22300));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_28_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_28_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_28_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_28_4  (
            .in0(N__21074),
            .in1(N__19352),
            .in2(_gnd_net_),
            .in3(N__19337),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__21964),
            .ce(N__21607),
            .sr(N__22300));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_28_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_28_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_28_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_28_5  (
            .in0(N__21057),
            .in1(N__19334),
            .in2(_gnd_net_),
            .in3(N__19319),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__21964),
            .ce(N__21607),
            .sr(N__22300));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_28_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_28_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_28_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_28_6  (
            .in0(N__21075),
            .in1(N__19683),
            .in2(_gnd_net_),
            .in3(N__19664),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__21964),
            .ce(N__21607),
            .sr(N__22300));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_28_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_28_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_28_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_28_7  (
            .in0(N__21058),
            .in1(N__19659),
            .in2(_gnd_net_),
            .in3(N__19640),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__21964),
            .ce(N__21607),
            .sr(N__22300));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_29_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_29_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_29_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_29_0  (
            .in0(N__21063),
            .in1(N__19635),
            .in2(_gnd_net_),
            .in3(N__19616),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_9_29_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__21961),
            .ce(N__21608),
            .sr(N__22303));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_29_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_29_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_29_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_29_1  (
            .in0(N__21076),
            .in1(N__19611),
            .in2(_gnd_net_),
            .in3(N__19592),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__21961),
            .ce(N__21608),
            .sr(N__22303));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_29_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_29_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_29_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_29_2  (
            .in0(N__21064),
            .in1(N__19587),
            .in2(_gnd_net_),
            .in3(N__19568),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__21961),
            .ce(N__21608),
            .sr(N__22303));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_29_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_29_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_29_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_29_3  (
            .in0(N__21077),
            .in1(N__19563),
            .in2(_gnd_net_),
            .in3(N__19544),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__21961),
            .ce(N__21608),
            .sr(N__22303));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_29_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_29_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_29_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_29_4  (
            .in0(N__21065),
            .in1(N__19541),
            .in2(_gnd_net_),
            .in3(N__19529),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__21961),
            .ce(N__21608),
            .sr(N__22303));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_29_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_29_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_29_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_29_5  (
            .in0(N__19523),
            .in1(N__21066),
            .in2(_gnd_net_),
            .in3(N__19526),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21961),
            .ce(N__21608),
            .sr(N__22303));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_10_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_10_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(N__21513),
            .in2(_gnd_net_),
            .in3(N__21479),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_138_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_10_12_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_10_12_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_10_12_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_10_12_5 (
            .in0(N__20186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22017),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_13_3.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_13_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_10_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20168),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22011),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_10_14_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_10_14_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_10_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_10_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20162),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22007),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_14_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_14_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_10_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20144),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22007),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_10_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_10_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_10_15_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__20138),
            .in2(_gnd_net_),
            .in3(N__20033),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21999),
            .ce(N__19945),
            .sr(N__22232));
    defparam \phase_controller_inst1.state_0_LC_10_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_10_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_10_16_0 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \phase_controller_inst1.state_0_LC_10_16_0  (
            .in0(N__21181),
            .in1(N__20249),
            .in2(N__20267),
            .in3(N__20209),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21994),
            .ce(),
            .sr(N__22235));
    defparam \phase_controller_slave.start_timer_tr_LC_10_16_1 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_LC_10_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_tr_LC_10_16_1 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \phase_controller_slave.start_timer_tr_LC_10_16_1  (
            .in0(N__19788),
            .in1(N__20237),
            .in2(N__20344),
            .in3(N__20216),
            .lcout(\phase_controller_slave.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21994),
            .ce(),
            .sr(N__22235));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_10_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_10_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_10_16_6 .LUT_INIT=16'b1010100010111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_10_16_6  (
            .in0(N__20266),
            .in1(N__19751),
            .in2(N__19742),
            .in3(N__19718),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21994),
            .ce(),
            .sr(N__22235));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_10_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_10_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__20262),
            .in2(_gnd_net_),
            .in3(N__20248),
            .lcout(\phase_controller_inst1.N_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_RNIR0JF_1_LC_10_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNIR0JF_1_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNIR0JF_1_LC_10_17_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.state_RNIR0JF_1_LC_10_17_2  (
            .in0(N__21170),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20208),
            .lcout(\phase_controller_inst1.T01_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_tr_RNO_1_LC_10_17_3 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_RNO_1_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_tr_RNO_1_LC_10_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_tr_RNO_1_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__21125),
            .in2(_gnd_net_),
            .in3(N__21240),
            .lcout(\phase_controller_slave.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_10_17_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_10_17_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_10_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_10_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20231),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21991),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_17_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__21548),
            .in2(_gnd_net_),
            .in3(N__20679),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_10_17_7 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_10_17_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_tr_RNO_0_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(N__20496),
            .in2(_gnd_net_),
            .in3(N__20463),
            .lcout(\phase_controller_slave.N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_1_LC_10_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_10_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_10_18_0 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_inst1.state_1_LC_10_18_0  (
            .in0(N__20438),
            .in1(N__20417),
            .in2(N__21180),
            .in3(N__20210),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21987),
            .ce(),
            .sr(N__22240));
    defparam \phase_controller_slave.state_0_LC_10_18_1 .C_ON=1'b0;
    defparam \phase_controller_slave.state_0_LC_10_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_0_LC_10_18_1 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_slave.state_0_LC_10_18_1  (
            .in0(N__21248),
            .in1(N__20497),
            .in2(N__21131),
            .in3(N__20464),
            .lcout(\phase_controller_slave.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21987),
            .ce(),
            .sr(N__22240));
    defparam \phase_controller_inst1.state_2_LC_10_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_10_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_10_18_2 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst1.state_2_LC_10_18_2  (
            .in0(N__20681),
            .in1(N__20436),
            .in2(N__21556),
            .in3(N__20416),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21987),
            .ce(),
            .sr(N__22240));
    defparam \phase_controller_inst1.T01_LC_10_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_LC_10_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T01_LC_10_18_3 .LUT_INIT=16'b1010101010101110;
    LogicCell40 \phase_controller_inst1.T01_LC_10_18_3  (
            .in0(N__20437),
            .in1(N__20450),
            .in2(N__21644),
            .in3(N__20854),
            .lcout(shift_flag_start),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21987),
            .ce(),
            .sr(N__22240));
    defparam \phase_controller_inst1.start_timer_tr_LC_10_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_10_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_10_18_4 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_10_18_4  (
            .in0(N__20855),
            .in1(N__21643),
            .in2(N__20778),
            .in3(N__20689),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21987),
            .ce(),
            .sr(N__22240));
    defparam \phase_controller_inst1.state_3_LC_10_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_10_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_10_18_5 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \phase_controller_inst1.state_3_LC_10_18_5  (
            .in0(N__20690),
            .in1(N__21552),
            .in2(N__21617),
            .in3(N__20680),
            .lcout(\phase_controller_inst1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21987),
            .ce(),
            .sr(N__22240));
    defparam \phase_controller_inst1.start_timer_hc_LC_10_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_10_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_10_18_6 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_10_18_6  (
            .in0(N__20663),
            .in1(N__21642),
            .in2(N__20594),
            .in3(N__20381),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21987),
            .ce(),
            .sr(N__22240));
    defparam \phase_controller_slave.state_4_LC_10_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.state_4_LC_10_18_7 .SEQ_MODE=4'b1011;
    defparam \phase_controller_slave.state_4_LC_10_18_7 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_slave.state_4_LC_10_18_7  (
            .in0(N__20299),
            .in1(N__20498),
            .in2(N__20333),
            .in3(N__20465),
            .lcout(\phase_controller_slave.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21987),
            .ce(),
            .sr(N__22240));
    defparam \phase_controller_slave.un1_start_LC_10_19_2 .C_ON=1'b0;
    defparam \phase_controller_slave.un1_start_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.un1_start_LC_10_19_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.un1_start_LC_10_19_2  (
            .in0(N__21709),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20449),
            .lcout(\phase_controller_slave.un1_startZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_10_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_10_19_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__20435),
            .in2(_gnd_net_),
            .in3(N__20410),
            .lcout(\phase_controller_inst1.N_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.state_2_LC_10_20_1 .C_ON=1'b0;
    defparam \phase_controller_slave.state_2_LC_10_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_2_LC_10_20_1 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_slave.state_2_LC_10_20_1  (
            .in0(N__20375),
            .in1(N__20287),
            .in2(N__21227),
            .in3(N__21204),
            .lcout(\phase_controller_slave.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21981),
            .ce(),
            .sr(N__22247));
    defparam \phase_controller_slave.state_3_LC_10_20_2 .C_ON=1'b0;
    defparam \phase_controller_slave.state_3_LC_10_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_3_LC_10_20_2 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \phase_controller_slave.state_3_LC_10_20_2  (
            .in0(N__20286),
            .in1(N__20374),
            .in2(N__20343),
            .in3(N__20300),
            .lcout(\phase_controller_slave.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21981),
            .ce(),
            .sr(N__22247));
    defparam \phase_controller_slave.state_1_LC_10_21_2 .C_ON=1'b0;
    defparam \phase_controller_slave.state_1_LC_10_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_1_LC_10_21_2 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_slave.state_1_LC_10_21_2  (
            .in0(N__21247),
            .in1(N__21226),
            .in2(N__21126),
            .in3(N__21206),
            .lcout(\phase_controller_slave.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21978),
            .ce(),
            .sr(N__22252));
    defparam \phase_controller_inst1.S2_LC_10_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_10_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_10_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21182),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21977),
            .ce(),
            .sr(N__22259));
    defparam \phase_controller_slave.S2_LC_10_25_5 .C_ON=1'b0;
    defparam \phase_controller_slave.S2_LC_10_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S2_LC_10_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.S2_LC_10_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21130),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21969),
            .ce(),
            .sr(N__22277));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_10_26_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_10_26_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_10_26_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_10_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21761),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_11_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_11_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_11_12_2 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_11_12_2  (
            .in0(N__21515),
            .in1(N__21497),
            .in2(_gnd_net_),
            .in3(N__21484),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22012),
            .ce(),
            .sr(N__22231));
    defparam \delay_measurement_inst.stop_timer_tr_LC_11_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_tr_LC_11_12_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_11_12_4  (
            .in0(N__21394),
            .in1(N__21419),
            .in2(_gnd_net_),
            .in3(N__21374),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22012),
            .ce(),
            .sr(N__22231));
    defparam \delay_measurement_inst.start_timer_tr_LC_11_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_tr_LC_11_12_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_11_12_5  (
            .in0(N__21418),
            .in1(N__21373),
            .in2(_gnd_net_),
            .in3(N__21393),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22012),
            .ce(),
            .sr(N__22231));
    defparam \delay_measurement_inst.prev_tr_sig_LC_11_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_tr_sig_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_tr_sig_LC_11_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.prev_tr_sig_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21420),
            .lcout(\delay_measurement_inst.prev_tr_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22012),
            .ce(),
            .sr(N__22231));
    defparam \delay_measurement_inst.tr_state_RNIFBI31_0_LC_11_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_RNIFBI31_0_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.tr_state_RNIFBI31_0_LC_11_13_0 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \delay_measurement_inst.tr_state_RNIFBI31_0_LC_11_13_0  (
            .in0(N__21371),
            .in1(N__21392),
            .in2(N__21422),
            .in3(N__20951),
            .lcout(\delay_measurement_inst.un1_tr_state_1_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_4_LC_11_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_11_17_3 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_11_17_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__21707),
            .in2(_gnd_net_),
            .in3(N__21638),
            .lcout(\phase_controller_inst1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21988),
            .ce(),
            .sr(N__22236));
    defparam \phase_controller_inst1.state_RNO_0_3_LC_11_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_11_18_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.state_RNO_0_3_LC_11_18_1  (
            .in0(N__21708),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21637),
            .lcout(\phase_controller_inst1.N_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_26_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_26_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_26_7 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_26_7  (
            .in0(N__22414),
            .in1(N__21785),
            .in2(_gnd_net_),
            .in3(N__21759),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_137_i_g ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S1_LC_11_28_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_11_28_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_11_28_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_11_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21563),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21959),
            .ce(),
            .sr(N__22288));
    defparam SB_DFF_inst_DELAY_TR2_LC_12_12_0.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR2_LC_12_12_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR2_LC_12_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR2_LC_12_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21428),
            .lcout(delay_tr_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22006),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_12_3 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_12_3  (
            .in0(N__21514),
            .in1(N__21496),
            .in2(_gnd_net_),
            .in3(N__21480),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_139_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR1_LC_12_12_5.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR1_LC_12_12_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR1_LC_12_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR1_LC_12_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21446),
            .lcout(delay_tr_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22006),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_state_0_LC_12_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_0_LC_12_13_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.tr_state_0_LC_12_13_2 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.tr_state_0_LC_12_13_2  (
            .in0(N__21421),
            .in1(N__21372),
            .in2(_gnd_net_),
            .in3(N__21395),
            .lcout(\delay_measurement_inst.tr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21998),
            .ce(N__21349),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.hc_state_0_LC_12_24_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_state_0_LC_12_24_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.hc_state_0_LC_12_24_1 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.hc_state_0_LC_12_24_1  (
            .in0(N__22377),
            .in1(N__22359),
            .in2(_gnd_net_),
            .in3(N__22071),
            .lcout(\delay_measurement_inst.hc_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21965),
            .ce(N__21338),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_12_25_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_12_25_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_hc_LC_12_25_4 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_12_25_4  (
            .in0(N__22379),
            .in1(N__22360),
            .in2(_gnd_net_),
            .in3(N__22076),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21962),
            .ce(),
            .sr(N__22269));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_26_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_26_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_26_4 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_12_26_4  (
            .in0(N__22415),
            .in1(N__21781),
            .in2(_gnd_net_),
            .in3(N__21760),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21960),
            .ce(),
            .sr(N__22274));
    defparam SB_DFF_inst_DELAY_HC1_LC_13_17_3.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC1_LC_13_17_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC1_LC_13_17_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_DELAY_HC1_LC_13_17_3 (
            .in0(N__22403),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(delay_hc_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21989),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC2_LC_13_22_0.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC2_LC_13_22_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC2_LC_13_22_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC2_LC_13_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22388),
            .lcout(delay_hc_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21975),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.prev_hc_sig_LC_13_24_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_hc_sig_LC_13_24_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_hc_sig_LC_13_24_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.prev_hc_sig_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(N__22075),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.prev_hc_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21970),
            .ce(),
            .sr(N__22253));
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_25_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_25_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_25_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_13_25_1  (
            .in0(N__22378),
            .in1(N__22361),
            .in2(N__22343),
            .in3(N__22070),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21966),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_26_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_26_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(N__21777),
            .in2(_gnd_net_),
            .in3(N__21755),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_136_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // MAIN
