-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Feb 27 2025 18:59:42

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    rgb_g : out std_logic;
    T01 : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    T23 : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    clock_output : out std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    T45 : out std_logic;
    T12 : out std_logic;
    s4_phy : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__49535\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49514\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49487\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49479\ : std_logic;
signal \N__49478\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49452\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49433\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49415\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49406\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49398\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49396\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49388\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49379\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49361\ : std_logic;
signal \N__49358\ : std_logic;
signal \N__49355\ : std_logic;
signal \N__49352\ : std_logic;
signal \N__49349\ : std_logic;
signal \N__49346\ : std_logic;
signal \N__49345\ : std_logic;
signal \N__49342\ : std_logic;
signal \N__49339\ : std_logic;
signal \N__49336\ : std_logic;
signal \N__49331\ : std_logic;
signal \N__49330\ : std_logic;
signal \N__49329\ : std_logic;
signal \N__49322\ : std_logic;
signal \N__49319\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49316\ : std_logic;
signal \N__49313\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49301\ : std_logic;
signal \N__49300\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49294\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49285\ : std_logic;
signal \N__49282\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49276\ : std_logic;
signal \N__49273\ : std_logic;
signal \N__49268\ : std_logic;
signal \N__49265\ : std_logic;
signal \N__49262\ : std_logic;
signal \N__49259\ : std_logic;
signal \N__49256\ : std_logic;
signal \N__49253\ : std_logic;
signal \N__49252\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49246\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49238\ : std_logic;
signal \N__49235\ : std_logic;
signal \N__49234\ : std_logic;
signal \N__49233\ : std_logic;
signal \N__49230\ : std_logic;
signal \N__49225\ : std_logic;
signal \N__49222\ : std_logic;
signal \N__49219\ : std_logic;
signal \N__49214\ : std_logic;
signal \N__49211\ : std_logic;
signal \N__49208\ : std_logic;
signal \N__49207\ : std_logic;
signal \N__49204\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49192\ : std_logic;
signal \N__49187\ : std_logic;
signal \N__49184\ : std_logic;
signal \N__49181\ : std_logic;
signal \N__49178\ : std_logic;
signal \N__49177\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49168\ : std_logic;
signal \N__49163\ : std_logic;
signal \N__49160\ : std_logic;
signal \N__49159\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49145\ : std_logic;
signal \N__49142\ : std_logic;
signal \N__49139\ : std_logic;
signal \N__49136\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49127\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49097\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49067\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49065\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49062\ : std_logic;
signal \N__49059\ : std_logic;
signal \N__49056\ : std_logic;
signal \N__49055\ : std_logic;
signal \N__49054\ : std_logic;
signal \N__49051\ : std_logic;
signal \N__49050\ : std_logic;
signal \N__49045\ : std_logic;
signal \N__49042\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49036\ : std_logic;
signal \N__49031\ : std_logic;
signal \N__49026\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49010\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49001\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48995\ : std_logic;
signal \N__48990\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48980\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48978\ : std_logic;
signal \N__48977\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48963\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48960\ : std_logic;
signal \N__48959\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48953\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48947\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48930\ : std_logic;
signal \N__48927\ : std_logic;
signal \N__48924\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48908\ : std_logic;
signal \N__48907\ : std_logic;
signal \N__48904\ : std_logic;
signal \N__48901\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48897\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48883\ : std_logic;
signal \N__48878\ : std_logic;
signal \N__48875\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48868\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48859\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48846\ : std_logic;
signal \N__48843\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48827\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48809\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48807\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48804\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48796\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48794\ : std_logic;
signal \N__48793\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48791\ : std_logic;
signal \N__48790\ : std_logic;
signal \N__48789\ : std_logic;
signal \N__48788\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48785\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48783\ : std_logic;
signal \N__48782\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48780\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48777\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48772\ : std_logic;
signal \N__48771\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48762\ : std_logic;
signal \N__48761\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48758\ : std_logic;
signal \N__48757\ : std_logic;
signal \N__48756\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48752\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48750\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48747\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48744\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48741\ : std_logic;
signal \N__48740\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48738\ : std_logic;
signal \N__48737\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48732\ : std_logic;
signal \N__48731\ : std_logic;
signal \N__48730\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48727\ : std_logic;
signal \N__48726\ : std_logic;
signal \N__48725\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48712\ : std_logic;
signal \N__48711\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48707\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48704\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48698\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48695\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48693\ : std_logic;
signal \N__48692\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48690\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48687\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48684\ : std_logic;
signal \N__48683\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48679\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48677\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48675\ : std_logic;
signal \N__48674\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48672\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48669\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48665\ : std_logic;
signal \N__48664\ : std_logic;
signal \N__48663\ : std_logic;
signal \N__48662\ : std_logic;
signal \N__48661\ : std_logic;
signal \N__48660\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48658\ : std_logic;
signal \N__48657\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48650\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48311\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48309\ : std_logic;
signal \N__48308\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48302\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48290\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48282\ : std_logic;
signal \N__48281\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48277\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48274\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48271\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48268\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48255\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48252\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48249\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48246\ : std_logic;
signal \N__48245\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48240\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48230\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48224\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48219\ : std_logic;
signal \N__48218\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48212\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48209\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48204\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48200\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48184\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48178\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48175\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48172\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48145\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48142\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48136\ : std_logic;
signal \N__48135\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48127\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48124\ : std_logic;
signal \N__48123\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47773\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47740\ : std_logic;
signal \N__47737\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47718\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47710\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47639\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47614\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47571\ : std_logic;
signal \N__47568\ : std_logic;
signal \N__47565\ : std_logic;
signal \N__47562\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47553\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47539\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47532\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47504\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47471\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47389\ : std_logic;
signal \N__47386\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47266\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47254\ : std_logic;
signal \N__47251\ : std_logic;
signal \N__47248\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47223\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47186\ : std_logic;
signal \N__47183\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47161\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47148\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47145\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47142\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47139\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47132\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47130\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47114\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47111\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47108\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47091\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47083\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47065\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47059\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47026\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46949\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46715\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46685\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46682\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46679\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46675\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46615\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46592\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46454\ : std_logic;
signal \N__46451\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46436\ : std_logic;
signal \N__46427\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46400\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46368\ : std_logic;
signal \N__46365\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46337\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46316\ : std_logic;
signal \N__46313\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46247\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46130\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46115\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46109\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45938\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45901\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45895\ : std_logic;
signal \N__45892\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45858\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45847\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45829\ : std_logic;
signal \N__45826\ : std_logic;
signal \N__45823\ : std_logic;
signal \N__45820\ : std_logic;
signal \N__45817\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45811\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45746\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45710\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45700\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45469\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45431\ : std_logic;
signal \N__45428\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45421\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45395\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45368\ : std_logic;
signal \N__45365\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45356\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45332\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45320\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45308\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45272\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45259\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45230\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45199\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45179\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45164\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45125\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45023\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45008\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44996\ : std_logic;
signal \N__44993\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44942\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44855\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44837\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44826\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44810\ : std_logic;
signal \N__44809\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44767\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44747\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44690\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44686\ : std_logic;
signal \N__44683\ : std_logic;
signal \N__44680\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44672\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44651\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44534\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44516\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44467\ : std_logic;
signal \N__44464\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44452\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44391\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44211\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44147\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44113\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44033\ : std_logic;
signal \N__44030\ : std_logic;
signal \N__44027\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44017\ : std_logic;
signal \N__44016\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43999\ : std_logic;
signal \N__43996\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43989\ : std_logic;
signal \N__43986\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43975\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43961\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43935\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43925\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43883\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43877\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43868\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43802\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43788\ : std_logic;
signal \N__43785\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43741\ : std_logic;
signal \N__43738\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43706\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43631\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43618\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43498\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43418\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43383\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43374\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43272\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43204\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43181\ : std_logic;
signal \N__43178\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43155\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43067\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43061\ : std_logic;
signal \N__43058\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42868\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42854\ : std_logic;
signal \N__42851\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42802\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42748\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42700\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42668\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42569\ : std_logic;
signal \N__42566\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42557\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42553\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42533\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42389\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42355\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42349\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42344\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42210\ : std_logic;
signal \N__42207\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42142\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42101\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41980\ : std_logic;
signal \N__41977\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41948\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41942\ : std_logic;
signal \N__41939\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41933\ : std_logic;
signal \N__41930\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41924\ : std_logic;
signal \N__41921\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41906\ : std_logic;
signal \N__41903\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41897\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41890\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41849\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41783\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41776\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41762\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41687\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41659\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41415\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41403\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41386\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41273\ : std_logic;
signal \N__41270\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41225\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41195\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41173\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41165\ : std_logic;
signal \N__41162\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41051\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41032\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40972\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40870\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40709\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40688\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40662\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40649\ : std_logic;
signal \N__40646\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40560\ : std_logic;
signal \N__40557\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40424\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40128\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40074\ : std_logic;
signal \N__40071\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40055\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39986\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39959\ : std_logic;
signal \N__39956\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39935\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39911\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39329\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39069\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38997\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38605\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38354\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38240\ : std_logic;
signal \N__38237\ : std_logic;
signal \N__38234\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38225\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38063\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37729\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36189\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\ : std_logic;
signal \rgb_drv_RNOZ0\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator\ : std_logic;
signal \bfn_3_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \bfn_3_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_17\ : std_logic;
signal \bfn_3_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_25\ : std_logic;
signal \bfn_3_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \N_38_i_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_77_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_7_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_7_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_7_23_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_8_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_8_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal s4_phy_c : std_logic;
signal \GB_BUFFER_clock_output_0_THRU_CO\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30\ : std_logic;
signal \current_shift_inst.control_input_18\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \elapsed_time_ns_1_RNIE03T9_0_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \elapsed_time_ns_1_RNIF13T9_0_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \elapsed_time_ns_1_RNIV2EN9_0_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \elapsed_time_ns_1_RNI04EN9_0_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \elapsed_time_ns_1_RNIDV2T9_0_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df30_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \current_shift_inst.control_input_axb_0_cascade_\ : std_logic;
signal \current_shift_inst.N_1288_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \bfn_10_20_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt18\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_11_23_0_\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_11_24_0_\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal s3_phy_c : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_12_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.state_RNIG7JFZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_start_g\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_199_i\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_198_i\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\ : std_logic;
signal \bfn_12_21_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_12_22_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_15\ : std_logic;
signal \pwm_generator_inst.threshold_3\ : std_logic;
signal \pwm_generator_inst.threshold_4\ : std_logic;
signal \pwm_generator_inst.threshold_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_1\ : std_logic;
signal \pwm_generator_inst.threshold_0\ : std_logic;
signal \pwm_generator_inst.threshold_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_8\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.threshold_9\ : std_logic;
signal \pll_inst.red_c_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\ : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.N_162_i_g\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.timer_s1.N_162_i\ : std_logic;
signal \current_shift_inst.timer_s1.N_163_i\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\ : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\ : std_logic;
signal \bfn_13_25_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_8\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_15\ : std_logic;
signal \bfn_13_28_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_23\ : std_logic;
signal \bfn_13_29_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_13_30_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_16\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal state_ns_i_a3_1 : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_0\ : std_logic;
signal \bfn_14_25_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_8\ : std_logic;
signal \bfn_14_26_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_14_27_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold\ : std_logic;
signal \bfn_14_28_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_axbZ0Z_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\ : std_logic;
signal \bfn_14_29_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\ : std_logic;
signal \bfn_14_30_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal s1_phy_c : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal state_3 : std_logic;
signal \T01_c\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \bfn_15_24_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \bfn_15_25_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \bfn_15_26_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\ : std_logic;
signal \phase_controller_inst1.state_RNIE87FZ0Z_2\ : std_logic;
signal \T45_c\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \T23_c\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal start_stop_c : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNIDC91B_0_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \elapsed_time_ns_1_RNIED91B_0_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \elapsed_time_ns_1_RNIFE91B_0_3\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_200_i\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_201_i\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \T12_c\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.state_RNI7NN7Z0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_10\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_18_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_18_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt18\ : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt30\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_start_g\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\ : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal pwm_duty_input_7 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal pwm_duty_input_8 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal pwm_duty_input_1 : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_159\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal \_gnd_net_\ : std_logic;
signal clock_output_0 : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal clock_output_wire : std_logic;
signal \T01_wire\ : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal \T23_wire\ : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal \T12_wire\ : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal \T45_wire\ : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    clock_output <= clock_output_wire;
    T01 <= \T01_wire\;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    T23 <= \T23_wire\;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    T12 <= \T12_wire\;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    T45 <= \T45_wire\;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ <= \N__26826\&\N__26834\&\N__26825\&\N__26832\&\N__26824\&\N__26831\&\N__26823\&\N__26833\&\N__26820\&\N__26827\&\N__26819\&\N__26828\&\N__26822\&\N__26829\&\N__26821\&\N__26830\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__37883\&'0'&\N__37882\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__30965\&\N__30958\&\N__30963\&\N__30957\&\N__30964\&\N__30956\&\N__30966\&\N__30953\&\N__30959\&\N__30952\&\N__30960\&\N__30954\&\N__30961\&\N__30955\&\N__30962\;
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__37790\&\N__37787\&'0'&'0'&'0'&\N__37785\&\N__37789\&\N__37786\&\N__37788\;
    \pwm_generator_inst.un2_threshold_2_1_16\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_2_1_15\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_2_14\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_2_13\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_2_12\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_2_11\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_2_10\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_2_9\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_2_8\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_2_7\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_2_6\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_2_5\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_2_4\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_2_3\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_2_2\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_2_1\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_2_0\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ <= '0'&\N__30967\&\N__30970\&\N__30968\&\N__30971\&\N__30969\&\N__48825\&\N__47666\&\N__47726\&\N__49207\&\N__49158\&\N__49083\&\N__47571\&\N__49256\&\N__49346\&\N__47636\;
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__37891\&\N__37888\&'0'&'0'&'0'&\N__37886\&\N__37890\&\N__37887\&\N__37889\;
    \pwm_generator_inst.un2_threshold_1_25\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_1_24\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_1_23\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_1_22\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_1_21\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_1_20\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_1_19\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_1_18\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_1_17\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_1_16\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_1_15\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(0);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ <= '0'&\N__26780\&\N__22846\&\N__20309\&\N__22921\&\N__22867\&\N__36830\&\N__33898\&\N__39389\&\N__33931\&\N__36931\&\N__36901\&\N__36316\&\N__22804\&\N__22900\&\N__47269\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__37797\&'0'&\N__37796\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(19);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(18);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(17);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(16);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.un1_integrator\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__20075\,
            RESETB => \N__30797\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clock_output_0
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__37884\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__37881\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__37791\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__37784\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__37909\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__37885\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__37798\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__37795\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__49533\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49535\,
            DIN => \N__49534\,
            DOUT => \N__49533\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49535\,
            PADOUT => \N__49534\,
            PADIN => \N__49533\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clock_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49524\,
            DIN => \N__49523\,
            DOUT => \N__49522\,
            PACKAGEPIN => clock_output_wire
        );

    \clock_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49524\,
            PADOUT => \N__49523\,
            PADIN => \N__49522\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21884\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T01_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49515\,
            DIN => \N__49514\,
            DOUT => \N__49513\,
            PACKAGEPIN => \T01_wire\
        );

    \T01_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49515\,
            PADOUT => \N__49514\,
            PADIN => \N__49513\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__39272\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49506\,
            DIN => \N__49505\,
            DOUT => \N__49504\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49506\,
            PADOUT => \N__49505\,
            PADIN => \N__49504\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49497\,
            DIN => \N__49496\,
            DOUT => \N__49495\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49497\,
            PADOUT => \N__49496\,
            PADIN => \N__49495\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T23_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49488\,
            DIN => \N__49487\,
            DOUT => \N__49486\,
            PACKAGEPIN => \T23_wire\
        );

    \T23_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49488\,
            PADOUT => \N__49487\,
            PADIN => \N__49486\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__42593\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49479\,
            DIN => \N__49478\,
            DOUT => \N__49477\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49479\,
            PADOUT => \N__49478\,
            PADIN => \N__49477\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__27389\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49470\,
            DIN => \N__49469\,
            DOUT => \N__49468\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49470\,
            PADOUT => \N__49469\,
            PADIN => \N__49468\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49461\,
            DIN => \N__49460\,
            DOUT => \N__49459\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49461\,
            PADOUT => \N__49460\,
            PADIN => \N__49459\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__43037\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T12_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49452\,
            DIN => \N__49451\,
            DOUT => \N__49450\,
            PACKAGEPIN => \T12_wire\
        );

    \T12_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49452\,
            PADOUT => \N__49451\,
            PADIN => \N__49450\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__44603\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49443\,
            DIN => \N__49442\,
            DOUT => \N__49441\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49443\,
            PADOUT => \N__49442\,
            PADIN => \N__49441\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49434\,
            DIN => \N__49433\,
            DOUT => \N__49432\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49434\,
            PADOUT => \N__49433\,
            PADIN => \N__49432\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__39362\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49425\,
            DIN => \N__49424\,
            DOUT => \N__49423\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49425\,
            PADOUT => \N__49424\,
            PADIN => \N__49423\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21893\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49416\,
            DIN => \N__49415\,
            DOUT => \N__49414\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49416\,
            PADOUT => \N__49415\,
            PADIN => \N__49414\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49407\,
            DIN => \N__49406\,
            DOUT => \N__49405\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49407\,
            PADOUT => \N__49406\,
            PADIN => \N__49405\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__27365\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T45_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49398\,
            DIN => \N__49397\,
            DOUT => \N__49396\,
            PACKAGEPIN => \T45_wire\
        );

    \T45_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49398\,
            PADOUT => \N__49397\,
            PADIN => \N__49396\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__42656\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49389\,
            DIN => \N__49388\,
            DOUT => \N__49387\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49389\,
            PADOUT => \N__49388\,
            PADIN => \N__49387\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49380\,
            DIN => \N__49379\,
            DOUT => \N__49378\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49380\,
            PADOUT => \N__49379\,
            PADIN => \N__49378\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11861\ : InMux
    port map (
            O => \N__49361\,
            I => \N__49358\
        );

    \I__11860\ : LocalMux
    port map (
            O => \N__49358\,
            I => \N__49355\
        );

    \I__11859\ : Span4Mux_h
    port map (
            O => \N__49355\,
            I => \N__49352\
        );

    \I__11858\ : Span4Mux_h
    port map (
            O => \N__49352\,
            I => \N__49349\
        );

    \I__11857\ : Odrv4
    port map (
            O => \N__49349\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__11856\ : InMux
    port map (
            O => \N__49346\,
            I => \N__49342\
        );

    \I__11855\ : InMux
    port map (
            O => \N__49345\,
            I => \N__49339\
        );

    \I__11854\ : LocalMux
    port map (
            O => \N__49342\,
            I => \N__49336\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__49339\,
            I => pwm_duty_input_1
        );

    \I__11852\ : Odrv4
    port map (
            O => \N__49336\,
            I => pwm_duty_input_1
        );

    \I__11851\ : InMux
    port map (
            O => \N__49331\,
            I => \N__49322\
        );

    \I__11850\ : InMux
    port map (
            O => \N__49330\,
            I => \N__49322\
        );

    \I__11849\ : InMux
    port map (
            O => \N__49329\,
            I => \N__49322\
        );

    \I__11848\ : LocalMux
    port map (
            O => \N__49322\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \I__11847\ : CascadeMux
    port map (
            O => \N__49319\,
            I => \N__49313\
        );

    \I__11846\ : InMux
    port map (
            O => \N__49318\,
            I => \N__49304\
        );

    \I__11845\ : InMux
    port map (
            O => \N__49317\,
            I => \N__49304\
        );

    \I__11844\ : InMux
    port map (
            O => \N__49316\,
            I => \N__49304\
        );

    \I__11843\ : InMux
    port map (
            O => \N__49313\,
            I => \N__49304\
        );

    \I__11842\ : LocalMux
    port map (
            O => \N__49304\,
            I => \N__49301\
        );

    \I__11841\ : Span4Mux_s3_h
    port map (
            O => \N__49301\,
            I => \N__49297\
        );

    \I__11840\ : InMux
    port map (
            O => \N__49300\,
            I => \N__49294\
        );

    \I__11839\ : Odrv4
    port map (
            O => \N__49297\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__11838\ : LocalMux
    port map (
            O => \N__49294\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__11837\ : CascadeMux
    port map (
            O => \N__49289\,
            I => \N__49285\
        );

    \I__11836\ : CascadeMux
    port map (
            O => \N__49288\,
            I => \N__49282\
        );

    \I__11835\ : InMux
    port map (
            O => \N__49285\,
            I => \N__49276\
        );

    \I__11834\ : InMux
    port map (
            O => \N__49282\,
            I => \N__49276\
        );

    \I__11833\ : InMux
    port map (
            O => \N__49281\,
            I => \N__49273\
        );

    \I__11832\ : LocalMux
    port map (
            O => \N__49276\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__11831\ : LocalMux
    port map (
            O => \N__49273\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__11830\ : InMux
    port map (
            O => \N__49268\,
            I => \N__49265\
        );

    \I__11829\ : LocalMux
    port map (
            O => \N__49265\,
            I => \N__49262\
        );

    \I__11828\ : Span12Mux_s3_h
    port map (
            O => \N__49262\,
            I => \N__49259\
        );

    \I__11827\ : Odrv12
    port map (
            O => \N__49259\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__11826\ : InMux
    port map (
            O => \N__49256\,
            I => \N__49253\
        );

    \I__11825\ : LocalMux
    port map (
            O => \N__49253\,
            I => \N__49249\
        );

    \I__11824\ : InMux
    port map (
            O => \N__49252\,
            I => \N__49246\
        );

    \I__11823\ : Span4Mux_s1_h
    port map (
            O => \N__49249\,
            I => \N__49243\
        );

    \I__11822\ : LocalMux
    port map (
            O => \N__49246\,
            I => pwm_duty_input_2
        );

    \I__11821\ : Odrv4
    port map (
            O => \N__49243\,
            I => pwm_duty_input_2
        );

    \I__11820\ : CascadeMux
    port map (
            O => \N__49238\,
            I => \N__49235\
        );

    \I__11819\ : InMux
    port map (
            O => \N__49235\,
            I => \N__49230\
        );

    \I__11818\ : InMux
    port map (
            O => \N__49234\,
            I => \N__49225\
        );

    \I__11817\ : InMux
    port map (
            O => \N__49233\,
            I => \N__49225\
        );

    \I__11816\ : LocalMux
    port map (
            O => \N__49230\,
            I => \N__49222\
        );

    \I__11815\ : LocalMux
    port map (
            O => \N__49225\,
            I => \N__49219\
        );

    \I__11814\ : Span4Mux_s2_h
    port map (
            O => \N__49222\,
            I => \N__49214\
        );

    \I__11813\ : Span4Mux_v
    port map (
            O => \N__49219\,
            I => \N__49214\
        );

    \I__11812\ : Span4Mux_h
    port map (
            O => \N__49214\,
            I => \N__49211\
        );

    \I__11811\ : Odrv4
    port map (
            O => \N__49211\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__11810\ : CascadeMux
    port map (
            O => \N__49208\,
            I => \N__49204\
        );

    \I__11809\ : InMux
    port map (
            O => \N__49207\,
            I => \N__49200\
        );

    \I__11808\ : InMux
    port map (
            O => \N__49204\,
            I => \N__49195\
        );

    \I__11807\ : InMux
    port map (
            O => \N__49203\,
            I => \N__49195\
        );

    \I__11806\ : LocalMux
    port map (
            O => \N__49200\,
            I => \N__49192\
        );

    \I__11805\ : LocalMux
    port map (
            O => \N__49195\,
            I => pwm_duty_input_6
        );

    \I__11804\ : Odrv4
    port map (
            O => \N__49192\,
            I => pwm_duty_input_6
        );

    \I__11803\ : CascadeMux
    port map (
            O => \N__49187\,
            I => \N__49184\
        );

    \I__11802\ : InMux
    port map (
            O => \N__49184\,
            I => \N__49181\
        );

    \I__11801\ : LocalMux
    port map (
            O => \N__49181\,
            I => \N__49178\
        );

    \I__11800\ : Span4Mux_v
    port map (
            O => \N__49178\,
            I => \N__49173\
        );

    \I__11799\ : InMux
    port map (
            O => \N__49177\,
            I => \N__49168\
        );

    \I__11798\ : InMux
    port map (
            O => \N__49176\,
            I => \N__49168\
        );

    \I__11797\ : Sp12to4
    port map (
            O => \N__49173\,
            I => \N__49163\
        );

    \I__11796\ : LocalMux
    port map (
            O => \N__49168\,
            I => \N__49163\
        );

    \I__11795\ : Odrv12
    port map (
            O => \N__49163\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__11794\ : InMux
    port map (
            O => \N__49160\,
            I => \N__49153\
        );

    \I__11793\ : InMux
    port map (
            O => \N__49159\,
            I => \N__49153\
        );

    \I__11792\ : InMux
    port map (
            O => \N__49158\,
            I => \N__49150\
        );

    \I__11791\ : LocalMux
    port map (
            O => \N__49153\,
            I => pwm_duty_input_5
        );

    \I__11790\ : LocalMux
    port map (
            O => \N__49150\,
            I => pwm_duty_input_5
        );

    \I__11789\ : InMux
    port map (
            O => \N__49145\,
            I => \N__49142\
        );

    \I__11788\ : LocalMux
    port map (
            O => \N__49142\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__11787\ : InMux
    port map (
            O => \N__49139\,
            I => \N__49136\
        );

    \I__11786\ : LocalMux
    port map (
            O => \N__49136\,
            I => \N__49133\
        );

    \I__11785\ : Odrv12
    port map (
            O => \N__49133\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__11784\ : CascadeMux
    port map (
            O => \N__49130\,
            I => \N__49127\
        );

    \I__11783\ : InMux
    port map (
            O => \N__49127\,
            I => \N__49122\
        );

    \I__11782\ : InMux
    port map (
            O => \N__49126\,
            I => \N__49117\
        );

    \I__11781\ : InMux
    port map (
            O => \N__49125\,
            I => \N__49117\
        );

    \I__11780\ : LocalMux
    port map (
            O => \N__49122\,
            I => \N__49111\
        );

    \I__11779\ : LocalMux
    port map (
            O => \N__49117\,
            I => \N__49111\
        );

    \I__11778\ : InMux
    port map (
            O => \N__49116\,
            I => \N__49108\
        );

    \I__11777\ : Span4Mux_s2_h
    port map (
            O => \N__49111\,
            I => \N__49103\
        );

    \I__11776\ : LocalMux
    port map (
            O => \N__49108\,
            I => \N__49103\
        );

    \I__11775\ : Span4Mux_h
    port map (
            O => \N__49103\,
            I => \N__49100\
        );

    \I__11774\ : Span4Mux_h
    port map (
            O => \N__49100\,
            I => \N__49097\
        );

    \I__11773\ : Odrv4
    port map (
            O => \N__49097\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__11772\ : CascadeMux
    port map (
            O => \N__49094\,
            I => \N__49091\
        );

    \I__11771\ : InMux
    port map (
            O => \N__49091\,
            I => \N__49088\
        );

    \I__11770\ : LocalMux
    port map (
            O => \N__49088\,
            I => \N__49084\
        );

    \I__11769\ : InMux
    port map (
            O => \N__49087\,
            I => \N__49080\
        );

    \I__11768\ : Span4Mux_h
    port map (
            O => \N__49084\,
            I => \N__49077\
        );

    \I__11767\ : InMux
    port map (
            O => \N__49083\,
            I => \N__49074\
        );

    \I__11766\ : LocalMux
    port map (
            O => \N__49080\,
            I => pwm_duty_input_4
        );

    \I__11765\ : Odrv4
    port map (
            O => \N__49077\,
            I => pwm_duty_input_4
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__49074\,
            I => pwm_duty_input_4
        );

    \I__11763\ : CascadeMux
    port map (
            O => \N__49067\,
            I => \N__49059\
        );

    \I__11762\ : CascadeMux
    port map (
            O => \N__49066\,
            I => \N__49056\
        );

    \I__11761\ : CascadeMux
    port map (
            O => \N__49065\,
            I => \N__49051\
        );

    \I__11760\ : InMux
    port map (
            O => \N__49064\,
            I => \N__49045\
        );

    \I__11759\ : InMux
    port map (
            O => \N__49063\,
            I => \N__49045\
        );

    \I__11758\ : InMux
    port map (
            O => \N__49062\,
            I => \N__49042\
        );

    \I__11757\ : InMux
    port map (
            O => \N__49059\,
            I => \N__49039\
        );

    \I__11756\ : InMux
    port map (
            O => \N__49056\,
            I => \N__49036\
        );

    \I__11755\ : InMux
    port map (
            O => \N__49055\,
            I => \N__49031\
        );

    \I__11754\ : InMux
    port map (
            O => \N__49054\,
            I => \N__49031\
        );

    \I__11753\ : InMux
    port map (
            O => \N__49051\,
            I => \N__49026\
        );

    \I__11752\ : InMux
    port map (
            O => \N__49050\,
            I => \N__49026\
        );

    \I__11751\ : LocalMux
    port map (
            O => \N__49045\,
            I => \N__49021\
        );

    \I__11750\ : LocalMux
    port map (
            O => \N__49042\,
            I => \N__49021\
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__49039\,
            I => \N__49018\
        );

    \I__11748\ : LocalMux
    port map (
            O => \N__49036\,
            I => \N__49015\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__49031\,
            I => \N__49010\
        );

    \I__11746\ : LocalMux
    port map (
            O => \N__49026\,
            I => \N__49010\
        );

    \I__11745\ : Span4Mux_v
    port map (
            O => \N__49021\,
            I => \N__49007\
        );

    \I__11744\ : Span4Mux_s3_h
    port map (
            O => \N__49018\,
            I => \N__49004\
        );

    \I__11743\ : Span4Mux_s3_h
    port map (
            O => \N__49015\,
            I => \N__49001\
        );

    \I__11742\ : Span4Mux_s3_h
    port map (
            O => \N__49010\,
            I => \N__48998\
        );

    \I__11741\ : Span4Mux_h
    port map (
            O => \N__49007\,
            I => \N__48995\
        );

    \I__11740\ : Span4Mux_h
    port map (
            O => \N__49004\,
            I => \N__48990\
        );

    \I__11739\ : Span4Mux_h
    port map (
            O => \N__49001\,
            I => \N__48990\
        );

    \I__11738\ : Span4Mux_h
    port map (
            O => \N__48998\,
            I => \N__48987\
        );

    \I__11737\ : Odrv4
    port map (
            O => \N__48995\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__11736\ : Odrv4
    port map (
            O => \N__48990\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__11735\ : Odrv4
    port map (
            O => \N__48987\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__11734\ : InMux
    port map (
            O => \N__48980\,
            I => \N__48973\
        );

    \I__11733\ : InMux
    port map (
            O => \N__48979\,
            I => \N__48968\
        );

    \I__11732\ : InMux
    port map (
            O => \N__48978\,
            I => \N__48968\
        );

    \I__11731\ : InMux
    port map (
            O => \N__48977\,
            I => \N__48963\
        );

    \I__11730\ : InMux
    port map (
            O => \N__48976\,
            I => \N__48963\
        );

    \I__11729\ : LocalMux
    port map (
            O => \N__48973\,
            I => \N__48953\
        );

    \I__11728\ : LocalMux
    port map (
            O => \N__48968\,
            I => \N__48953\
        );

    \I__11727\ : LocalMux
    port map (
            O => \N__48963\,
            I => \N__48950\
        );

    \I__11726\ : InMux
    port map (
            O => \N__48962\,
            I => \N__48947\
        );

    \I__11725\ : InMux
    port map (
            O => \N__48961\,
            I => \N__48940\
        );

    \I__11724\ : InMux
    port map (
            O => \N__48960\,
            I => \N__48940\
        );

    \I__11723\ : InMux
    port map (
            O => \N__48959\,
            I => \N__48940\
        );

    \I__11722\ : InMux
    port map (
            O => \N__48958\,
            I => \N__48937\
        );

    \I__11721\ : Span4Mux_v
    port map (
            O => \N__48953\,
            I => \N__48930\
        );

    \I__11720\ : Span4Mux_s1_h
    port map (
            O => \N__48950\,
            I => \N__48930\
        );

    \I__11719\ : LocalMux
    port map (
            O => \N__48947\,
            I => \N__48930\
        );

    \I__11718\ : LocalMux
    port map (
            O => \N__48940\,
            I => \N__48927\
        );

    \I__11717\ : LocalMux
    port map (
            O => \N__48937\,
            I => \N__48924\
        );

    \I__11716\ : Span4Mux_h
    port map (
            O => \N__48930\,
            I => \N__48919\
        );

    \I__11715\ : Span4Mux_h
    port map (
            O => \N__48927\,
            I => \N__48919\
        );

    \I__11714\ : Span4Mux_h
    port map (
            O => \N__48924\,
            I => \N__48916\
        );

    \I__11713\ : Span4Mux_h
    port map (
            O => \N__48919\,
            I => \N__48913\
        );

    \I__11712\ : Odrv4
    port map (
            O => \N__48916\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__11711\ : Odrv4
    port map (
            O => \N__48913\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__11710\ : CascadeMux
    port map (
            O => \N__48908\,
            I => \N__48904\
        );

    \I__11709\ : CascadeMux
    port map (
            O => \N__48907\,
            I => \N__48901\
        );

    \I__11708\ : InMux
    port map (
            O => \N__48904\,
            I => \N__48897\
        );

    \I__11707\ : InMux
    port map (
            O => \N__48901\,
            I => \N__48894\
        );

    \I__11706\ : InMux
    port map (
            O => \N__48900\,
            I => \N__48891\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__48897\,
            I => \N__48888\
        );

    \I__11704\ : LocalMux
    port map (
            O => \N__48894\,
            I => \N__48883\
        );

    \I__11703\ : LocalMux
    port map (
            O => \N__48891\,
            I => \N__48883\
        );

    \I__11702\ : Span4Mux_s3_h
    port map (
            O => \N__48888\,
            I => \N__48878\
        );

    \I__11701\ : Span4Mux_v
    port map (
            O => \N__48883\,
            I => \N__48878\
        );

    \I__11700\ : Span4Mux_h
    port map (
            O => \N__48878\,
            I => \N__48875\
        );

    \I__11699\ : Odrv4
    port map (
            O => \N__48875\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__11698\ : InMux
    port map (
            O => \N__48872\,
            I => \N__48864\
        );

    \I__11697\ : InMux
    port map (
            O => \N__48871\,
            I => \N__48859\
        );

    \I__11696\ : InMux
    port map (
            O => \N__48870\,
            I => \N__48859\
        );

    \I__11695\ : InMux
    port map (
            O => \N__48869\,
            I => \N__48852\
        );

    \I__11694\ : InMux
    port map (
            O => \N__48868\,
            I => \N__48852\
        );

    \I__11693\ : InMux
    port map (
            O => \N__48867\,
            I => \N__48852\
        );

    \I__11692\ : LocalMux
    port map (
            O => \N__48864\,
            I => \N__48846\
        );

    \I__11691\ : LocalMux
    port map (
            O => \N__48859\,
            I => \N__48846\
        );

    \I__11690\ : LocalMux
    port map (
            O => \N__48852\,
            I => \N__48843\
        );

    \I__11689\ : InMux
    port map (
            O => \N__48851\,
            I => \N__48840\
        );

    \I__11688\ : Span4Mux_v
    port map (
            O => \N__48846\,
            I => \N__48833\
        );

    \I__11687\ : Span4Mux_s1_h
    port map (
            O => \N__48843\,
            I => \N__48833\
        );

    \I__11686\ : LocalMux
    port map (
            O => \N__48840\,
            I => \N__48833\
        );

    \I__11685\ : Span4Mux_h
    port map (
            O => \N__48833\,
            I => \N__48830\
        );

    \I__11684\ : Odrv4
    port map (
            O => \N__48830\,
            I => \current_shift_inst.PI_CTRL.N_159\
        );

    \I__11683\ : InMux
    port map (
            O => \N__48827\,
            I => \N__48820\
        );

    \I__11682\ : InMux
    port map (
            O => \N__48826\,
            I => \N__48820\
        );

    \I__11681\ : InMux
    port map (
            O => \N__48825\,
            I => \N__48817\
        );

    \I__11680\ : LocalMux
    port map (
            O => \N__48820\,
            I => pwm_duty_input_9
        );

    \I__11679\ : LocalMux
    port map (
            O => \N__48817\,
            I => pwm_duty_input_9
        );

    \I__11678\ : InMux
    port map (
            O => \N__48812\,
            I => \N__48809\
        );

    \I__11677\ : LocalMux
    port map (
            O => \N__48809\,
            I => \N__48643\
        );

    \I__11676\ : ClkMux
    port map (
            O => \N__48808\,
            I => \N__48314\
        );

    \I__11675\ : ClkMux
    port map (
            O => \N__48807\,
            I => \N__48314\
        );

    \I__11674\ : ClkMux
    port map (
            O => \N__48806\,
            I => \N__48314\
        );

    \I__11673\ : ClkMux
    port map (
            O => \N__48805\,
            I => \N__48314\
        );

    \I__11672\ : ClkMux
    port map (
            O => \N__48804\,
            I => \N__48314\
        );

    \I__11671\ : ClkMux
    port map (
            O => \N__48803\,
            I => \N__48314\
        );

    \I__11670\ : ClkMux
    port map (
            O => \N__48802\,
            I => \N__48314\
        );

    \I__11669\ : ClkMux
    port map (
            O => \N__48801\,
            I => \N__48314\
        );

    \I__11668\ : ClkMux
    port map (
            O => \N__48800\,
            I => \N__48314\
        );

    \I__11667\ : ClkMux
    port map (
            O => \N__48799\,
            I => \N__48314\
        );

    \I__11666\ : ClkMux
    port map (
            O => \N__48798\,
            I => \N__48314\
        );

    \I__11665\ : ClkMux
    port map (
            O => \N__48797\,
            I => \N__48314\
        );

    \I__11664\ : ClkMux
    port map (
            O => \N__48796\,
            I => \N__48314\
        );

    \I__11663\ : ClkMux
    port map (
            O => \N__48795\,
            I => \N__48314\
        );

    \I__11662\ : ClkMux
    port map (
            O => \N__48794\,
            I => \N__48314\
        );

    \I__11661\ : ClkMux
    port map (
            O => \N__48793\,
            I => \N__48314\
        );

    \I__11660\ : ClkMux
    port map (
            O => \N__48792\,
            I => \N__48314\
        );

    \I__11659\ : ClkMux
    port map (
            O => \N__48791\,
            I => \N__48314\
        );

    \I__11658\ : ClkMux
    port map (
            O => \N__48790\,
            I => \N__48314\
        );

    \I__11657\ : ClkMux
    port map (
            O => \N__48789\,
            I => \N__48314\
        );

    \I__11656\ : ClkMux
    port map (
            O => \N__48788\,
            I => \N__48314\
        );

    \I__11655\ : ClkMux
    port map (
            O => \N__48787\,
            I => \N__48314\
        );

    \I__11654\ : ClkMux
    port map (
            O => \N__48786\,
            I => \N__48314\
        );

    \I__11653\ : ClkMux
    port map (
            O => \N__48785\,
            I => \N__48314\
        );

    \I__11652\ : ClkMux
    port map (
            O => \N__48784\,
            I => \N__48314\
        );

    \I__11651\ : ClkMux
    port map (
            O => \N__48783\,
            I => \N__48314\
        );

    \I__11650\ : ClkMux
    port map (
            O => \N__48782\,
            I => \N__48314\
        );

    \I__11649\ : ClkMux
    port map (
            O => \N__48781\,
            I => \N__48314\
        );

    \I__11648\ : ClkMux
    port map (
            O => \N__48780\,
            I => \N__48314\
        );

    \I__11647\ : ClkMux
    port map (
            O => \N__48779\,
            I => \N__48314\
        );

    \I__11646\ : ClkMux
    port map (
            O => \N__48778\,
            I => \N__48314\
        );

    \I__11645\ : ClkMux
    port map (
            O => \N__48777\,
            I => \N__48314\
        );

    \I__11644\ : ClkMux
    port map (
            O => \N__48776\,
            I => \N__48314\
        );

    \I__11643\ : ClkMux
    port map (
            O => \N__48775\,
            I => \N__48314\
        );

    \I__11642\ : ClkMux
    port map (
            O => \N__48774\,
            I => \N__48314\
        );

    \I__11641\ : ClkMux
    port map (
            O => \N__48773\,
            I => \N__48314\
        );

    \I__11640\ : ClkMux
    port map (
            O => \N__48772\,
            I => \N__48314\
        );

    \I__11639\ : ClkMux
    port map (
            O => \N__48771\,
            I => \N__48314\
        );

    \I__11638\ : ClkMux
    port map (
            O => \N__48770\,
            I => \N__48314\
        );

    \I__11637\ : ClkMux
    port map (
            O => \N__48769\,
            I => \N__48314\
        );

    \I__11636\ : ClkMux
    port map (
            O => \N__48768\,
            I => \N__48314\
        );

    \I__11635\ : ClkMux
    port map (
            O => \N__48767\,
            I => \N__48314\
        );

    \I__11634\ : ClkMux
    port map (
            O => \N__48766\,
            I => \N__48314\
        );

    \I__11633\ : ClkMux
    port map (
            O => \N__48765\,
            I => \N__48314\
        );

    \I__11632\ : ClkMux
    port map (
            O => \N__48764\,
            I => \N__48314\
        );

    \I__11631\ : ClkMux
    port map (
            O => \N__48763\,
            I => \N__48314\
        );

    \I__11630\ : ClkMux
    port map (
            O => \N__48762\,
            I => \N__48314\
        );

    \I__11629\ : ClkMux
    port map (
            O => \N__48761\,
            I => \N__48314\
        );

    \I__11628\ : ClkMux
    port map (
            O => \N__48760\,
            I => \N__48314\
        );

    \I__11627\ : ClkMux
    port map (
            O => \N__48759\,
            I => \N__48314\
        );

    \I__11626\ : ClkMux
    port map (
            O => \N__48758\,
            I => \N__48314\
        );

    \I__11625\ : ClkMux
    port map (
            O => \N__48757\,
            I => \N__48314\
        );

    \I__11624\ : ClkMux
    port map (
            O => \N__48756\,
            I => \N__48314\
        );

    \I__11623\ : ClkMux
    port map (
            O => \N__48755\,
            I => \N__48314\
        );

    \I__11622\ : ClkMux
    port map (
            O => \N__48754\,
            I => \N__48314\
        );

    \I__11621\ : ClkMux
    port map (
            O => \N__48753\,
            I => \N__48314\
        );

    \I__11620\ : ClkMux
    port map (
            O => \N__48752\,
            I => \N__48314\
        );

    \I__11619\ : ClkMux
    port map (
            O => \N__48751\,
            I => \N__48314\
        );

    \I__11618\ : ClkMux
    port map (
            O => \N__48750\,
            I => \N__48314\
        );

    \I__11617\ : ClkMux
    port map (
            O => \N__48749\,
            I => \N__48314\
        );

    \I__11616\ : ClkMux
    port map (
            O => \N__48748\,
            I => \N__48314\
        );

    \I__11615\ : ClkMux
    port map (
            O => \N__48747\,
            I => \N__48314\
        );

    \I__11614\ : ClkMux
    port map (
            O => \N__48746\,
            I => \N__48314\
        );

    \I__11613\ : ClkMux
    port map (
            O => \N__48745\,
            I => \N__48314\
        );

    \I__11612\ : ClkMux
    port map (
            O => \N__48744\,
            I => \N__48314\
        );

    \I__11611\ : ClkMux
    port map (
            O => \N__48743\,
            I => \N__48314\
        );

    \I__11610\ : ClkMux
    port map (
            O => \N__48742\,
            I => \N__48314\
        );

    \I__11609\ : ClkMux
    port map (
            O => \N__48741\,
            I => \N__48314\
        );

    \I__11608\ : ClkMux
    port map (
            O => \N__48740\,
            I => \N__48314\
        );

    \I__11607\ : ClkMux
    port map (
            O => \N__48739\,
            I => \N__48314\
        );

    \I__11606\ : ClkMux
    port map (
            O => \N__48738\,
            I => \N__48314\
        );

    \I__11605\ : ClkMux
    port map (
            O => \N__48737\,
            I => \N__48314\
        );

    \I__11604\ : ClkMux
    port map (
            O => \N__48736\,
            I => \N__48314\
        );

    \I__11603\ : ClkMux
    port map (
            O => \N__48735\,
            I => \N__48314\
        );

    \I__11602\ : ClkMux
    port map (
            O => \N__48734\,
            I => \N__48314\
        );

    \I__11601\ : ClkMux
    port map (
            O => \N__48733\,
            I => \N__48314\
        );

    \I__11600\ : ClkMux
    port map (
            O => \N__48732\,
            I => \N__48314\
        );

    \I__11599\ : ClkMux
    port map (
            O => \N__48731\,
            I => \N__48314\
        );

    \I__11598\ : ClkMux
    port map (
            O => \N__48730\,
            I => \N__48314\
        );

    \I__11597\ : ClkMux
    port map (
            O => \N__48729\,
            I => \N__48314\
        );

    \I__11596\ : ClkMux
    port map (
            O => \N__48728\,
            I => \N__48314\
        );

    \I__11595\ : ClkMux
    port map (
            O => \N__48727\,
            I => \N__48314\
        );

    \I__11594\ : ClkMux
    port map (
            O => \N__48726\,
            I => \N__48314\
        );

    \I__11593\ : ClkMux
    port map (
            O => \N__48725\,
            I => \N__48314\
        );

    \I__11592\ : ClkMux
    port map (
            O => \N__48724\,
            I => \N__48314\
        );

    \I__11591\ : ClkMux
    port map (
            O => \N__48723\,
            I => \N__48314\
        );

    \I__11590\ : ClkMux
    port map (
            O => \N__48722\,
            I => \N__48314\
        );

    \I__11589\ : ClkMux
    port map (
            O => \N__48721\,
            I => \N__48314\
        );

    \I__11588\ : ClkMux
    port map (
            O => \N__48720\,
            I => \N__48314\
        );

    \I__11587\ : ClkMux
    port map (
            O => \N__48719\,
            I => \N__48314\
        );

    \I__11586\ : ClkMux
    port map (
            O => \N__48718\,
            I => \N__48314\
        );

    \I__11585\ : ClkMux
    port map (
            O => \N__48717\,
            I => \N__48314\
        );

    \I__11584\ : ClkMux
    port map (
            O => \N__48716\,
            I => \N__48314\
        );

    \I__11583\ : ClkMux
    port map (
            O => \N__48715\,
            I => \N__48314\
        );

    \I__11582\ : ClkMux
    port map (
            O => \N__48714\,
            I => \N__48314\
        );

    \I__11581\ : ClkMux
    port map (
            O => \N__48713\,
            I => \N__48314\
        );

    \I__11580\ : ClkMux
    port map (
            O => \N__48712\,
            I => \N__48314\
        );

    \I__11579\ : ClkMux
    port map (
            O => \N__48711\,
            I => \N__48314\
        );

    \I__11578\ : ClkMux
    port map (
            O => \N__48710\,
            I => \N__48314\
        );

    \I__11577\ : ClkMux
    port map (
            O => \N__48709\,
            I => \N__48314\
        );

    \I__11576\ : ClkMux
    port map (
            O => \N__48708\,
            I => \N__48314\
        );

    \I__11575\ : ClkMux
    port map (
            O => \N__48707\,
            I => \N__48314\
        );

    \I__11574\ : ClkMux
    port map (
            O => \N__48706\,
            I => \N__48314\
        );

    \I__11573\ : ClkMux
    port map (
            O => \N__48705\,
            I => \N__48314\
        );

    \I__11572\ : ClkMux
    port map (
            O => \N__48704\,
            I => \N__48314\
        );

    \I__11571\ : ClkMux
    port map (
            O => \N__48703\,
            I => \N__48314\
        );

    \I__11570\ : ClkMux
    port map (
            O => \N__48702\,
            I => \N__48314\
        );

    \I__11569\ : ClkMux
    port map (
            O => \N__48701\,
            I => \N__48314\
        );

    \I__11568\ : ClkMux
    port map (
            O => \N__48700\,
            I => \N__48314\
        );

    \I__11567\ : ClkMux
    port map (
            O => \N__48699\,
            I => \N__48314\
        );

    \I__11566\ : ClkMux
    port map (
            O => \N__48698\,
            I => \N__48314\
        );

    \I__11565\ : ClkMux
    port map (
            O => \N__48697\,
            I => \N__48314\
        );

    \I__11564\ : ClkMux
    port map (
            O => \N__48696\,
            I => \N__48314\
        );

    \I__11563\ : ClkMux
    port map (
            O => \N__48695\,
            I => \N__48314\
        );

    \I__11562\ : ClkMux
    port map (
            O => \N__48694\,
            I => \N__48314\
        );

    \I__11561\ : ClkMux
    port map (
            O => \N__48693\,
            I => \N__48314\
        );

    \I__11560\ : ClkMux
    port map (
            O => \N__48692\,
            I => \N__48314\
        );

    \I__11559\ : ClkMux
    port map (
            O => \N__48691\,
            I => \N__48314\
        );

    \I__11558\ : ClkMux
    port map (
            O => \N__48690\,
            I => \N__48314\
        );

    \I__11557\ : ClkMux
    port map (
            O => \N__48689\,
            I => \N__48314\
        );

    \I__11556\ : ClkMux
    port map (
            O => \N__48688\,
            I => \N__48314\
        );

    \I__11555\ : ClkMux
    port map (
            O => \N__48687\,
            I => \N__48314\
        );

    \I__11554\ : ClkMux
    port map (
            O => \N__48686\,
            I => \N__48314\
        );

    \I__11553\ : ClkMux
    port map (
            O => \N__48685\,
            I => \N__48314\
        );

    \I__11552\ : ClkMux
    port map (
            O => \N__48684\,
            I => \N__48314\
        );

    \I__11551\ : ClkMux
    port map (
            O => \N__48683\,
            I => \N__48314\
        );

    \I__11550\ : ClkMux
    port map (
            O => \N__48682\,
            I => \N__48314\
        );

    \I__11549\ : ClkMux
    port map (
            O => \N__48681\,
            I => \N__48314\
        );

    \I__11548\ : ClkMux
    port map (
            O => \N__48680\,
            I => \N__48314\
        );

    \I__11547\ : ClkMux
    port map (
            O => \N__48679\,
            I => \N__48314\
        );

    \I__11546\ : ClkMux
    port map (
            O => \N__48678\,
            I => \N__48314\
        );

    \I__11545\ : ClkMux
    port map (
            O => \N__48677\,
            I => \N__48314\
        );

    \I__11544\ : ClkMux
    port map (
            O => \N__48676\,
            I => \N__48314\
        );

    \I__11543\ : ClkMux
    port map (
            O => \N__48675\,
            I => \N__48314\
        );

    \I__11542\ : ClkMux
    port map (
            O => \N__48674\,
            I => \N__48314\
        );

    \I__11541\ : ClkMux
    port map (
            O => \N__48673\,
            I => \N__48314\
        );

    \I__11540\ : ClkMux
    port map (
            O => \N__48672\,
            I => \N__48314\
        );

    \I__11539\ : ClkMux
    port map (
            O => \N__48671\,
            I => \N__48314\
        );

    \I__11538\ : ClkMux
    port map (
            O => \N__48670\,
            I => \N__48314\
        );

    \I__11537\ : ClkMux
    port map (
            O => \N__48669\,
            I => \N__48314\
        );

    \I__11536\ : ClkMux
    port map (
            O => \N__48668\,
            I => \N__48314\
        );

    \I__11535\ : ClkMux
    port map (
            O => \N__48667\,
            I => \N__48314\
        );

    \I__11534\ : ClkMux
    port map (
            O => \N__48666\,
            I => \N__48314\
        );

    \I__11533\ : ClkMux
    port map (
            O => \N__48665\,
            I => \N__48314\
        );

    \I__11532\ : ClkMux
    port map (
            O => \N__48664\,
            I => \N__48314\
        );

    \I__11531\ : ClkMux
    port map (
            O => \N__48663\,
            I => \N__48314\
        );

    \I__11530\ : ClkMux
    port map (
            O => \N__48662\,
            I => \N__48314\
        );

    \I__11529\ : ClkMux
    port map (
            O => \N__48661\,
            I => \N__48314\
        );

    \I__11528\ : ClkMux
    port map (
            O => \N__48660\,
            I => \N__48314\
        );

    \I__11527\ : ClkMux
    port map (
            O => \N__48659\,
            I => \N__48314\
        );

    \I__11526\ : ClkMux
    port map (
            O => \N__48658\,
            I => \N__48314\
        );

    \I__11525\ : ClkMux
    port map (
            O => \N__48657\,
            I => \N__48314\
        );

    \I__11524\ : ClkMux
    port map (
            O => \N__48656\,
            I => \N__48314\
        );

    \I__11523\ : ClkMux
    port map (
            O => \N__48655\,
            I => \N__48314\
        );

    \I__11522\ : ClkMux
    port map (
            O => \N__48654\,
            I => \N__48314\
        );

    \I__11521\ : ClkMux
    port map (
            O => \N__48653\,
            I => \N__48314\
        );

    \I__11520\ : ClkMux
    port map (
            O => \N__48652\,
            I => \N__48314\
        );

    \I__11519\ : ClkMux
    port map (
            O => \N__48651\,
            I => \N__48314\
        );

    \I__11518\ : ClkMux
    port map (
            O => \N__48650\,
            I => \N__48314\
        );

    \I__11517\ : ClkMux
    port map (
            O => \N__48649\,
            I => \N__48314\
        );

    \I__11516\ : ClkMux
    port map (
            O => \N__48648\,
            I => \N__48314\
        );

    \I__11515\ : ClkMux
    port map (
            O => \N__48647\,
            I => \N__48314\
        );

    \I__11514\ : ClkMux
    port map (
            O => \N__48646\,
            I => \N__48314\
        );

    \I__11513\ : Glb2LocalMux
    port map (
            O => \N__48643\,
            I => \N__48314\
        );

    \I__11512\ : GlobalMux
    port map (
            O => \N__48314\,
            I => clock_output_0
        );

    \I__11511\ : InMux
    port map (
            O => \N__48311\,
            I => \N__48305\
        );

    \I__11510\ : InMux
    port map (
            O => \N__48310\,
            I => \N__48302\
        );

    \I__11509\ : InMux
    port map (
            O => \N__48309\,
            I => \N__48299\
        );

    \I__11508\ : InMux
    port map (
            O => \N__48308\,
            I => \N__48296\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__48305\,
            I => \N__48293\
        );

    \I__11506\ : LocalMux
    port map (
            O => \N__48302\,
            I => \N__48290\
        );

    \I__11505\ : LocalMux
    port map (
            O => \N__48299\,
            I => \N__48287\
        );

    \I__11504\ : LocalMux
    port map (
            O => \N__48296\,
            I => \N__48283\
        );

    \I__11503\ : Glb2LocalMux
    port map (
            O => \N__48293\,
            I => \N__47786\
        );

    \I__11502\ : Glb2LocalMux
    port map (
            O => \N__48290\,
            I => \N__47786\
        );

    \I__11501\ : Glb2LocalMux
    port map (
            O => \N__48287\,
            I => \N__47786\
        );

    \I__11500\ : SRMux
    port map (
            O => \N__48286\,
            I => \N__47786\
        );

    \I__11499\ : Glb2LocalMux
    port map (
            O => \N__48283\,
            I => \N__47786\
        );

    \I__11498\ : SRMux
    port map (
            O => \N__48282\,
            I => \N__47786\
        );

    \I__11497\ : SRMux
    port map (
            O => \N__48281\,
            I => \N__47786\
        );

    \I__11496\ : SRMux
    port map (
            O => \N__48280\,
            I => \N__47786\
        );

    \I__11495\ : SRMux
    port map (
            O => \N__48279\,
            I => \N__47786\
        );

    \I__11494\ : SRMux
    port map (
            O => \N__48278\,
            I => \N__47786\
        );

    \I__11493\ : SRMux
    port map (
            O => \N__48277\,
            I => \N__47786\
        );

    \I__11492\ : SRMux
    port map (
            O => \N__48276\,
            I => \N__47786\
        );

    \I__11491\ : SRMux
    port map (
            O => \N__48275\,
            I => \N__47786\
        );

    \I__11490\ : SRMux
    port map (
            O => \N__48274\,
            I => \N__47786\
        );

    \I__11489\ : SRMux
    port map (
            O => \N__48273\,
            I => \N__47786\
        );

    \I__11488\ : SRMux
    port map (
            O => \N__48272\,
            I => \N__47786\
        );

    \I__11487\ : SRMux
    port map (
            O => \N__48271\,
            I => \N__47786\
        );

    \I__11486\ : SRMux
    port map (
            O => \N__48270\,
            I => \N__47786\
        );

    \I__11485\ : SRMux
    port map (
            O => \N__48269\,
            I => \N__47786\
        );

    \I__11484\ : SRMux
    port map (
            O => \N__48268\,
            I => \N__47786\
        );

    \I__11483\ : SRMux
    port map (
            O => \N__48267\,
            I => \N__47786\
        );

    \I__11482\ : SRMux
    port map (
            O => \N__48266\,
            I => \N__47786\
        );

    \I__11481\ : SRMux
    port map (
            O => \N__48265\,
            I => \N__47786\
        );

    \I__11480\ : SRMux
    port map (
            O => \N__48264\,
            I => \N__47786\
        );

    \I__11479\ : SRMux
    port map (
            O => \N__48263\,
            I => \N__47786\
        );

    \I__11478\ : SRMux
    port map (
            O => \N__48262\,
            I => \N__47786\
        );

    \I__11477\ : SRMux
    port map (
            O => \N__48261\,
            I => \N__47786\
        );

    \I__11476\ : SRMux
    port map (
            O => \N__48260\,
            I => \N__47786\
        );

    \I__11475\ : SRMux
    port map (
            O => \N__48259\,
            I => \N__47786\
        );

    \I__11474\ : SRMux
    port map (
            O => \N__48258\,
            I => \N__47786\
        );

    \I__11473\ : SRMux
    port map (
            O => \N__48257\,
            I => \N__47786\
        );

    \I__11472\ : SRMux
    port map (
            O => \N__48256\,
            I => \N__47786\
        );

    \I__11471\ : SRMux
    port map (
            O => \N__48255\,
            I => \N__47786\
        );

    \I__11470\ : SRMux
    port map (
            O => \N__48254\,
            I => \N__47786\
        );

    \I__11469\ : SRMux
    port map (
            O => \N__48253\,
            I => \N__47786\
        );

    \I__11468\ : SRMux
    port map (
            O => \N__48252\,
            I => \N__47786\
        );

    \I__11467\ : SRMux
    port map (
            O => \N__48251\,
            I => \N__47786\
        );

    \I__11466\ : SRMux
    port map (
            O => \N__48250\,
            I => \N__47786\
        );

    \I__11465\ : SRMux
    port map (
            O => \N__48249\,
            I => \N__47786\
        );

    \I__11464\ : SRMux
    port map (
            O => \N__48248\,
            I => \N__47786\
        );

    \I__11463\ : SRMux
    port map (
            O => \N__48247\,
            I => \N__47786\
        );

    \I__11462\ : SRMux
    port map (
            O => \N__48246\,
            I => \N__47786\
        );

    \I__11461\ : SRMux
    port map (
            O => \N__48245\,
            I => \N__47786\
        );

    \I__11460\ : SRMux
    port map (
            O => \N__48244\,
            I => \N__47786\
        );

    \I__11459\ : SRMux
    port map (
            O => \N__48243\,
            I => \N__47786\
        );

    \I__11458\ : SRMux
    port map (
            O => \N__48242\,
            I => \N__47786\
        );

    \I__11457\ : SRMux
    port map (
            O => \N__48241\,
            I => \N__47786\
        );

    \I__11456\ : SRMux
    port map (
            O => \N__48240\,
            I => \N__47786\
        );

    \I__11455\ : SRMux
    port map (
            O => \N__48239\,
            I => \N__47786\
        );

    \I__11454\ : SRMux
    port map (
            O => \N__48238\,
            I => \N__47786\
        );

    \I__11453\ : SRMux
    port map (
            O => \N__48237\,
            I => \N__47786\
        );

    \I__11452\ : SRMux
    port map (
            O => \N__48236\,
            I => \N__47786\
        );

    \I__11451\ : SRMux
    port map (
            O => \N__48235\,
            I => \N__47786\
        );

    \I__11450\ : SRMux
    port map (
            O => \N__48234\,
            I => \N__47786\
        );

    \I__11449\ : SRMux
    port map (
            O => \N__48233\,
            I => \N__47786\
        );

    \I__11448\ : SRMux
    port map (
            O => \N__48232\,
            I => \N__47786\
        );

    \I__11447\ : SRMux
    port map (
            O => \N__48231\,
            I => \N__47786\
        );

    \I__11446\ : SRMux
    port map (
            O => \N__48230\,
            I => \N__47786\
        );

    \I__11445\ : SRMux
    port map (
            O => \N__48229\,
            I => \N__47786\
        );

    \I__11444\ : SRMux
    port map (
            O => \N__48228\,
            I => \N__47786\
        );

    \I__11443\ : SRMux
    port map (
            O => \N__48227\,
            I => \N__47786\
        );

    \I__11442\ : SRMux
    port map (
            O => \N__48226\,
            I => \N__47786\
        );

    \I__11441\ : SRMux
    port map (
            O => \N__48225\,
            I => \N__47786\
        );

    \I__11440\ : SRMux
    port map (
            O => \N__48224\,
            I => \N__47786\
        );

    \I__11439\ : SRMux
    port map (
            O => \N__48223\,
            I => \N__47786\
        );

    \I__11438\ : SRMux
    port map (
            O => \N__48222\,
            I => \N__47786\
        );

    \I__11437\ : SRMux
    port map (
            O => \N__48221\,
            I => \N__47786\
        );

    \I__11436\ : SRMux
    port map (
            O => \N__48220\,
            I => \N__47786\
        );

    \I__11435\ : SRMux
    port map (
            O => \N__48219\,
            I => \N__47786\
        );

    \I__11434\ : SRMux
    port map (
            O => \N__48218\,
            I => \N__47786\
        );

    \I__11433\ : SRMux
    port map (
            O => \N__48217\,
            I => \N__47786\
        );

    \I__11432\ : SRMux
    port map (
            O => \N__48216\,
            I => \N__47786\
        );

    \I__11431\ : SRMux
    port map (
            O => \N__48215\,
            I => \N__47786\
        );

    \I__11430\ : SRMux
    port map (
            O => \N__48214\,
            I => \N__47786\
        );

    \I__11429\ : SRMux
    port map (
            O => \N__48213\,
            I => \N__47786\
        );

    \I__11428\ : SRMux
    port map (
            O => \N__48212\,
            I => \N__47786\
        );

    \I__11427\ : SRMux
    port map (
            O => \N__48211\,
            I => \N__47786\
        );

    \I__11426\ : SRMux
    port map (
            O => \N__48210\,
            I => \N__47786\
        );

    \I__11425\ : SRMux
    port map (
            O => \N__48209\,
            I => \N__47786\
        );

    \I__11424\ : SRMux
    port map (
            O => \N__48208\,
            I => \N__47786\
        );

    \I__11423\ : SRMux
    port map (
            O => \N__48207\,
            I => \N__47786\
        );

    \I__11422\ : SRMux
    port map (
            O => \N__48206\,
            I => \N__47786\
        );

    \I__11421\ : SRMux
    port map (
            O => \N__48205\,
            I => \N__47786\
        );

    \I__11420\ : SRMux
    port map (
            O => \N__48204\,
            I => \N__47786\
        );

    \I__11419\ : SRMux
    port map (
            O => \N__48203\,
            I => \N__47786\
        );

    \I__11418\ : SRMux
    port map (
            O => \N__48202\,
            I => \N__47786\
        );

    \I__11417\ : SRMux
    port map (
            O => \N__48201\,
            I => \N__47786\
        );

    \I__11416\ : SRMux
    port map (
            O => \N__48200\,
            I => \N__47786\
        );

    \I__11415\ : SRMux
    port map (
            O => \N__48199\,
            I => \N__47786\
        );

    \I__11414\ : SRMux
    port map (
            O => \N__48198\,
            I => \N__47786\
        );

    \I__11413\ : SRMux
    port map (
            O => \N__48197\,
            I => \N__47786\
        );

    \I__11412\ : SRMux
    port map (
            O => \N__48196\,
            I => \N__47786\
        );

    \I__11411\ : SRMux
    port map (
            O => \N__48195\,
            I => \N__47786\
        );

    \I__11410\ : SRMux
    port map (
            O => \N__48194\,
            I => \N__47786\
        );

    \I__11409\ : SRMux
    port map (
            O => \N__48193\,
            I => \N__47786\
        );

    \I__11408\ : SRMux
    port map (
            O => \N__48192\,
            I => \N__47786\
        );

    \I__11407\ : SRMux
    port map (
            O => \N__48191\,
            I => \N__47786\
        );

    \I__11406\ : SRMux
    port map (
            O => \N__48190\,
            I => \N__47786\
        );

    \I__11405\ : SRMux
    port map (
            O => \N__48189\,
            I => \N__47786\
        );

    \I__11404\ : SRMux
    port map (
            O => \N__48188\,
            I => \N__47786\
        );

    \I__11403\ : SRMux
    port map (
            O => \N__48187\,
            I => \N__47786\
        );

    \I__11402\ : SRMux
    port map (
            O => \N__48186\,
            I => \N__47786\
        );

    \I__11401\ : SRMux
    port map (
            O => \N__48185\,
            I => \N__47786\
        );

    \I__11400\ : SRMux
    port map (
            O => \N__48184\,
            I => \N__47786\
        );

    \I__11399\ : SRMux
    port map (
            O => \N__48183\,
            I => \N__47786\
        );

    \I__11398\ : SRMux
    port map (
            O => \N__48182\,
            I => \N__47786\
        );

    \I__11397\ : SRMux
    port map (
            O => \N__48181\,
            I => \N__47786\
        );

    \I__11396\ : SRMux
    port map (
            O => \N__48180\,
            I => \N__47786\
        );

    \I__11395\ : SRMux
    port map (
            O => \N__48179\,
            I => \N__47786\
        );

    \I__11394\ : SRMux
    port map (
            O => \N__48178\,
            I => \N__47786\
        );

    \I__11393\ : SRMux
    port map (
            O => \N__48177\,
            I => \N__47786\
        );

    \I__11392\ : SRMux
    port map (
            O => \N__48176\,
            I => \N__47786\
        );

    \I__11391\ : SRMux
    port map (
            O => \N__48175\,
            I => \N__47786\
        );

    \I__11390\ : SRMux
    port map (
            O => \N__48174\,
            I => \N__47786\
        );

    \I__11389\ : SRMux
    port map (
            O => \N__48173\,
            I => \N__47786\
        );

    \I__11388\ : SRMux
    port map (
            O => \N__48172\,
            I => \N__47786\
        );

    \I__11387\ : SRMux
    port map (
            O => \N__48171\,
            I => \N__47786\
        );

    \I__11386\ : SRMux
    port map (
            O => \N__48170\,
            I => \N__47786\
        );

    \I__11385\ : SRMux
    port map (
            O => \N__48169\,
            I => \N__47786\
        );

    \I__11384\ : SRMux
    port map (
            O => \N__48168\,
            I => \N__47786\
        );

    \I__11383\ : SRMux
    port map (
            O => \N__48167\,
            I => \N__47786\
        );

    \I__11382\ : SRMux
    port map (
            O => \N__48166\,
            I => \N__47786\
        );

    \I__11381\ : SRMux
    port map (
            O => \N__48165\,
            I => \N__47786\
        );

    \I__11380\ : SRMux
    port map (
            O => \N__48164\,
            I => \N__47786\
        );

    \I__11379\ : SRMux
    port map (
            O => \N__48163\,
            I => \N__47786\
        );

    \I__11378\ : SRMux
    port map (
            O => \N__48162\,
            I => \N__47786\
        );

    \I__11377\ : SRMux
    port map (
            O => \N__48161\,
            I => \N__47786\
        );

    \I__11376\ : SRMux
    port map (
            O => \N__48160\,
            I => \N__47786\
        );

    \I__11375\ : SRMux
    port map (
            O => \N__48159\,
            I => \N__47786\
        );

    \I__11374\ : SRMux
    port map (
            O => \N__48158\,
            I => \N__47786\
        );

    \I__11373\ : SRMux
    port map (
            O => \N__48157\,
            I => \N__47786\
        );

    \I__11372\ : SRMux
    port map (
            O => \N__48156\,
            I => \N__47786\
        );

    \I__11371\ : SRMux
    port map (
            O => \N__48155\,
            I => \N__47786\
        );

    \I__11370\ : SRMux
    port map (
            O => \N__48154\,
            I => \N__47786\
        );

    \I__11369\ : SRMux
    port map (
            O => \N__48153\,
            I => \N__47786\
        );

    \I__11368\ : SRMux
    port map (
            O => \N__48152\,
            I => \N__47786\
        );

    \I__11367\ : SRMux
    port map (
            O => \N__48151\,
            I => \N__47786\
        );

    \I__11366\ : SRMux
    port map (
            O => \N__48150\,
            I => \N__47786\
        );

    \I__11365\ : SRMux
    port map (
            O => \N__48149\,
            I => \N__47786\
        );

    \I__11364\ : SRMux
    port map (
            O => \N__48148\,
            I => \N__47786\
        );

    \I__11363\ : SRMux
    port map (
            O => \N__48147\,
            I => \N__47786\
        );

    \I__11362\ : SRMux
    port map (
            O => \N__48146\,
            I => \N__47786\
        );

    \I__11361\ : SRMux
    port map (
            O => \N__48145\,
            I => \N__47786\
        );

    \I__11360\ : SRMux
    port map (
            O => \N__48144\,
            I => \N__47786\
        );

    \I__11359\ : SRMux
    port map (
            O => \N__48143\,
            I => \N__47786\
        );

    \I__11358\ : SRMux
    port map (
            O => \N__48142\,
            I => \N__47786\
        );

    \I__11357\ : SRMux
    port map (
            O => \N__48141\,
            I => \N__47786\
        );

    \I__11356\ : SRMux
    port map (
            O => \N__48140\,
            I => \N__47786\
        );

    \I__11355\ : SRMux
    port map (
            O => \N__48139\,
            I => \N__47786\
        );

    \I__11354\ : SRMux
    port map (
            O => \N__48138\,
            I => \N__47786\
        );

    \I__11353\ : SRMux
    port map (
            O => \N__48137\,
            I => \N__47786\
        );

    \I__11352\ : SRMux
    port map (
            O => \N__48136\,
            I => \N__47786\
        );

    \I__11351\ : SRMux
    port map (
            O => \N__48135\,
            I => \N__47786\
        );

    \I__11350\ : SRMux
    port map (
            O => \N__48134\,
            I => \N__47786\
        );

    \I__11349\ : SRMux
    port map (
            O => \N__48133\,
            I => \N__47786\
        );

    \I__11348\ : SRMux
    port map (
            O => \N__48132\,
            I => \N__47786\
        );

    \I__11347\ : SRMux
    port map (
            O => \N__48131\,
            I => \N__47786\
        );

    \I__11346\ : SRMux
    port map (
            O => \N__48130\,
            I => \N__47786\
        );

    \I__11345\ : SRMux
    port map (
            O => \N__48129\,
            I => \N__47786\
        );

    \I__11344\ : SRMux
    port map (
            O => \N__48128\,
            I => \N__47786\
        );

    \I__11343\ : SRMux
    port map (
            O => \N__48127\,
            I => \N__47786\
        );

    \I__11342\ : SRMux
    port map (
            O => \N__48126\,
            I => \N__47786\
        );

    \I__11341\ : SRMux
    port map (
            O => \N__48125\,
            I => \N__47786\
        );

    \I__11340\ : SRMux
    port map (
            O => \N__48124\,
            I => \N__47786\
        );

    \I__11339\ : SRMux
    port map (
            O => \N__48123\,
            I => \N__47786\
        );

    \I__11338\ : SRMux
    port map (
            O => \N__48122\,
            I => \N__47786\
        );

    \I__11337\ : SRMux
    port map (
            O => \N__48121\,
            I => \N__47786\
        );

    \I__11336\ : GlobalMux
    port map (
            O => \N__47786\,
            I => \N__47783\
        );

    \I__11335\ : gio2CtrlBuf
    port map (
            O => \N__47783\,
            I => red_c_g
        );

    \I__11334\ : InMux
    port map (
            O => \N__47780\,
            I => \N__47777\
        );

    \I__11333\ : LocalMux
    port map (
            O => \N__47777\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__11332\ : InMux
    port map (
            O => \N__47774\,
            I => \N__47765\
        );

    \I__11331\ : InMux
    port map (
            O => \N__47773\,
            I => \N__47765\
        );

    \I__11330\ : InMux
    port map (
            O => \N__47772\,
            I => \N__47765\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__47765\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__11328\ : CascadeMux
    port map (
            O => \N__47762\,
            I => \N__47759\
        );

    \I__11327\ : InMux
    port map (
            O => \N__47759\,
            I => \N__47754\
        );

    \I__11326\ : InMux
    port map (
            O => \N__47758\,
            I => \N__47749\
        );

    \I__11325\ : InMux
    port map (
            O => \N__47757\,
            I => \N__47749\
        );

    \I__11324\ : LocalMux
    port map (
            O => \N__47754\,
            I => \N__47746\
        );

    \I__11323\ : LocalMux
    port map (
            O => \N__47749\,
            I => \N__47743\
        );

    \I__11322\ : Span4Mux_v
    port map (
            O => \N__47746\,
            I => \N__47740\
        );

    \I__11321\ : Span4Mux_h
    port map (
            O => \N__47743\,
            I => \N__47737\
        );

    \I__11320\ : Sp12to4
    port map (
            O => \N__47740\,
            I => \N__47734\
        );

    \I__11319\ : Span4Mux_h
    port map (
            O => \N__47737\,
            I => \N__47731\
        );

    \I__11318\ : Odrv12
    port map (
            O => \N__47734\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__11317\ : Odrv4
    port map (
            O => \N__47731\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__11316\ : InMux
    port map (
            O => \N__47726\,
            I => \N__47723\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__47723\,
            I => \N__47718\
        );

    \I__11314\ : InMux
    port map (
            O => \N__47722\,
            I => \N__47713\
        );

    \I__11313\ : InMux
    port map (
            O => \N__47721\,
            I => \N__47713\
        );

    \I__11312\ : Span4Mux_s0_h
    port map (
            O => \N__47718\,
            I => \N__47710\
        );

    \I__11311\ : LocalMux
    port map (
            O => \N__47713\,
            I => pwm_duty_input_7
        );

    \I__11310\ : Odrv4
    port map (
            O => \N__47710\,
            I => pwm_duty_input_7
        );

    \I__11309\ : CascadeMux
    port map (
            O => \N__47705\,
            I => \N__47701\
        );

    \I__11308\ : CascadeMux
    port map (
            O => \N__47704\,
            I => \N__47698\
        );

    \I__11307\ : InMux
    port map (
            O => \N__47701\,
            I => \N__47695\
        );

    \I__11306\ : InMux
    port map (
            O => \N__47698\,
            I => \N__47692\
        );

    \I__11305\ : LocalMux
    port map (
            O => \N__47695\,
            I => \N__47688\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__47692\,
            I => \N__47685\
        );

    \I__11303\ : InMux
    port map (
            O => \N__47691\,
            I => \N__47682\
        );

    \I__11302\ : Span4Mux_h
    port map (
            O => \N__47688\,
            I => \N__47679\
        );

    \I__11301\ : Span12Mux_s1_h
    port map (
            O => \N__47685\,
            I => \N__47674\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__47682\,
            I => \N__47674\
        );

    \I__11299\ : Span4Mux_h
    port map (
            O => \N__47679\,
            I => \N__47671\
        );

    \I__11298\ : Odrv12
    port map (
            O => \N__47674\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__11297\ : Odrv4
    port map (
            O => \N__47671\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__11296\ : InMux
    port map (
            O => \N__47666\,
            I => \N__47661\
        );

    \I__11295\ : InMux
    port map (
            O => \N__47665\,
            I => \N__47656\
        );

    \I__11294\ : InMux
    port map (
            O => \N__47664\,
            I => \N__47656\
        );

    \I__11293\ : LocalMux
    port map (
            O => \N__47661\,
            I => \N__47653\
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__47656\,
            I => pwm_duty_input_8
        );

    \I__11291\ : Odrv4
    port map (
            O => \N__47653\,
            I => pwm_duty_input_8
        );

    \I__11290\ : InMux
    port map (
            O => \N__47648\,
            I => \N__47645\
        );

    \I__11289\ : LocalMux
    port map (
            O => \N__47645\,
            I => \N__47642\
        );

    \I__11288\ : Span4Mux_h
    port map (
            O => \N__47642\,
            I => \N__47639\
        );

    \I__11287\ : Odrv4
    port map (
            O => \N__47639\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__11286\ : InMux
    port map (
            O => \N__47636\,
            I => \N__47632\
        );

    \I__11285\ : InMux
    port map (
            O => \N__47635\,
            I => \N__47629\
        );

    \I__11284\ : LocalMux
    port map (
            O => \N__47632\,
            I => \N__47626\
        );

    \I__11283\ : LocalMux
    port map (
            O => \N__47629\,
            I => pwm_duty_input_0
        );

    \I__11282\ : Odrv4
    port map (
            O => \N__47626\,
            I => pwm_duty_input_0
        );

    \I__11281\ : InMux
    port map (
            O => \N__47621\,
            I => \N__47617\
        );

    \I__11280\ : InMux
    port map (
            O => \N__47620\,
            I => \N__47614\
        );

    \I__11279\ : LocalMux
    port map (
            O => \N__47617\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__11278\ : LocalMux
    port map (
            O => \N__47614\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__11277\ : InMux
    port map (
            O => \N__47609\,
            I => \N__47606\
        );

    \I__11276\ : LocalMux
    port map (
            O => \N__47606\,
            I => \N__47601\
        );

    \I__11275\ : InMux
    port map (
            O => \N__47605\,
            I => \N__47598\
        );

    \I__11274\ : InMux
    port map (
            O => \N__47604\,
            I => \N__47595\
        );

    \I__11273\ : Span4Mux_v
    port map (
            O => \N__47601\,
            I => \N__47590\
        );

    \I__11272\ : LocalMux
    port map (
            O => \N__47598\,
            I => \N__47590\
        );

    \I__11271\ : LocalMux
    port map (
            O => \N__47595\,
            I => \N__47587\
        );

    \I__11270\ : Span4Mux_h
    port map (
            O => \N__47590\,
            I => \N__47584\
        );

    \I__11269\ : Span12Mux_s4_h
    port map (
            O => \N__47587\,
            I => \N__47581\
        );

    \I__11268\ : Span4Mux_h
    port map (
            O => \N__47584\,
            I => \N__47578\
        );

    \I__11267\ : Odrv12
    port map (
            O => \N__47581\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__11266\ : Odrv4
    port map (
            O => \N__47578\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__11265\ : InMux
    port map (
            O => \N__47573\,
            I => \N__47568\
        );

    \I__11264\ : InMux
    port map (
            O => \N__47572\,
            I => \N__47565\
        );

    \I__11263\ : InMux
    port map (
            O => \N__47571\,
            I => \N__47562\
        );

    \I__11262\ : LocalMux
    port map (
            O => \N__47568\,
            I => \N__47559\
        );

    \I__11261\ : LocalMux
    port map (
            O => \N__47565\,
            I => \N__47556\
        );

    \I__11260\ : LocalMux
    port map (
            O => \N__47562\,
            I => \N__47553\
        );

    \I__11259\ : Odrv4
    port map (
            O => \N__47559\,
            I => pwm_duty_input_3
        );

    \I__11258\ : Odrv4
    port map (
            O => \N__47556\,
            I => pwm_duty_input_3
        );

    \I__11257\ : Odrv4
    port map (
            O => \N__47553\,
            I => pwm_duty_input_3
        );

    \I__11256\ : InMux
    port map (
            O => \N__47546\,
            I => \N__47532\
        );

    \I__11255\ : InMux
    port map (
            O => \N__47545\,
            I => \N__47532\
        );

    \I__11254\ : InMux
    port map (
            O => \N__47544\,
            I => \N__47517\
        );

    \I__11253\ : InMux
    port map (
            O => \N__47543\,
            I => \N__47517\
        );

    \I__11252\ : InMux
    port map (
            O => \N__47542\,
            I => \N__47517\
        );

    \I__11251\ : InMux
    port map (
            O => \N__47541\,
            I => \N__47517\
        );

    \I__11250\ : InMux
    port map (
            O => \N__47540\,
            I => \N__47517\
        );

    \I__11249\ : InMux
    port map (
            O => \N__47539\,
            I => \N__47517\
        );

    \I__11248\ : InMux
    port map (
            O => \N__47538\,
            I => \N__47517\
        );

    \I__11247\ : InMux
    port map (
            O => \N__47537\,
            I => \N__47514\
        );

    \I__11246\ : LocalMux
    port map (
            O => \N__47532\,
            I => \N__47509\
        );

    \I__11245\ : LocalMux
    port map (
            O => \N__47517\,
            I => \N__47509\
        );

    \I__11244\ : LocalMux
    port map (
            O => \N__47514\,
            I => \N__47504\
        );

    \I__11243\ : Span12Mux_s7_v
    port map (
            O => \N__47509\,
            I => \N__47504\
        );

    \I__11242\ : Odrv12
    port map (
            O => \N__47504\,
            I => \pwm_generator_inst.N_16\
        );

    \I__11241\ : InMux
    port map (
            O => \N__47501\,
            I => \N__47498\
        );

    \I__11240\ : LocalMux
    port map (
            O => \N__47498\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4\
        );

    \I__11239\ : CascadeMux
    port map (
            O => \N__47495\,
            I => \current_shift_inst.PI_CTRL.N_27_cascade_\
        );

    \I__11238\ : InMux
    port map (
            O => \N__47492\,
            I => \N__47489\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__47489\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\
        );

    \I__11236\ : InMux
    port map (
            O => \N__47486\,
            I => \N__47483\
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__47483\,
            I => \current_shift_inst.PI_CTRL.N_98\
        );

    \I__11234\ : CascadeMux
    port map (
            O => \N__47480\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\
        );

    \I__11233\ : InMux
    port map (
            O => \N__47477\,
            I => \N__47464\
        );

    \I__11232\ : InMux
    port map (
            O => \N__47476\,
            I => \N__47464\
        );

    \I__11231\ : InMux
    port map (
            O => \N__47475\,
            I => \N__47448\
        );

    \I__11230\ : InMux
    port map (
            O => \N__47474\,
            I => \N__47448\
        );

    \I__11229\ : InMux
    port map (
            O => \N__47473\,
            I => \N__47448\
        );

    \I__11228\ : InMux
    port map (
            O => \N__47472\,
            I => \N__47448\
        );

    \I__11227\ : InMux
    port map (
            O => \N__47471\,
            I => \N__47448\
        );

    \I__11226\ : InMux
    port map (
            O => \N__47470\,
            I => \N__47448\
        );

    \I__11225\ : InMux
    port map (
            O => \N__47469\,
            I => \N__47448\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__47464\,
            I => \N__47445\
        );

    \I__11223\ : InMux
    port map (
            O => \N__47463\,
            I => \N__47442\
        );

    \I__11222\ : LocalMux
    port map (
            O => \N__47448\,
            I => \N__47439\
        );

    \I__11221\ : Span4Mux_v
    port map (
            O => \N__47445\,
            I => \N__47434\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__47442\,
            I => \N__47434\
        );

    \I__11219\ : Span4Mux_h
    port map (
            O => \N__47439\,
            I => \N__47431\
        );

    \I__11218\ : Span4Mux_h
    port map (
            O => \N__47434\,
            I => \N__47428\
        );

    \I__11217\ : Span4Mux_h
    port map (
            O => \N__47431\,
            I => \N__47425\
        );

    \I__11216\ : Sp12to4
    port map (
            O => \N__47428\,
            I => \N__47422\
        );

    \I__11215\ : Span4Mux_h
    port map (
            O => \N__47425\,
            I => \N__47419\
        );

    \I__11214\ : Odrv12
    port map (
            O => \N__47422\,
            I => \pwm_generator_inst.N_17\
        );

    \I__11213\ : Odrv4
    port map (
            O => \N__47419\,
            I => \pwm_generator_inst.N_17\
        );

    \I__11212\ : CascadeMux
    port map (
            O => \N__47414\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\
        );

    \I__11211\ : InMux
    port map (
            O => \N__47411\,
            I => \N__47408\
        );

    \I__11210\ : LocalMux
    port map (
            O => \N__47408\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\
        );

    \I__11209\ : CascadeMux
    port map (
            O => \N__47405\,
            I => \N__47401\
        );

    \I__11208\ : InMux
    port map (
            O => \N__47404\,
            I => \N__47396\
        );

    \I__11207\ : InMux
    port map (
            O => \N__47401\,
            I => \N__47396\
        );

    \I__11206\ : LocalMux
    port map (
            O => \N__47396\,
            I => \N__47392\
        );

    \I__11205\ : InMux
    port map (
            O => \N__47395\,
            I => \N__47389\
        );

    \I__11204\ : Span4Mux_h
    port map (
            O => \N__47392\,
            I => \N__47386\
        );

    \I__11203\ : LocalMux
    port map (
            O => \N__47389\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__11202\ : Odrv4
    port map (
            O => \N__47386\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__11201\ : CascadeMux
    port map (
            O => \N__47381\,
            I => \N__47377\
        );

    \I__11200\ : InMux
    port map (
            O => \N__47380\,
            I => \N__47372\
        );

    \I__11199\ : InMux
    port map (
            O => \N__47377\,
            I => \N__47372\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__47372\,
            I => \N__47368\
        );

    \I__11197\ : InMux
    port map (
            O => \N__47371\,
            I => \N__47365\
        );

    \I__11196\ : Span4Mux_h
    port map (
            O => \N__47368\,
            I => \N__47362\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__47365\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__11194\ : Odrv4
    port map (
            O => \N__47362\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__11193\ : InMux
    port map (
            O => \N__47357\,
            I => \N__47354\
        );

    \I__11192\ : LocalMux
    port map (
            O => \N__47354\,
            I => \N__47351\
        );

    \I__11191\ : Odrv4
    port map (
            O => \N__47351\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\
        );

    \I__11190\ : InMux
    port map (
            O => \N__47348\,
            I => \N__47343\
        );

    \I__11189\ : InMux
    port map (
            O => \N__47347\,
            I => \N__47340\
        );

    \I__11188\ : InMux
    port map (
            O => \N__47346\,
            I => \N__47337\
        );

    \I__11187\ : LocalMux
    port map (
            O => \N__47343\,
            I => \N__47334\
        );

    \I__11186\ : LocalMux
    port map (
            O => \N__47340\,
            I => \N__47331\
        );

    \I__11185\ : LocalMux
    port map (
            O => \N__47337\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__11184\ : Odrv12
    port map (
            O => \N__47334\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__11183\ : Odrv4
    port map (
            O => \N__47331\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__11182\ : InMux
    port map (
            O => \N__47324\,
            I => \N__47320\
        );

    \I__11181\ : InMux
    port map (
            O => \N__47323\,
            I => \N__47316\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__47320\,
            I => \N__47313\
        );

    \I__11179\ : InMux
    port map (
            O => \N__47319\,
            I => \N__47310\
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__47316\,
            I => \N__47307\
        );

    \I__11177\ : Span4Mux_h
    port map (
            O => \N__47313\,
            I => \N__47304\
        );

    \I__11176\ : LocalMux
    port map (
            O => \N__47310\,
            I => \N__47299\
        );

    \I__11175\ : Span4Mux_h
    port map (
            O => \N__47307\,
            I => \N__47299\
        );

    \I__11174\ : Span4Mux_h
    port map (
            O => \N__47304\,
            I => \N__47295\
        );

    \I__11173\ : Span4Mux_h
    port map (
            O => \N__47299\,
            I => \N__47292\
        );

    \I__11172\ : InMux
    port map (
            O => \N__47298\,
            I => \N__47289\
        );

    \I__11171\ : Odrv4
    port map (
            O => \N__47295\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__11170\ : Odrv4
    port map (
            O => \N__47292\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__11169\ : LocalMux
    port map (
            O => \N__47289\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__11168\ : InMux
    port map (
            O => \N__47282\,
            I => \N__47276\
        );

    \I__11167\ : InMux
    port map (
            O => \N__47281\,
            I => \N__47276\
        );

    \I__11166\ : LocalMux
    port map (
            O => \N__47276\,
            I => \N__47273\
        );

    \I__11165\ : Odrv12
    port map (
            O => \N__47273\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\
        );

    \I__11164\ : InMux
    port map (
            O => \N__47270\,
            I => \N__47266\
        );

    \I__11163\ : InMux
    port map (
            O => \N__47269\,
            I => \N__47263\
        );

    \I__11162\ : LocalMux
    port map (
            O => \N__47266\,
            I => \N__47260\
        );

    \I__11161\ : LocalMux
    port map (
            O => \N__47263\,
            I => \N__47257\
        );

    \I__11160\ : Sp12to4
    port map (
            O => \N__47260\,
            I => \N__47254\
        );

    \I__11159\ : Span4Mux_v
    port map (
            O => \N__47257\,
            I => \N__47251\
        );

    \I__11158\ : Span12Mux_v
    port map (
            O => \N__47254\,
            I => \N__47248\
        );

    \I__11157\ : Sp12to4
    port map (
            O => \N__47251\,
            I => \N__47245\
        );

    \I__11156\ : Odrv12
    port map (
            O => \N__47248\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__11155\ : Odrv12
    port map (
            O => \N__47245\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__11154\ : InMux
    port map (
            O => \N__47240\,
            I => \N__47237\
        );

    \I__11153\ : LocalMux
    port map (
            O => \N__47237\,
            I => \N__47234\
        );

    \I__11152\ : Odrv4
    port map (
            O => \N__47234\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__11151\ : InMux
    port map (
            O => \N__47231\,
            I => \N__47227\
        );

    \I__11150\ : InMux
    port map (
            O => \N__47230\,
            I => \N__47223\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__47227\,
            I => \N__47220\
        );

    \I__11148\ : InMux
    port map (
            O => \N__47226\,
            I => \N__47217\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__47223\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__11146\ : Odrv12
    port map (
            O => \N__47220\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__11145\ : LocalMux
    port map (
            O => \N__47217\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__11144\ : InMux
    port map (
            O => \N__47210\,
            I => \N__47206\
        );

    \I__11143\ : InMux
    port map (
            O => \N__47209\,
            I => \N__47202\
        );

    \I__11142\ : LocalMux
    port map (
            O => \N__47206\,
            I => \N__47199\
        );

    \I__11141\ : InMux
    port map (
            O => \N__47205\,
            I => \N__47196\
        );

    \I__11140\ : LocalMux
    port map (
            O => \N__47202\,
            I => \N__47192\
        );

    \I__11139\ : Span4Mux_h
    port map (
            O => \N__47199\,
            I => \N__47189\
        );

    \I__11138\ : LocalMux
    port map (
            O => \N__47196\,
            I => \N__47186\
        );

    \I__11137\ : CascadeMux
    port map (
            O => \N__47195\,
            I => \N__47183\
        );

    \I__11136\ : Span4Mux_v
    port map (
            O => \N__47192\,
            I => \N__47178\
        );

    \I__11135\ : Span4Mux_h
    port map (
            O => \N__47189\,
            I => \N__47178\
        );

    \I__11134\ : Span12Mux_v
    port map (
            O => \N__47186\,
            I => \N__47175\
        );

    \I__11133\ : InMux
    port map (
            O => \N__47183\,
            I => \N__47172\
        );

    \I__11132\ : Odrv4
    port map (
            O => \N__47178\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__11131\ : Odrv12
    port map (
            O => \N__47175\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__11130\ : LocalMux
    port map (
            O => \N__47172\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__11129\ : InMux
    port map (
            O => \N__47165\,
            I => \N__47157\
        );

    \I__11128\ : InMux
    port map (
            O => \N__47164\,
            I => \N__47154\
        );

    \I__11127\ : InMux
    port map (
            O => \N__47163\,
            I => \N__47151\
        );

    \I__11126\ : InMux
    port map (
            O => \N__47162\,
            I => \N__47148\
        );

    \I__11125\ : InMux
    port map (
            O => \N__47161\,
            I => \N__47125\
        );

    \I__11124\ : InMux
    port map (
            O => \N__47160\,
            I => \N__47125\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__47157\,
            I => \N__47103\
        );

    \I__11122\ : LocalMux
    port map (
            O => \N__47154\,
            I => \N__47096\
        );

    \I__11121\ : LocalMux
    port map (
            O => \N__47151\,
            I => \N__47096\
        );

    \I__11120\ : LocalMux
    port map (
            O => \N__47148\,
            I => \N__47096\
        );

    \I__11119\ : InMux
    port map (
            O => \N__47147\,
            I => \N__47091\
        );

    \I__11118\ : InMux
    port map (
            O => \N__47146\,
            I => \N__47091\
        );

    \I__11117\ : CascadeMux
    port map (
            O => \N__47145\,
            I => \N__47085\
        );

    \I__11116\ : InMux
    port map (
            O => \N__47144\,
            I => \N__47072\
        );

    \I__11115\ : InMux
    port map (
            O => \N__47143\,
            I => \N__47072\
        );

    \I__11114\ : InMux
    port map (
            O => \N__47142\,
            I => \N__47072\
        );

    \I__11113\ : InMux
    port map (
            O => \N__47141\,
            I => \N__47072\
        );

    \I__11112\ : InMux
    port map (
            O => \N__47140\,
            I => \N__47067\
        );

    \I__11111\ : InMux
    port map (
            O => \N__47139\,
            I => \N__47067\
        );

    \I__11110\ : InMux
    port map (
            O => \N__47138\,
            I => \N__47048\
        );

    \I__11109\ : InMux
    port map (
            O => \N__47137\,
            I => \N__47045\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47136\,
            I => \N__47034\
        );

    \I__11107\ : InMux
    port map (
            O => \N__47135\,
            I => \N__47034\
        );

    \I__11106\ : InMux
    port map (
            O => \N__47134\,
            I => \N__47034\
        );

    \I__11105\ : InMux
    port map (
            O => \N__47133\,
            I => \N__47034\
        );

    \I__11104\ : InMux
    port map (
            O => \N__47132\,
            I => \N__47034\
        );

    \I__11103\ : InMux
    port map (
            O => \N__47131\,
            I => \N__47029\
        );

    \I__11102\ : InMux
    port map (
            O => \N__47130\,
            I => \N__47029\
        );

    \I__11101\ : LocalMux
    port map (
            O => \N__47125\,
            I => \N__47026\
        );

    \I__11100\ : InMux
    port map (
            O => \N__47124\,
            I => \N__47021\
        );

    \I__11099\ : InMux
    port map (
            O => \N__47123\,
            I => \N__47021\
        );

    \I__11098\ : InMux
    port map (
            O => \N__47122\,
            I => \N__47018\
        );

    \I__11097\ : InMux
    port map (
            O => \N__47121\,
            I => \N__47013\
        );

    \I__11096\ : InMux
    port map (
            O => \N__47120\,
            I => \N__47013\
        );

    \I__11095\ : InMux
    port map (
            O => \N__47119\,
            I => \N__47004\
        );

    \I__11094\ : InMux
    port map (
            O => \N__47118\,
            I => \N__47004\
        );

    \I__11093\ : InMux
    port map (
            O => \N__47117\,
            I => \N__47004\
        );

    \I__11092\ : InMux
    port map (
            O => \N__47116\,
            I => \N__47004\
        );

    \I__11091\ : InMux
    port map (
            O => \N__47115\,
            I => \N__46995\
        );

    \I__11090\ : InMux
    port map (
            O => \N__47114\,
            I => \N__46995\
        );

    \I__11089\ : InMux
    port map (
            O => \N__47113\,
            I => \N__46995\
        );

    \I__11088\ : InMux
    port map (
            O => \N__47112\,
            I => \N__46995\
        );

    \I__11087\ : InMux
    port map (
            O => \N__47111\,
            I => \N__46985\
        );

    \I__11086\ : InMux
    port map (
            O => \N__47110\,
            I => \N__46985\
        );

    \I__11085\ : InMux
    port map (
            O => \N__47109\,
            I => \N__46978\
        );

    \I__11084\ : InMux
    port map (
            O => \N__47108\,
            I => \N__46978\
        );

    \I__11083\ : InMux
    port map (
            O => \N__47107\,
            I => \N__46978\
        );

    \I__11082\ : InMux
    port map (
            O => \N__47106\,
            I => \N__46971\
        );

    \I__11081\ : Span4Mux_v
    port map (
            O => \N__47103\,
            I => \N__46964\
        );

    \I__11080\ : Span4Mux_v
    port map (
            O => \N__47096\,
            I => \N__46964\
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__47091\,
            I => \N__46964\
        );

    \I__11078\ : InMux
    port map (
            O => \N__47090\,
            I => \N__46957\
        );

    \I__11077\ : InMux
    port map (
            O => \N__47089\,
            I => \N__46957\
        );

    \I__11076\ : InMux
    port map (
            O => \N__47088\,
            I => \N__46957\
        );

    \I__11075\ : InMux
    port map (
            O => \N__47085\,
            I => \N__46954\
        );

    \I__11074\ : InMux
    port map (
            O => \N__47084\,
            I => \N__46949\
        );

    \I__11073\ : InMux
    port map (
            O => \N__47083\,
            I => \N__46949\
        );

    \I__11072\ : InMux
    port map (
            O => \N__47082\,
            I => \N__46946\
        );

    \I__11071\ : InMux
    port map (
            O => \N__47081\,
            I => \N__46943\
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__47072\,
            I => \N__46940\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__47067\,
            I => \N__46937\
        );

    \I__11068\ : InMux
    port map (
            O => \N__47066\,
            I => \N__46916\
        );

    \I__11067\ : InMux
    port map (
            O => \N__47065\,
            I => \N__46916\
        );

    \I__11066\ : InMux
    port map (
            O => \N__47064\,
            I => \N__46907\
        );

    \I__11065\ : InMux
    port map (
            O => \N__47063\,
            I => \N__46907\
        );

    \I__11064\ : InMux
    port map (
            O => \N__47062\,
            I => \N__46907\
        );

    \I__11063\ : InMux
    port map (
            O => \N__47061\,
            I => \N__46907\
        );

    \I__11062\ : InMux
    port map (
            O => \N__47060\,
            I => \N__46900\
        );

    \I__11061\ : InMux
    port map (
            O => \N__47059\,
            I => \N__46900\
        );

    \I__11060\ : InMux
    port map (
            O => \N__47058\,
            I => \N__46900\
        );

    \I__11059\ : InMux
    port map (
            O => \N__47057\,
            I => \N__46893\
        );

    \I__11058\ : InMux
    port map (
            O => \N__47056\,
            I => \N__46893\
        );

    \I__11057\ : InMux
    port map (
            O => \N__47055\,
            I => \N__46893\
        );

    \I__11056\ : InMux
    port map (
            O => \N__47054\,
            I => \N__46884\
        );

    \I__11055\ : InMux
    port map (
            O => \N__47053\,
            I => \N__46884\
        );

    \I__11054\ : InMux
    port map (
            O => \N__47052\,
            I => \N__46884\
        );

    \I__11053\ : InMux
    port map (
            O => \N__47051\,
            I => \N__46884\
        );

    \I__11052\ : LocalMux
    port map (
            O => \N__47048\,
            I => \N__46877\
        );

    \I__11051\ : LocalMux
    port map (
            O => \N__47045\,
            I => \N__46877\
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__47034\,
            I => \N__46877\
        );

    \I__11049\ : LocalMux
    port map (
            O => \N__47029\,
            I => \N__46870\
        );

    \I__11048\ : Span4Mux_v
    port map (
            O => \N__47026\,
            I => \N__46870\
        );

    \I__11047\ : LocalMux
    port map (
            O => \N__47021\,
            I => \N__46870\
        );

    \I__11046\ : LocalMux
    port map (
            O => \N__47018\,
            I => \N__46861\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__47013\,
            I => \N__46861\
        );

    \I__11044\ : LocalMux
    port map (
            O => \N__47004\,
            I => \N__46861\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__46995\,
            I => \N__46861\
        );

    \I__11042\ : InMux
    port map (
            O => \N__46994\,
            I => \N__46850\
        );

    \I__11041\ : InMux
    port map (
            O => \N__46993\,
            I => \N__46850\
        );

    \I__11040\ : InMux
    port map (
            O => \N__46992\,
            I => \N__46850\
        );

    \I__11039\ : InMux
    port map (
            O => \N__46991\,
            I => \N__46850\
        );

    \I__11038\ : InMux
    port map (
            O => \N__46990\,
            I => \N__46850\
        );

    \I__11037\ : LocalMux
    port map (
            O => \N__46985\,
            I => \N__46845\
        );

    \I__11036\ : LocalMux
    port map (
            O => \N__46978\,
            I => \N__46845\
        );

    \I__11035\ : InMux
    port map (
            O => \N__46977\,
            I => \N__46842\
        );

    \I__11034\ : InMux
    port map (
            O => \N__46976\,
            I => \N__46834\
        );

    \I__11033\ : InMux
    port map (
            O => \N__46975\,
            I => \N__46834\
        );

    \I__11032\ : InMux
    port map (
            O => \N__46974\,
            I => \N__46834\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__46971\,
            I => \N__46823\
        );

    \I__11030\ : Span4Mux_h
    port map (
            O => \N__46964\,
            I => \N__46823\
        );

    \I__11029\ : LocalMux
    port map (
            O => \N__46957\,
            I => \N__46823\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__46954\,
            I => \N__46823\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__46949\,
            I => \N__46823\
        );

    \I__11026\ : LocalMux
    port map (
            O => \N__46946\,
            I => \N__46814\
        );

    \I__11025\ : LocalMux
    port map (
            O => \N__46943\,
            I => \N__46814\
        );

    \I__11024\ : Span4Mux_h
    port map (
            O => \N__46940\,
            I => \N__46814\
        );

    \I__11023\ : Span4Mux_h
    port map (
            O => \N__46937\,
            I => \N__46814\
        );

    \I__11022\ : InMux
    port map (
            O => \N__46936\,
            I => \N__46811\
        );

    \I__11021\ : InMux
    port map (
            O => \N__46935\,
            I => \N__46808\
        );

    \I__11020\ : InMux
    port map (
            O => \N__46934\,
            I => \N__46801\
        );

    \I__11019\ : InMux
    port map (
            O => \N__46933\,
            I => \N__46801\
        );

    \I__11018\ : InMux
    port map (
            O => \N__46932\,
            I => \N__46801\
        );

    \I__11017\ : InMux
    port map (
            O => \N__46931\,
            I => \N__46796\
        );

    \I__11016\ : InMux
    port map (
            O => \N__46930\,
            I => \N__46796\
        );

    \I__11015\ : InMux
    port map (
            O => \N__46929\,
            I => \N__46785\
        );

    \I__11014\ : InMux
    port map (
            O => \N__46928\,
            I => \N__46785\
        );

    \I__11013\ : InMux
    port map (
            O => \N__46927\,
            I => \N__46785\
        );

    \I__11012\ : InMux
    port map (
            O => \N__46926\,
            I => \N__46785\
        );

    \I__11011\ : InMux
    port map (
            O => \N__46925\,
            I => \N__46785\
        );

    \I__11010\ : InMux
    port map (
            O => \N__46924\,
            I => \N__46776\
        );

    \I__11009\ : InMux
    port map (
            O => \N__46923\,
            I => \N__46776\
        );

    \I__11008\ : InMux
    port map (
            O => \N__46922\,
            I => \N__46776\
        );

    \I__11007\ : InMux
    port map (
            O => \N__46921\,
            I => \N__46776\
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__46916\,
            I => \N__46773\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__46907\,
            I => \N__46764\
        );

    \I__11004\ : LocalMux
    port map (
            O => \N__46900\,
            I => \N__46764\
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__46893\,
            I => \N__46764\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__46884\,
            I => \N__46764\
        );

    \I__11001\ : Span4Mux_v
    port map (
            O => \N__46877\,
            I => \N__46757\
        );

    \I__11000\ : Span4Mux_v
    port map (
            O => \N__46870\,
            I => \N__46757\
        );

    \I__10999\ : Span4Mux_v
    port map (
            O => \N__46861\,
            I => \N__46757\
        );

    \I__10998\ : LocalMux
    port map (
            O => \N__46850\,
            I => \N__46750\
        );

    \I__10997\ : Span12Mux_v
    port map (
            O => \N__46845\,
            I => \N__46750\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__46842\,
            I => \N__46750\
        );

    \I__10995\ : InMux
    port map (
            O => \N__46841\,
            I => \N__46747\
        );

    \I__10994\ : LocalMux
    port map (
            O => \N__46834\,
            I => \N__46740\
        );

    \I__10993\ : Span4Mux_v
    port map (
            O => \N__46823\,
            I => \N__46740\
        );

    \I__10992\ : Span4Mux_v
    port map (
            O => \N__46814\,
            I => \N__46740\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__46811\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__46808\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__46801\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__46796\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__10987\ : LocalMux
    port map (
            O => \N__46785\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__10986\ : LocalMux
    port map (
            O => \N__46776\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__10985\ : Odrv4
    port map (
            O => \N__46773\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__10984\ : Odrv4
    port map (
            O => \N__46764\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__10983\ : Odrv4
    port map (
            O => \N__46757\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__10982\ : Odrv12
    port map (
            O => \N__46750\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__10981\ : LocalMux
    port map (
            O => \N__46747\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__10980\ : Odrv4
    port map (
            O => \N__46740\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__10979\ : InMux
    port map (
            O => \N__46715\,
            I => \N__46709\
        );

    \I__10978\ : InMux
    port map (
            O => \N__46714\,
            I => \N__46709\
        );

    \I__10977\ : LocalMux
    port map (
            O => \N__46709\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\
        );

    \I__10976\ : CEMux
    port map (
            O => \N__46706\,
            I => \N__46703\
        );

    \I__10975\ : LocalMux
    port map (
            O => \N__46703\,
            I => \N__46691\
        );

    \I__10974\ : CEMux
    port map (
            O => \N__46702\,
            I => \N__46688\
        );

    \I__10973\ : InMux
    port map (
            O => \N__46701\,
            I => \N__46672\
        );

    \I__10972\ : CEMux
    port map (
            O => \N__46700\,
            I => \N__46669\
        );

    \I__10971\ : CEMux
    port map (
            O => \N__46699\,
            I => \N__46666\
        );

    \I__10970\ : CEMux
    port map (
            O => \N__46698\,
            I => \N__46658\
        );

    \I__10969\ : InMux
    port map (
            O => \N__46697\,
            I => \N__46648\
        );

    \I__10968\ : InMux
    port map (
            O => \N__46696\,
            I => \N__46648\
        );

    \I__10967\ : InMux
    port map (
            O => \N__46695\,
            I => \N__46648\
        );

    \I__10966\ : InMux
    port map (
            O => \N__46694\,
            I => \N__46648\
        );

    \I__10965\ : Span4Mux_v
    port map (
            O => \N__46691\,
            I => \N__46643\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__46688\,
            I => \N__46643\
        );

    \I__10963\ : CEMux
    port map (
            O => \N__46687\,
            I => \N__46640\
        );

    \I__10962\ : CEMux
    port map (
            O => \N__46686\,
            I => \N__46637\
        );

    \I__10961\ : InMux
    port map (
            O => \N__46685\,
            I => \N__46628\
        );

    \I__10960\ : InMux
    port map (
            O => \N__46684\,
            I => \N__46628\
        );

    \I__10959\ : InMux
    port map (
            O => \N__46683\,
            I => \N__46628\
        );

    \I__10958\ : InMux
    port map (
            O => \N__46682\,
            I => \N__46628\
        );

    \I__10957\ : InMux
    port map (
            O => \N__46681\,
            I => \N__46619\
        );

    \I__10956\ : InMux
    port map (
            O => \N__46680\,
            I => \N__46619\
        );

    \I__10955\ : InMux
    port map (
            O => \N__46679\,
            I => \N__46619\
        );

    \I__10954\ : InMux
    port map (
            O => \N__46678\,
            I => \N__46619\
        );

    \I__10953\ : CEMux
    port map (
            O => \N__46677\,
            I => \N__46616\
        );

    \I__10952\ : CEMux
    port map (
            O => \N__46676\,
            I => \N__46611\
        );

    \I__10951\ : CEMux
    port map (
            O => \N__46675\,
            I => \N__46598\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__46672\,
            I => \N__46595\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__46669\,
            I => \N__46586\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__46666\,
            I => \N__46583\
        );

    \I__10947\ : CEMux
    port map (
            O => \N__46665\,
            I => \N__46580\
        );

    \I__10946\ : InMux
    port map (
            O => \N__46664\,
            I => \N__46571\
        );

    \I__10945\ : InMux
    port map (
            O => \N__46663\,
            I => \N__46571\
        );

    \I__10944\ : InMux
    port map (
            O => \N__46662\,
            I => \N__46571\
        );

    \I__10943\ : InMux
    port map (
            O => \N__46661\,
            I => \N__46571\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__46658\,
            I => \N__46568\
        );

    \I__10941\ : CEMux
    port map (
            O => \N__46657\,
            I => \N__46565\
        );

    \I__10940\ : LocalMux
    port map (
            O => \N__46648\,
            I => \N__46562\
        );

    \I__10939\ : Span4Mux_h
    port map (
            O => \N__46643\,
            I => \N__46557\
        );

    \I__10938\ : LocalMux
    port map (
            O => \N__46640\,
            I => \N__46557\
        );

    \I__10937\ : LocalMux
    port map (
            O => \N__46637\,
            I => \N__46554\
        );

    \I__10936\ : LocalMux
    port map (
            O => \N__46628\,
            I => \N__46547\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__46619\,
            I => \N__46547\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__46616\,
            I => \N__46547\
        );

    \I__10933\ : CEMux
    port map (
            O => \N__46615\,
            I => \N__46544\
        );

    \I__10932\ : CEMux
    port map (
            O => \N__46614\,
            I => \N__46541\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__46611\,
            I => \N__46538\
        );

    \I__10930\ : InMux
    port map (
            O => \N__46610\,
            I => \N__46531\
        );

    \I__10929\ : InMux
    port map (
            O => \N__46609\,
            I => \N__46531\
        );

    \I__10928\ : InMux
    port map (
            O => \N__46608\,
            I => \N__46531\
        );

    \I__10927\ : InMux
    port map (
            O => \N__46607\,
            I => \N__46522\
        );

    \I__10926\ : InMux
    port map (
            O => \N__46606\,
            I => \N__46522\
        );

    \I__10925\ : InMux
    port map (
            O => \N__46605\,
            I => \N__46522\
        );

    \I__10924\ : InMux
    port map (
            O => \N__46604\,
            I => \N__46522\
        );

    \I__10923\ : InMux
    port map (
            O => \N__46603\,
            I => \N__46515\
        );

    \I__10922\ : InMux
    port map (
            O => \N__46602\,
            I => \N__46515\
        );

    \I__10921\ : InMux
    port map (
            O => \N__46601\,
            I => \N__46515\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__46598\,
            I => \N__46512\
        );

    \I__10919\ : Span4Mux_h
    port map (
            O => \N__46595\,
            I => \N__46509\
        );

    \I__10918\ : InMux
    port map (
            O => \N__46594\,
            I => \N__46500\
        );

    \I__10917\ : InMux
    port map (
            O => \N__46593\,
            I => \N__46500\
        );

    \I__10916\ : InMux
    port map (
            O => \N__46592\,
            I => \N__46500\
        );

    \I__10915\ : InMux
    port map (
            O => \N__46591\,
            I => \N__46500\
        );

    \I__10914\ : CEMux
    port map (
            O => \N__46590\,
            I => \N__46497\
        );

    \I__10913\ : CEMux
    port map (
            O => \N__46589\,
            I => \N__46494\
        );

    \I__10912\ : Span4Mux_h
    port map (
            O => \N__46586\,
            I => \N__46477\
        );

    \I__10911\ : Span4Mux_h
    port map (
            O => \N__46583\,
            I => \N__46477\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__46580\,
            I => \N__46477\
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__46571\,
            I => \N__46477\
        );

    \I__10908\ : Span4Mux_v
    port map (
            O => \N__46568\,
            I => \N__46477\
        );

    \I__10907\ : LocalMux
    port map (
            O => \N__46565\,
            I => \N__46477\
        );

    \I__10906\ : Span4Mux_h
    port map (
            O => \N__46562\,
            I => \N__46477\
        );

    \I__10905\ : Span4Mux_v
    port map (
            O => \N__46557\,
            I => \N__46477\
        );

    \I__10904\ : Span4Mux_v
    port map (
            O => \N__46554\,
            I => \N__46474\
        );

    \I__10903\ : Span4Mux_h
    port map (
            O => \N__46547\,
            I => \N__46471\
        );

    \I__10902\ : LocalMux
    port map (
            O => \N__46544\,
            I => \N__46468\
        );

    \I__10901\ : LocalMux
    port map (
            O => \N__46541\,
            I => \N__46465\
        );

    \I__10900\ : Span4Mux_v
    port map (
            O => \N__46538\,
            I => \N__46454\
        );

    \I__10899\ : LocalMux
    port map (
            O => \N__46531\,
            I => \N__46454\
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__46522\,
            I => \N__46454\
        );

    \I__10897\ : LocalMux
    port map (
            O => \N__46515\,
            I => \N__46454\
        );

    \I__10896\ : Span4Mux_h
    port map (
            O => \N__46512\,
            I => \N__46454\
        );

    \I__10895\ : Span4Mux_v
    port map (
            O => \N__46509\,
            I => \N__46451\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__46500\,
            I => \N__46448\
        );

    \I__10893\ : LocalMux
    port map (
            O => \N__46497\,
            I => \N__46439\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__46494\,
            I => \N__46439\
        );

    \I__10891\ : Span4Mux_v
    port map (
            O => \N__46477\,
            I => \N__46439\
        );

    \I__10890\ : Span4Mux_s3_h
    port map (
            O => \N__46474\,
            I => \N__46439\
        );

    \I__10889\ : Span4Mux_v
    port map (
            O => \N__46471\,
            I => \N__46436\
        );

    \I__10888\ : Span4Mux_h
    port map (
            O => \N__46468\,
            I => \N__46427\
        );

    \I__10887\ : Span4Mux_h
    port map (
            O => \N__46465\,
            I => \N__46427\
        );

    \I__10886\ : Span4Mux_v
    port map (
            O => \N__46454\,
            I => \N__46427\
        );

    \I__10885\ : Span4Mux_h
    port map (
            O => \N__46451\,
            I => \N__46427\
        );

    \I__10884\ : Span4Mux_v
    port map (
            O => \N__46448\,
            I => \N__46422\
        );

    \I__10883\ : Span4Mux_h
    port map (
            O => \N__46439\,
            I => \N__46422\
        );

    \I__10882\ : Odrv4
    port map (
            O => \N__46436\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__10881\ : Odrv4
    port map (
            O => \N__46427\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__10880\ : Odrv4
    port map (
            O => \N__46422\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__10879\ : CascadeMux
    port map (
            O => \N__46415\,
            I => \N__46410\
        );

    \I__10878\ : CascadeMux
    port map (
            O => \N__46414\,
            I => \N__46407\
        );

    \I__10877\ : InMux
    port map (
            O => \N__46413\,
            I => \N__46400\
        );

    \I__10876\ : InMux
    port map (
            O => \N__46410\,
            I => \N__46400\
        );

    \I__10875\ : InMux
    port map (
            O => \N__46407\,
            I => \N__46400\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__46400\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__10873\ : InMux
    port map (
            O => \N__46397\,
            I => \N__46391\
        );

    \I__10872\ : InMux
    port map (
            O => \N__46396\,
            I => \N__46388\
        );

    \I__10871\ : InMux
    port map (
            O => \N__46395\,
            I => \N__46385\
        );

    \I__10870\ : InMux
    port map (
            O => \N__46394\,
            I => \N__46382\
        );

    \I__10869\ : LocalMux
    port map (
            O => \N__46391\,
            I => \N__46379\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__46388\,
            I => \N__46374\
        );

    \I__10867\ : LocalMux
    port map (
            O => \N__46385\,
            I => \N__46374\
        );

    \I__10866\ : LocalMux
    port map (
            O => \N__46382\,
            I => \N__46371\
        );

    \I__10865\ : Span4Mux_h
    port map (
            O => \N__46379\,
            I => \N__46368\
        );

    \I__10864\ : Span4Mux_h
    port map (
            O => \N__46374\,
            I => \N__46365\
        );

    \I__10863\ : Span4Mux_v
    port map (
            O => \N__46371\,
            I => \N__46362\
        );

    \I__10862\ : Odrv4
    port map (
            O => \N__46368\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__10861\ : Odrv4
    port map (
            O => \N__46365\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__10860\ : Odrv4
    port map (
            O => \N__46362\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__10859\ : InMux
    port map (
            O => \N__46355\,
            I => \N__46350\
        );

    \I__10858\ : InMux
    port map (
            O => \N__46354\,
            I => \N__46347\
        );

    \I__10857\ : InMux
    port map (
            O => \N__46353\,
            I => \N__46344\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__46350\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__46347\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__46344\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__10853\ : InMux
    port map (
            O => \N__46337\,
            I => \N__46332\
        );

    \I__10852\ : InMux
    port map (
            O => \N__46336\,
            I => \N__46329\
        );

    \I__10851\ : InMux
    port map (
            O => \N__46335\,
            I => \N__46326\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__46332\,
            I => \N__46323\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__46329\,
            I => \N__46320\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__46326\,
            I => \N__46316\
        );

    \I__10847\ : Span4Mux_h
    port map (
            O => \N__46323\,
            I => \N__46313\
        );

    \I__10846\ : Span4Mux_h
    port map (
            O => \N__46320\,
            I => \N__46310\
        );

    \I__10845\ : InMux
    port map (
            O => \N__46319\,
            I => \N__46307\
        );

    \I__10844\ : Odrv4
    port map (
            O => \N__46316\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__10843\ : Odrv4
    port map (
            O => \N__46313\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__10842\ : Odrv4
    port map (
            O => \N__46310\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__46307\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__10840\ : InMux
    port map (
            O => \N__46298\,
            I => \N__46295\
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__46295\,
            I => \N__46292\
        );

    \I__10838\ : Span4Mux_h
    port map (
            O => \N__46292\,
            I => \N__46288\
        );

    \I__10837\ : InMux
    port map (
            O => \N__46291\,
            I => \N__46284\
        );

    \I__10836\ : Span4Mux_h
    port map (
            O => \N__46288\,
            I => \N__46281\
        );

    \I__10835\ : InMux
    port map (
            O => \N__46287\,
            I => \N__46278\
        );

    \I__10834\ : LocalMux
    port map (
            O => \N__46284\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__10833\ : Odrv4
    port map (
            O => \N__46281\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__46278\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__10831\ : InMux
    port map (
            O => \N__46271\,
            I => \N__46268\
        );

    \I__10830\ : LocalMux
    port map (
            O => \N__46268\,
            I => \N__46264\
        );

    \I__10829\ : InMux
    port map (
            O => \N__46267\,
            I => \N__46261\
        );

    \I__10828\ : Sp12to4
    port map (
            O => \N__46264\,
            I => \N__46256\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__46261\,
            I => \N__46256\
        );

    \I__10826\ : Odrv12
    port map (
            O => \N__46256\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__10825\ : CascadeMux
    port map (
            O => \N__46253\,
            I => \N__46250\
        );

    \I__10824\ : InMux
    port map (
            O => \N__46250\,
            I => \N__46247\
        );

    \I__10823\ : LocalMux
    port map (
            O => \N__46247\,
            I => \N__46243\
        );

    \I__10822\ : InMux
    port map (
            O => \N__46246\,
            I => \N__46239\
        );

    \I__10821\ : Span4Mux_v
    port map (
            O => \N__46243\,
            I => \N__46235\
        );

    \I__10820\ : InMux
    port map (
            O => \N__46242\,
            I => \N__46232\
        );

    \I__10819\ : LocalMux
    port map (
            O => \N__46239\,
            I => \N__46229\
        );

    \I__10818\ : InMux
    port map (
            O => \N__46238\,
            I => \N__46225\
        );

    \I__10817\ : Span4Mux_v
    port map (
            O => \N__46235\,
            I => \N__46222\
        );

    \I__10816\ : LocalMux
    port map (
            O => \N__46232\,
            I => \N__46219\
        );

    \I__10815\ : Span4Mux_v
    port map (
            O => \N__46229\,
            I => \N__46216\
        );

    \I__10814\ : InMux
    port map (
            O => \N__46228\,
            I => \N__46213\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__46225\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__10812\ : Odrv4
    port map (
            O => \N__46222\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__10811\ : Odrv12
    port map (
            O => \N__46219\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__10810\ : Odrv4
    port map (
            O => \N__46216\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__46213\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__10808\ : InMux
    port map (
            O => \N__46202\,
            I => \N__46198\
        );

    \I__10807\ : InMux
    port map (
            O => \N__46201\,
            I => \N__46195\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__46198\,
            I => \N__46192\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__46195\,
            I => \N__46186\
        );

    \I__10804\ : Span4Mux_h
    port map (
            O => \N__46192\,
            I => \N__46183\
        );

    \I__10803\ : InMux
    port map (
            O => \N__46191\,
            I => \N__46178\
        );

    \I__10802\ : InMux
    port map (
            O => \N__46190\,
            I => \N__46178\
        );

    \I__10801\ : InMux
    port map (
            O => \N__46189\,
            I => \N__46175\
        );

    \I__10800\ : Span12Mux_s9_h
    port map (
            O => \N__46186\,
            I => \N__46168\
        );

    \I__10799\ : Sp12to4
    port map (
            O => \N__46183\,
            I => \N__46168\
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__46178\,
            I => \N__46168\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__46175\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__10796\ : Odrv12
    port map (
            O => \N__46168\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__10795\ : InMux
    port map (
            O => \N__46163\,
            I => \N__46160\
        );

    \I__10794\ : LocalMux
    port map (
            O => \N__46160\,
            I => \N__46156\
        );

    \I__10793\ : InMux
    port map (
            O => \N__46159\,
            I => \N__46153\
        );

    \I__10792\ : Span4Mux_v
    port map (
            O => \N__46156\,
            I => \N__46150\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__46153\,
            I => \N__46146\
        );

    \I__10790\ : Span4Mux_v
    port map (
            O => \N__46150\,
            I => \N__46143\
        );

    \I__10789\ : InMux
    port map (
            O => \N__46149\,
            I => \N__46140\
        );

    \I__10788\ : Span4Mux_v
    port map (
            O => \N__46146\,
            I => \N__46137\
        );

    \I__10787\ : Odrv4
    port map (
            O => \N__46143\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__10786\ : LocalMux
    port map (
            O => \N__46140\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__10785\ : Odrv4
    port map (
            O => \N__46137\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__10784\ : InMux
    port map (
            O => \N__46130\,
            I => \N__46124\
        );

    \I__10783\ : InMux
    port map (
            O => \N__46129\,
            I => \N__46124\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__46124\,
            I => \N__46121\
        );

    \I__10781\ : Odrv12
    port map (
            O => \N__46121\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\
        );

    \I__10780\ : CEMux
    port map (
            O => \N__46118\,
            I => \N__46082\
        );

    \I__10779\ : CEMux
    port map (
            O => \N__46117\,
            I => \N__46082\
        );

    \I__10778\ : CEMux
    port map (
            O => \N__46116\,
            I => \N__46082\
        );

    \I__10777\ : CEMux
    port map (
            O => \N__46115\,
            I => \N__46082\
        );

    \I__10776\ : CEMux
    port map (
            O => \N__46114\,
            I => \N__46082\
        );

    \I__10775\ : CEMux
    port map (
            O => \N__46113\,
            I => \N__46082\
        );

    \I__10774\ : CEMux
    port map (
            O => \N__46112\,
            I => \N__46082\
        );

    \I__10773\ : CEMux
    port map (
            O => \N__46111\,
            I => \N__46082\
        );

    \I__10772\ : CEMux
    port map (
            O => \N__46110\,
            I => \N__46082\
        );

    \I__10771\ : CEMux
    port map (
            O => \N__46109\,
            I => \N__46082\
        );

    \I__10770\ : CEMux
    port map (
            O => \N__46108\,
            I => \N__46082\
        );

    \I__10769\ : CEMux
    port map (
            O => \N__46107\,
            I => \N__46082\
        );

    \I__10768\ : GlobalMux
    port map (
            O => \N__46082\,
            I => \N__46079\
        );

    \I__10767\ : gio2CtrlBuf
    port map (
            O => \N__46079\,
            I => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \I__10766\ : InMux
    port map (
            O => \N__46076\,
            I => \N__46072\
        );

    \I__10765\ : InMux
    port map (
            O => \N__46075\,
            I => \N__46069\
        );

    \I__10764\ : LocalMux
    port map (
            O => \N__46072\,
            I => \N__46065\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__46069\,
            I => \N__46062\
        );

    \I__10762\ : InMux
    port map (
            O => \N__46068\,
            I => \N__46059\
        );

    \I__10761\ : Span4Mux_h
    port map (
            O => \N__46065\,
            I => \N__46056\
        );

    \I__10760\ : Span4Mux_h
    port map (
            O => \N__46062\,
            I => \N__46053\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__46059\,
            I => \N__46048\
        );

    \I__10758\ : Span4Mux_v
    port map (
            O => \N__46056\,
            I => \N__46048\
        );

    \I__10757\ : Span4Mux_v
    port map (
            O => \N__46053\,
            I => \N__46045\
        );

    \I__10756\ : Span4Mux_h
    port map (
            O => \N__46048\,
            I => \N__46041\
        );

    \I__10755\ : Span4Mux_h
    port map (
            O => \N__46045\,
            I => \N__46038\
        );

    \I__10754\ : InMux
    port map (
            O => \N__46044\,
            I => \N__46035\
        );

    \I__10753\ : Odrv4
    port map (
            O => \N__46041\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__10752\ : Odrv4
    port map (
            O => \N__46038\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__46035\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__10750\ : InMux
    port map (
            O => \N__46028\,
            I => \N__46025\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__46025\,
            I => \N__46021\
        );

    \I__10748\ : InMux
    port map (
            O => \N__46024\,
            I => \N__46017\
        );

    \I__10747\ : Span4Mux_h
    port map (
            O => \N__46021\,
            I => \N__46014\
        );

    \I__10746\ : InMux
    port map (
            O => \N__46020\,
            I => \N__46011\
        );

    \I__10745\ : LocalMux
    port map (
            O => \N__46017\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__10744\ : Odrv4
    port map (
            O => \N__46014\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__46011\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__10742\ : InMux
    port map (
            O => \N__46004\,
            I => \N__46001\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__46001\,
            I => \N__45997\
        );

    \I__10740\ : InMux
    port map (
            O => \N__46000\,
            I => \N__45993\
        );

    \I__10739\ : Span4Mux_h
    port map (
            O => \N__45997\,
            I => \N__45990\
        );

    \I__10738\ : InMux
    port map (
            O => \N__45996\,
            I => \N__45987\
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__45993\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__10736\ : Odrv4
    port map (
            O => \N__45990\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__45987\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__10734\ : InMux
    port map (
            O => \N__45980\,
            I => \N__45977\
        );

    \I__10733\ : LocalMux
    port map (
            O => \N__45977\,
            I => \N__45971\
        );

    \I__10732\ : InMux
    port map (
            O => \N__45976\,
            I => \N__45968\
        );

    \I__10731\ : InMux
    port map (
            O => \N__45975\,
            I => \N__45965\
        );

    \I__10730\ : InMux
    port map (
            O => \N__45974\,
            I => \N__45962\
        );

    \I__10729\ : Span4Mux_h
    port map (
            O => \N__45971\,
            I => \N__45957\
        );

    \I__10728\ : LocalMux
    port map (
            O => \N__45968\,
            I => \N__45957\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__45965\,
            I => \N__45954\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__45962\,
            I => \N__45949\
        );

    \I__10725\ : Span4Mux_h
    port map (
            O => \N__45957\,
            I => \N__45949\
        );

    \I__10724\ : Odrv4
    port map (
            O => \N__45954\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__10723\ : Odrv4
    port map (
            O => \N__45949\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__10722\ : CascadeMux
    port map (
            O => \N__45944\,
            I => \N__45941\
        );

    \I__10721\ : InMux
    port map (
            O => \N__45941\,
            I => \N__45938\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__45938\,
            I => \N__45935\
        );

    \I__10719\ : Odrv4
    port map (
            O => \N__45935\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__10718\ : CascadeMux
    port map (
            O => \N__45932\,
            I => \N__45929\
        );

    \I__10717\ : InMux
    port map (
            O => \N__45929\,
            I => \N__45926\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__45926\,
            I => \N__45923\
        );

    \I__10715\ : Odrv12
    port map (
            O => \N__45923\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt22\
        );

    \I__10714\ : InMux
    port map (
            O => \N__45920\,
            I => \N__45914\
        );

    \I__10713\ : InMux
    port map (
            O => \N__45919\,
            I => \N__45914\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__45914\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\
        );

    \I__10711\ : InMux
    port map (
            O => \N__45911\,
            I => \N__45908\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__45908\,
            I => \N__45904\
        );

    \I__10709\ : InMux
    port map (
            O => \N__45907\,
            I => \N__45901\
        );

    \I__10708\ : Odrv4
    port map (
            O => \N__45904\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\
        );

    \I__10707\ : LocalMux
    port map (
            O => \N__45901\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\
        );

    \I__10706\ : InMux
    port map (
            O => \N__45896\,
            I => \N__45892\
        );

    \I__10705\ : InMux
    port map (
            O => \N__45895\,
            I => \N__45888\
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__45892\,
            I => \N__45885\
        );

    \I__10703\ : InMux
    port map (
            O => \N__45891\,
            I => \N__45882\
        );

    \I__10702\ : LocalMux
    port map (
            O => \N__45888\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10701\ : Odrv4
    port map (
            O => \N__45885\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10700\ : LocalMux
    port map (
            O => \N__45882\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10699\ : CascadeMux
    port map (
            O => \N__45875\,
            I => \N__45870\
        );

    \I__10698\ : CascadeMux
    port map (
            O => \N__45874\,
            I => \N__45867\
        );

    \I__10697\ : InMux
    port map (
            O => \N__45873\,
            I => \N__45864\
        );

    \I__10696\ : InMux
    port map (
            O => \N__45870\,
            I => \N__45861\
        );

    \I__10695\ : InMux
    port map (
            O => \N__45867\,
            I => \N__45858\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__45864\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__45861\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__45858\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10691\ : InMux
    port map (
            O => \N__45851\,
            I => \N__45847\
        );

    \I__10690\ : InMux
    port map (
            O => \N__45850\,
            I => \N__45844\
        );

    \I__10689\ : LocalMux
    port map (
            O => \N__45847\,
            I => \N__45841\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__45844\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\
        );

    \I__10687\ : Odrv4
    port map (
            O => \N__45841\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\
        );

    \I__10686\ : InMux
    port map (
            O => \N__45836\,
            I => \N__45833\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__45833\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\
        );

    \I__10684\ : CascadeMux
    port map (
            O => \N__45830\,
            I => \N__45826\
        );

    \I__10683\ : InMux
    port map (
            O => \N__45829\,
            I => \N__45823\
        );

    \I__10682\ : InMux
    port map (
            O => \N__45826\,
            I => \N__45820\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__45823\,
            I => \N__45817\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__45820\,
            I => \N__45814\
        );

    \I__10679\ : Span4Mux_h
    port map (
            O => \N__45817\,
            I => \N__45811\
        );

    \I__10678\ : Odrv4
    port map (
            O => \N__45814\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt30\
        );

    \I__10677\ : Odrv4
    port map (
            O => \N__45811\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt30\
        );

    \I__10676\ : InMux
    port map (
            O => \N__45806\,
            I => \N__45803\
        );

    \I__10675\ : LocalMux
    port map (
            O => \N__45803\,
            I => \N__45799\
        );

    \I__10674\ : InMux
    port map (
            O => \N__45802\,
            I => \N__45796\
        );

    \I__10673\ : Odrv12
    port map (
            O => \N__45799\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__10672\ : LocalMux
    port map (
            O => \N__45796\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__10671\ : CascadeMux
    port map (
            O => \N__45791\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\
        );

    \I__10670\ : InMux
    port map (
            O => \N__45788\,
            I => \N__45782\
        );

    \I__10669\ : InMux
    port map (
            O => \N__45787\,
            I => \N__45777\
        );

    \I__10668\ : InMux
    port map (
            O => \N__45786\,
            I => \N__45777\
        );

    \I__10667\ : CascadeMux
    port map (
            O => \N__45785\,
            I => \N__45774\
        );

    \I__10666\ : LocalMux
    port map (
            O => \N__45782\,
            I => \N__45771\
        );

    \I__10665\ : LocalMux
    port map (
            O => \N__45777\,
            I => \N__45768\
        );

    \I__10664\ : InMux
    port map (
            O => \N__45774\,
            I => \N__45765\
        );

    \I__10663\ : Span4Mux_h
    port map (
            O => \N__45771\,
            I => \N__45758\
        );

    \I__10662\ : Span4Mux_h
    port map (
            O => \N__45768\,
            I => \N__45758\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__45765\,
            I => \N__45758\
        );

    \I__10660\ : Odrv4
    port map (
            O => \N__45758\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__10659\ : InMux
    port map (
            O => \N__45755\,
            I => \N__45752\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__45752\,
            I => \N__45749\
        );

    \I__10657\ : Odrv4
    port map (
            O => \N__45749\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\
        );

    \I__10656\ : InMux
    port map (
            O => \N__45746\,
            I => \N__45737\
        );

    \I__10655\ : InMux
    port map (
            O => \N__45745\,
            I => \N__45737\
        );

    \I__10654\ : InMux
    port map (
            O => \N__45744\,
            I => \N__45737\
        );

    \I__10653\ : LocalMux
    port map (
            O => \N__45737\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__10652\ : CascadeMux
    port map (
            O => \N__45734\,
            I => \N__45730\
        );

    \I__10651\ : InMux
    port map (
            O => \N__45733\,
            I => \N__45725\
        );

    \I__10650\ : InMux
    port map (
            O => \N__45730\,
            I => \N__45718\
        );

    \I__10649\ : InMux
    port map (
            O => \N__45729\,
            I => \N__45718\
        );

    \I__10648\ : InMux
    port map (
            O => \N__45728\,
            I => \N__45718\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__45725\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__10646\ : LocalMux
    port map (
            O => \N__45718\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__10645\ : InMux
    port map (
            O => \N__45713\,
            I => \N__45707\
        );

    \I__10644\ : InMux
    port map (
            O => \N__45712\,
            I => \N__45700\
        );

    \I__10643\ : InMux
    port map (
            O => \N__45711\,
            I => \N__45700\
        );

    \I__10642\ : InMux
    port map (
            O => \N__45710\,
            I => \N__45700\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__45707\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__45700\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__10639\ : CascadeMux
    port map (
            O => \N__45695\,
            I => \N__45692\
        );

    \I__10638\ : InMux
    port map (
            O => \N__45692\,
            I => \N__45689\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__45689\,
            I => \N__45686\
        );

    \I__10636\ : Span4Mux_h
    port map (
            O => \N__45686\,
            I => \N__45683\
        );

    \I__10635\ : Odrv4
    port map (
            O => \N__45683\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df30\
        );

    \I__10634\ : InMux
    port map (
            O => \N__45680\,
            I => \N__45677\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__45677\,
            I => \N__45674\
        );

    \I__10632\ : Odrv12
    port map (
            O => \N__45674\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__10631\ : CascadeMux
    port map (
            O => \N__45671\,
            I => \N__45668\
        );

    \I__10630\ : InMux
    port map (
            O => \N__45668\,
            I => \N__45665\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__45665\,
            I => \N__45662\
        );

    \I__10628\ : Span4Mux_h
    port map (
            O => \N__45662\,
            I => \N__45659\
        );

    \I__10627\ : Odrv4
    port map (
            O => \N__45659\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt26\
        );

    \I__10626\ : InMux
    port map (
            O => \N__45656\,
            I => \N__45653\
        );

    \I__10625\ : LocalMux
    port map (
            O => \N__45653\,
            I => \N__45650\
        );

    \I__10624\ : Odrv4
    port map (
            O => \N__45650\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\
        );

    \I__10623\ : CascadeMux
    port map (
            O => \N__45647\,
            I => \N__45644\
        );

    \I__10622\ : InMux
    port map (
            O => \N__45644\,
            I => \N__45641\
        );

    \I__10621\ : LocalMux
    port map (
            O => \N__45641\,
            I => \N__45638\
        );

    \I__10620\ : Span4Mux_v
    port map (
            O => \N__45638\,
            I => \N__45635\
        );

    \I__10619\ : Odrv4
    port map (
            O => \N__45635\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt28\
        );

    \I__10618\ : InMux
    port map (
            O => \N__45632\,
            I => \N__45629\
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__45629\,
            I => \N__45626\
        );

    \I__10616\ : Odrv4
    port map (
            O => \N__45626\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\
        );

    \I__10615\ : InMux
    port map (
            O => \N__45623\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_28\
        );

    \I__10614\ : InMux
    port map (
            O => \N__45620\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30\
        );

    \I__10613\ : InMux
    port map (
            O => \N__45617\,
            I => \N__45614\
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__45614\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt24\
        );

    \I__10611\ : CascadeMux
    port map (
            O => \N__45611\,
            I => \N__45607\
        );

    \I__10610\ : InMux
    port map (
            O => \N__45610\,
            I => \N__45603\
        );

    \I__10609\ : InMux
    port map (
            O => \N__45607\,
            I => \N__45598\
        );

    \I__10608\ : InMux
    port map (
            O => \N__45606\,
            I => \N__45598\
        );

    \I__10607\ : LocalMux
    port map (
            O => \N__45603\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__45598\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__10605\ : CascadeMux
    port map (
            O => \N__45593\,
            I => \N__45589\
        );

    \I__10604\ : InMux
    port map (
            O => \N__45592\,
            I => \N__45584\
        );

    \I__10603\ : InMux
    port map (
            O => \N__45589\,
            I => \N__45584\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__45584\,
            I => \N__45581\
        );

    \I__10601\ : Odrv12
    port map (
            O => \N__45581\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\
        );

    \I__10600\ : InMux
    port map (
            O => \N__45578\,
            I => \N__45573\
        );

    \I__10599\ : InMux
    port map (
            O => \N__45577\,
            I => \N__45568\
        );

    \I__10598\ : InMux
    port map (
            O => \N__45576\,
            I => \N__45568\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__45573\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__10596\ : LocalMux
    port map (
            O => \N__45568\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__10595\ : CascadeMux
    port map (
            O => \N__45563\,
            I => \N__45560\
        );

    \I__10594\ : InMux
    port map (
            O => \N__45560\,
            I => \N__45557\
        );

    \I__10593\ : LocalMux
    port map (
            O => \N__45557\,
            I => \N__45554\
        );

    \I__10592\ : Odrv4
    port map (
            O => \N__45554\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\
        );

    \I__10591\ : InMux
    port map (
            O => \N__45551\,
            I => \N__45547\
        );

    \I__10590\ : InMux
    port map (
            O => \N__45550\,
            I => \N__45544\
        );

    \I__10589\ : LocalMux
    port map (
            O => \N__45547\,
            I => \N__45541\
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__45544\,
            I => \N__45535\
        );

    \I__10587\ : Span4Mux_v
    port map (
            O => \N__45541\,
            I => \N__45535\
        );

    \I__10586\ : InMux
    port map (
            O => \N__45540\,
            I => \N__45532\
        );

    \I__10585\ : Odrv4
    port map (
            O => \N__45535\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__45532\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__10583\ : InMux
    port map (
            O => \N__45527\,
            I => \N__45524\
        );

    \I__10582\ : LocalMux
    port map (
            O => \N__45524\,
            I => \N__45519\
        );

    \I__10581\ : InMux
    port map (
            O => \N__45523\,
            I => \N__45516\
        );

    \I__10580\ : InMux
    port map (
            O => \N__45522\,
            I => \N__45513\
        );

    \I__10579\ : Span4Mux_v
    port map (
            O => \N__45519\,
            I => \N__45508\
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__45516\,
            I => \N__45508\
        );

    \I__10577\ : LocalMux
    port map (
            O => \N__45513\,
            I => \N__45504\
        );

    \I__10576\ : Span4Mux_h
    port map (
            O => \N__45508\,
            I => \N__45501\
        );

    \I__10575\ : InMux
    port map (
            O => \N__45507\,
            I => \N__45498\
        );

    \I__10574\ : Odrv12
    port map (
            O => \N__45504\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__10573\ : Odrv4
    port map (
            O => \N__45501\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__10572\ : LocalMux
    port map (
            O => \N__45498\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__10571\ : InMux
    port map (
            O => \N__45491\,
            I => \N__45488\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__45488\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__10569\ : InMux
    port map (
            O => \N__45485\,
            I => \N__45482\
        );

    \I__10568\ : LocalMux
    port map (
            O => \N__45482\,
            I => \N__45479\
        );

    \I__10567\ : Odrv12
    port map (
            O => \N__45479\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__10566\ : InMux
    port map (
            O => \N__45476\,
            I => \N__45472\
        );

    \I__10565\ : InMux
    port map (
            O => \N__45475\,
            I => \N__45469\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__45472\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__45469\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__10562\ : CascadeMux
    port map (
            O => \N__45464\,
            I => \N__45461\
        );

    \I__10561\ : InMux
    port map (
            O => \N__45461\,
            I => \N__45458\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__45458\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__10559\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45451\
        );

    \I__10558\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45448\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__45451\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__45448\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__10555\ : InMux
    port map (
            O => \N__45443\,
            I => \N__45440\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__45440\,
            I => \N__45437\
        );

    \I__10553\ : Span4Mux_h
    port map (
            O => \N__45437\,
            I => \N__45434\
        );

    \I__10552\ : Odrv4
    port map (
            O => \N__45434\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__10551\ : CascadeMux
    port map (
            O => \N__45431\,
            I => \N__45428\
        );

    \I__10550\ : InMux
    port map (
            O => \N__45428\,
            I => \N__45425\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__45425\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__10548\ : InMux
    port map (
            O => \N__45422\,
            I => \N__45418\
        );

    \I__10547\ : InMux
    port map (
            O => \N__45421\,
            I => \N__45415\
        );

    \I__10546\ : LocalMux
    port map (
            O => \N__45418\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__45415\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__10544\ : CascadeMux
    port map (
            O => \N__45410\,
            I => \N__45407\
        );

    \I__10543\ : InMux
    port map (
            O => \N__45407\,
            I => \N__45404\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__45404\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__10541\ : InMux
    port map (
            O => \N__45401\,
            I => \N__45398\
        );

    \I__10540\ : LocalMux
    port map (
            O => \N__45398\,
            I => \N__45395\
        );

    \I__10539\ : Odrv4
    port map (
            O => \N__45395\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__10538\ : InMux
    port map (
            O => \N__45392\,
            I => \N__45388\
        );

    \I__10537\ : InMux
    port map (
            O => \N__45391\,
            I => \N__45385\
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__45388\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__10535\ : LocalMux
    port map (
            O => \N__45385\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__10534\ : CascadeMux
    port map (
            O => \N__45380\,
            I => \N__45377\
        );

    \I__10533\ : InMux
    port map (
            O => \N__45377\,
            I => \N__45374\
        );

    \I__10532\ : LocalMux
    port map (
            O => \N__45374\,
            I => \N__45371\
        );

    \I__10531\ : Odrv4
    port map (
            O => \N__45371\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__10530\ : InMux
    port map (
            O => \N__45368\,
            I => \N__45365\
        );

    \I__10529\ : LocalMux
    port map (
            O => \N__45365\,
            I => \N__45362\
        );

    \I__10528\ : Span4Mux_h
    port map (
            O => \N__45362\,
            I => \N__45359\
        );

    \I__10527\ : Odrv4
    port map (
            O => \N__45359\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\
        );

    \I__10526\ : CascadeMux
    port map (
            O => \N__45356\,
            I => \N__45353\
        );

    \I__10525\ : InMux
    port map (
            O => \N__45353\,
            I => \N__45350\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__45350\,
            I => \N__45347\
        );

    \I__10523\ : Span4Mux_h
    port map (
            O => \N__45347\,
            I => \N__45344\
        );

    \I__10522\ : Odrv4
    port map (
            O => \N__45344\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt16\
        );

    \I__10521\ : InMux
    port map (
            O => \N__45341\,
            I => \N__45338\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__45338\,
            I => \N__45335\
        );

    \I__10519\ : Span4Mux_v
    port map (
            O => \N__45335\,
            I => \N__45332\
        );

    \I__10518\ : Odrv4
    port map (
            O => \N__45332\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\
        );

    \I__10517\ : CascadeMux
    port map (
            O => \N__45329\,
            I => \N__45326\
        );

    \I__10516\ : InMux
    port map (
            O => \N__45326\,
            I => \N__45323\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__45323\,
            I => \N__45320\
        );

    \I__10514\ : Span4Mux_v
    port map (
            O => \N__45320\,
            I => \N__45317\
        );

    \I__10513\ : Odrv4
    port map (
            O => \N__45317\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt18\
        );

    \I__10512\ : InMux
    port map (
            O => \N__45314\,
            I => \N__45311\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__45311\,
            I => \N__45308\
        );

    \I__10510\ : Odrv4
    port map (
            O => \N__45308\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\
        );

    \I__10509\ : CascadeMux
    port map (
            O => \N__45305\,
            I => \N__45302\
        );

    \I__10508\ : InMux
    port map (
            O => \N__45302\,
            I => \N__45299\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__45299\,
            I => \N__45296\
        );

    \I__10506\ : Odrv4
    port map (
            O => \N__45296\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt20\
        );

    \I__10505\ : CascadeMux
    port map (
            O => \N__45293\,
            I => \N__45290\
        );

    \I__10504\ : InMux
    port map (
            O => \N__45290\,
            I => \N__45287\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__45287\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__10502\ : InMux
    port map (
            O => \N__45284\,
            I => \N__45280\
        );

    \I__10501\ : InMux
    port map (
            O => \N__45283\,
            I => \N__45277\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__45280\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__45277\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__10498\ : InMux
    port map (
            O => \N__45272\,
            I => \N__45269\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__45269\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__10496\ : InMux
    port map (
            O => \N__45266\,
            I => \N__45262\
        );

    \I__10495\ : InMux
    port map (
            O => \N__45265\,
            I => \N__45259\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__45262\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__45259\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__10492\ : CascadeMux
    port map (
            O => \N__45254\,
            I => \N__45251\
        );

    \I__10491\ : InMux
    port map (
            O => \N__45251\,
            I => \N__45248\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__45248\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__10489\ : InMux
    port map (
            O => \N__45245\,
            I => \N__45242\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__45242\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__10487\ : InMux
    port map (
            O => \N__45239\,
            I => \N__45236\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__45236\,
            I => \N__45233\
        );

    \I__10485\ : Odrv12
    port map (
            O => \N__45233\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__10484\ : InMux
    port map (
            O => \N__45230\,
            I => \N__45226\
        );

    \I__10483\ : InMux
    port map (
            O => \N__45229\,
            I => \N__45223\
        );

    \I__10482\ : LocalMux
    port map (
            O => \N__45226\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__10481\ : LocalMux
    port map (
            O => \N__45223\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__10480\ : CascadeMux
    port map (
            O => \N__45218\,
            I => \N__45215\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45215\,
            I => \N__45212\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__45212\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__10477\ : InMux
    port map (
            O => \N__45209\,
            I => \N__45206\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__45206\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__10475\ : InMux
    port map (
            O => \N__45203\,
            I => \N__45199\
        );

    \I__10474\ : InMux
    port map (
            O => \N__45202\,
            I => \N__45196\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__45199\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__45196\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__10471\ : CascadeMux
    port map (
            O => \N__45191\,
            I => \N__45188\
        );

    \I__10470\ : InMux
    port map (
            O => \N__45188\,
            I => \N__45185\
        );

    \I__10469\ : LocalMux
    port map (
            O => \N__45185\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__10468\ : InMux
    port map (
            O => \N__45182\,
            I => \N__45179\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__45179\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__10466\ : InMux
    port map (
            O => \N__45176\,
            I => \N__45172\
        );

    \I__10465\ : InMux
    port map (
            O => \N__45175\,
            I => \N__45169\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__45172\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__10463\ : LocalMux
    port map (
            O => \N__45169\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__10462\ : CascadeMux
    port map (
            O => \N__45164\,
            I => \N__45161\
        );

    \I__10461\ : InMux
    port map (
            O => \N__45161\,
            I => \N__45158\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__45158\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__10459\ : InMux
    port map (
            O => \N__45155\,
            I => \N__45152\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__45152\,
            I => \N__45149\
        );

    \I__10457\ : Odrv12
    port map (
            O => \N__45149\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__10456\ : InMux
    port map (
            O => \N__45146\,
            I => \N__45142\
        );

    \I__10455\ : InMux
    port map (
            O => \N__45145\,
            I => \N__45139\
        );

    \I__10454\ : LocalMux
    port map (
            O => \N__45142\,
            I => \N__45136\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__45139\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__10452\ : Odrv4
    port map (
            O => \N__45136\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__10451\ : CascadeMux
    port map (
            O => \N__45131\,
            I => \N__45128\
        );

    \I__10450\ : InMux
    port map (
            O => \N__45128\,
            I => \N__45125\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__45125\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__10448\ : InMux
    port map (
            O => \N__45122\,
            I => \N__45118\
        );

    \I__10447\ : InMux
    port map (
            O => \N__45121\,
            I => \N__45115\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__45118\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__45115\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__10444\ : InMux
    port map (
            O => \N__45110\,
            I => \N__45107\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__45107\,
            I => \N__45104\
        );

    \I__10442\ : Odrv4
    port map (
            O => \N__45104\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__10441\ : CascadeMux
    port map (
            O => \N__45101\,
            I => \N__45098\
        );

    \I__10440\ : InMux
    port map (
            O => \N__45098\,
            I => \N__45095\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__45095\,
            I => \N__45092\
        );

    \I__10438\ : Odrv4
    port map (
            O => \N__45092\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__10437\ : InMux
    port map (
            O => \N__45089\,
            I => \N__45085\
        );

    \I__10436\ : InMux
    port map (
            O => \N__45088\,
            I => \N__45082\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__45085\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__45082\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__10433\ : InMux
    port map (
            O => \N__45077\,
            I => \N__45073\
        );

    \I__10432\ : InMux
    port map (
            O => \N__45076\,
            I => \N__45069\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__45073\,
            I => \N__45066\
        );

    \I__10430\ : InMux
    port map (
            O => \N__45072\,
            I => \N__45063\
        );

    \I__10429\ : LocalMux
    port map (
            O => \N__45069\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__10428\ : Odrv4
    port map (
            O => \N__45066\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__45063\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__10426\ : InMux
    port map (
            O => \N__45056\,
            I => \N__45052\
        );

    \I__10425\ : InMux
    port map (
            O => \N__45055\,
            I => \N__45049\
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__45052\,
            I => \N__45045\
        );

    \I__10423\ : LocalMux
    port map (
            O => \N__45049\,
            I => \N__45042\
        );

    \I__10422\ : InMux
    port map (
            O => \N__45048\,
            I => \N__45039\
        );

    \I__10421\ : Span4Mux_v
    port map (
            O => \N__45045\,
            I => \N__45036\
        );

    \I__10420\ : Span4Mux_h
    port map (
            O => \N__45042\,
            I => \N__45033\
        );

    \I__10419\ : LocalMux
    port map (
            O => \N__45039\,
            I => \N__45030\
        );

    \I__10418\ : Span4Mux_v
    port map (
            O => \N__45036\,
            I => \N__45026\
        );

    \I__10417\ : Span4Mux_v
    port map (
            O => \N__45033\,
            I => \N__45023\
        );

    \I__10416\ : Span12Mux_v
    port map (
            O => \N__45030\,
            I => \N__45020\
        );

    \I__10415\ : InMux
    port map (
            O => \N__45029\,
            I => \N__45017\
        );

    \I__10414\ : Odrv4
    port map (
            O => \N__45026\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__10413\ : Odrv4
    port map (
            O => \N__45023\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__10412\ : Odrv12
    port map (
            O => \N__45020\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__10411\ : LocalMux
    port map (
            O => \N__45017\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__10410\ : InMux
    port map (
            O => \N__45008\,
            I => \N__45005\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__45005\,
            I => \N__44999\
        );

    \I__10408\ : InMux
    port map (
            O => \N__45004\,
            I => \N__44996\
        );

    \I__10407\ : InMux
    port map (
            O => \N__45003\,
            I => \N__44993\
        );

    \I__10406\ : InMux
    port map (
            O => \N__45002\,
            I => \N__44990\
        );

    \I__10405\ : Span4Mux_h
    port map (
            O => \N__44999\,
            I => \N__44987\
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__44996\,
            I => \N__44982\
        );

    \I__10403\ : LocalMux
    port map (
            O => \N__44993\,
            I => \N__44982\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__44990\,
            I => \N__44979\
        );

    \I__10401\ : Span4Mux_v
    port map (
            O => \N__44987\,
            I => \N__44976\
        );

    \I__10400\ : Span4Mux_v
    port map (
            O => \N__44982\,
            I => \N__44971\
        );

    \I__10399\ : Span4Mux_h
    port map (
            O => \N__44979\,
            I => \N__44971\
        );

    \I__10398\ : Odrv4
    port map (
            O => \N__44976\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__10397\ : Odrv4
    port map (
            O => \N__44971\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__10396\ : InMux
    port map (
            O => \N__44966\,
            I => \N__44961\
        );

    \I__10395\ : InMux
    port map (
            O => \N__44965\,
            I => \N__44958\
        );

    \I__10394\ : InMux
    port map (
            O => \N__44964\,
            I => \N__44955\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__44961\,
            I => \N__44952\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__44958\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__44955\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__10390\ : Odrv4
    port map (
            O => \N__44952\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__10389\ : InMux
    port map (
            O => \N__44945\,
            I => \N__44942\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__44942\,
            I => \N__44938\
        );

    \I__10387\ : InMux
    port map (
            O => \N__44941\,
            I => \N__44934\
        );

    \I__10386\ : Span4Mux_h
    port map (
            O => \N__44938\,
            I => \N__44931\
        );

    \I__10385\ : InMux
    port map (
            O => \N__44937\,
            I => \N__44928\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__44934\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__10383\ : Odrv4
    port map (
            O => \N__44931\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__44928\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__10381\ : InMux
    port map (
            O => \N__44921\,
            I => \N__44916\
        );

    \I__10380\ : InMux
    port map (
            O => \N__44920\,
            I => \N__44912\
        );

    \I__10379\ : InMux
    port map (
            O => \N__44919\,
            I => \N__44909\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__44916\,
            I => \N__44906\
        );

    \I__10377\ : InMux
    port map (
            O => \N__44915\,
            I => \N__44903\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__44912\,
            I => \N__44898\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__44909\,
            I => \N__44898\
        );

    \I__10374\ : Span4Mux_v
    port map (
            O => \N__44906\,
            I => \N__44893\
        );

    \I__10373\ : LocalMux
    port map (
            O => \N__44903\,
            I => \N__44893\
        );

    \I__10372\ : Span4Mux_v
    port map (
            O => \N__44898\,
            I => \N__44890\
        );

    \I__10371\ : Span4Mux_h
    port map (
            O => \N__44893\,
            I => \N__44887\
        );

    \I__10370\ : Odrv4
    port map (
            O => \N__44890\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__10369\ : Odrv4
    port map (
            O => \N__44887\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__10368\ : InMux
    port map (
            O => \N__44882\,
            I => \N__44879\
        );

    \I__10367\ : LocalMux
    port map (
            O => \N__44879\,
            I => \N__44874\
        );

    \I__10366\ : InMux
    port map (
            O => \N__44878\,
            I => \N__44871\
        );

    \I__10365\ : InMux
    port map (
            O => \N__44877\,
            I => \N__44868\
        );

    \I__10364\ : Span4Mux_h
    port map (
            O => \N__44874\,
            I => \N__44865\
        );

    \I__10363\ : LocalMux
    port map (
            O => \N__44871\,
            I => \N__44862\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__44868\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__10361\ : Odrv4
    port map (
            O => \N__44865\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__10360\ : Odrv12
    port map (
            O => \N__44862\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__10359\ : InMux
    port map (
            O => \N__44855\,
            I => \N__44850\
        );

    \I__10358\ : InMux
    port map (
            O => \N__44854\,
            I => \N__44846\
        );

    \I__10357\ : InMux
    port map (
            O => \N__44853\,
            I => \N__44843\
        );

    \I__10356\ : LocalMux
    port map (
            O => \N__44850\,
            I => \N__44840\
        );

    \I__10355\ : InMux
    port map (
            O => \N__44849\,
            I => \N__44837\
        );

    \I__10354\ : LocalMux
    port map (
            O => \N__44846\,
            I => \N__44834\
        );

    \I__10353\ : LocalMux
    port map (
            O => \N__44843\,
            I => \N__44831\
        );

    \I__10352\ : Span4Mux_v
    port map (
            O => \N__44840\,
            I => \N__44826\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__44837\,
            I => \N__44826\
        );

    \I__10350\ : Span4Mux_v
    port map (
            O => \N__44834\,
            I => \N__44823\
        );

    \I__10349\ : Span4Mux_v
    port map (
            O => \N__44831\,
            I => \N__44818\
        );

    \I__10348\ : Span4Mux_h
    port map (
            O => \N__44826\,
            I => \N__44818\
        );

    \I__10347\ : Odrv4
    port map (
            O => \N__44823\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__10346\ : Odrv4
    port map (
            O => \N__44818\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__10345\ : InMux
    port map (
            O => \N__44813\,
            I => \N__44810\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__44810\,
            I => \N__44806\
        );

    \I__10343\ : InMux
    port map (
            O => \N__44809\,
            I => \N__44802\
        );

    \I__10342\ : Span4Mux_h
    port map (
            O => \N__44806\,
            I => \N__44799\
        );

    \I__10341\ : InMux
    port map (
            O => \N__44805\,
            I => \N__44796\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__44802\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__10339\ : Odrv4
    port map (
            O => \N__44799\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__44796\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__10337\ : InMux
    port map (
            O => \N__44789\,
            I => \N__44784\
        );

    \I__10336\ : InMux
    port map (
            O => \N__44788\,
            I => \N__44781\
        );

    \I__10335\ : InMux
    port map (
            O => \N__44787\,
            I => \N__44778\
        );

    \I__10334\ : LocalMux
    port map (
            O => \N__44784\,
            I => \N__44773\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__44781\,
            I => \N__44773\
        );

    \I__10332\ : LocalMux
    port map (
            O => \N__44778\,
            I => \N__44770\
        );

    \I__10331\ : Span4Mux_h
    port map (
            O => \N__44773\,
            I => \N__44767\
        );

    \I__10330\ : Span4Mux_h
    port map (
            O => \N__44770\,
            I => \N__44763\
        );

    \I__10329\ : Span4Mux_v
    port map (
            O => \N__44767\,
            I => \N__44760\
        );

    \I__10328\ : InMux
    port map (
            O => \N__44766\,
            I => \N__44757\
        );

    \I__10327\ : Odrv4
    port map (
            O => \N__44763\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__10326\ : Odrv4
    port map (
            O => \N__44760\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__44757\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__10324\ : CascadeMux
    port map (
            O => \N__44750\,
            I => \N__44747\
        );

    \I__10323\ : InMux
    port map (
            O => \N__44747\,
            I => \N__44741\
        );

    \I__10322\ : InMux
    port map (
            O => \N__44746\,
            I => \N__44741\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__44741\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__10320\ : CascadeMux
    port map (
            O => \N__44738\,
            I => \N__44735\
        );

    \I__10319\ : InMux
    port map (
            O => \N__44735\,
            I => \N__44730\
        );

    \I__10318\ : InMux
    port map (
            O => \N__44734\,
            I => \N__44727\
        );

    \I__10317\ : CascadeMux
    port map (
            O => \N__44733\,
            I => \N__44724\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__44730\,
            I => \N__44721\
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__44727\,
            I => \N__44718\
        );

    \I__10314\ : InMux
    port map (
            O => \N__44724\,
            I => \N__44715\
        );

    \I__10313\ : Span12Mux_h
    port map (
            O => \N__44721\,
            I => \N__44712\
        );

    \I__10312\ : Span4Mux_h
    port map (
            O => \N__44718\,
            I => \N__44709\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__44715\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10310\ : Odrv12
    port map (
            O => \N__44712\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10309\ : Odrv4
    port map (
            O => \N__44709\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10308\ : InMux
    port map (
            O => \N__44702\,
            I => \N__44699\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__44699\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__10306\ : CascadeMux
    port map (
            O => \N__44696\,
            I => \N__44693\
        );

    \I__10305\ : InMux
    port map (
            O => \N__44693\,
            I => \N__44690\
        );

    \I__10304\ : LocalMux
    port map (
            O => \N__44690\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__10303\ : InMux
    port map (
            O => \N__44687\,
            I => \N__44683\
        );

    \I__10302\ : InMux
    port map (
            O => \N__44686\,
            I => \N__44680\
        );

    \I__10301\ : LocalMux
    port map (
            O => \N__44683\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__44680\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__10299\ : CascadeMux
    port map (
            O => \N__44675\,
            I => \N__44672\
        );

    \I__10298\ : InMux
    port map (
            O => \N__44672\,
            I => \N__44669\
        );

    \I__10297\ : LocalMux
    port map (
            O => \N__44669\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__10296\ : InMux
    port map (
            O => \N__44666\,
            I => \N__44663\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__44663\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__10294\ : CascadeMux
    port map (
            O => \N__44660\,
            I => \N__44657\
        );

    \I__10293\ : InMux
    port map (
            O => \N__44657\,
            I => \N__44654\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__44654\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__10291\ : InMux
    port map (
            O => \N__44651\,
            I => \N__44647\
        );

    \I__10290\ : InMux
    port map (
            O => \N__44650\,
            I => \N__44644\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__44647\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__44644\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__10287\ : InMux
    port map (
            O => \N__44639\,
            I => \N__44636\
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__44636\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__10285\ : InMux
    port map (
            O => \N__44633\,
            I => \N__44628\
        );

    \I__10284\ : CascadeMux
    port map (
            O => \N__44632\,
            I => \N__44624\
        );

    \I__10283\ : InMux
    port map (
            O => \N__44631\,
            I => \N__44621\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__44628\,
            I => \N__44618\
        );

    \I__10281\ : InMux
    port map (
            O => \N__44627\,
            I => \N__44613\
        );

    \I__10280\ : InMux
    port map (
            O => \N__44624\,
            I => \N__44613\
        );

    \I__10279\ : LocalMux
    port map (
            O => \N__44621\,
            I => \N__44606\
        );

    \I__10278\ : Span4Mux_h
    port map (
            O => \N__44618\,
            I => \N__44606\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__44613\,
            I => \N__44606\
        );

    \I__10276\ : Odrv4
    port map (
            O => \N__44606\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__10275\ : IoInMux
    port map (
            O => \N__44603\,
            I => \N__44600\
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__44600\,
            I => \N__44597\
        );

    \I__10273\ : Span4Mux_s1_v
    port map (
            O => \N__44597\,
            I => \N__44594\
        );

    \I__10272\ : Span4Mux_v
    port map (
            O => \N__44594\,
            I => \N__44591\
        );

    \I__10271\ : Span4Mux_v
    port map (
            O => \N__44591\,
            I => \N__44587\
        );

    \I__10270\ : InMux
    port map (
            O => \N__44590\,
            I => \N__44584\
        );

    \I__10269\ : Odrv4
    port map (
            O => \N__44587\,
            I => \T12_c\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__44584\,
            I => \T12_c\
        );

    \I__10267\ : InMux
    port map (
            O => \N__44579\,
            I => \N__44572\
        );

    \I__10266\ : InMux
    port map (
            O => \N__44578\,
            I => \N__44572\
        );

    \I__10265\ : InMux
    port map (
            O => \N__44577\,
            I => \N__44569\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__44572\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__10263\ : LocalMux
    port map (
            O => \N__44569\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__10262\ : InMux
    port map (
            O => \N__44564\,
            I => \N__44560\
        );

    \I__10261\ : InMux
    port map (
            O => \N__44563\,
            I => \N__44557\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__44560\,
            I => \N__44554\
        );

    \I__10259\ : LocalMux
    port map (
            O => \N__44557\,
            I => \N__44551\
        );

    \I__10258\ : Span4Mux_h
    port map (
            O => \N__44554\,
            I => \N__44546\
        );

    \I__10257\ : Span4Mux_v
    port map (
            O => \N__44551\,
            I => \N__44546\
        );

    \I__10256\ : Odrv4
    port map (
            O => \N__44546\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0\
        );

    \I__10255\ : InMux
    port map (
            O => \N__44543\,
            I => \N__44540\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__44540\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__10253\ : InMux
    port map (
            O => \N__44537\,
            I => \N__44534\
        );

    \I__10252\ : LocalMux
    port map (
            O => \N__44534\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__10251\ : CascadeMux
    port map (
            O => \N__44531\,
            I => \N__44528\
        );

    \I__10250\ : InMux
    port map (
            O => \N__44528\,
            I => \N__44525\
        );

    \I__10249\ : LocalMux
    port map (
            O => \N__44525\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__10248\ : InMux
    port map (
            O => \N__44522\,
            I => \N__44519\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__44519\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__10246\ : InMux
    port map (
            O => \N__44516\,
            I => \N__44513\
        );

    \I__10245\ : LocalMux
    port map (
            O => \N__44513\,
            I => \N__44510\
        );

    \I__10244\ : Span4Mux_v
    port map (
            O => \N__44510\,
            I => \N__44506\
        );

    \I__10243\ : InMux
    port map (
            O => \N__44509\,
            I => \N__44503\
        );

    \I__10242\ : Odrv4
    port map (
            O => \N__44506\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__44503\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__10240\ : InMux
    port map (
            O => \N__44498\,
            I => \N__44495\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__44495\,
            I => \N__44492\
        );

    \I__10238\ : Span4Mux_v
    port map (
            O => \N__44492\,
            I => \N__44488\
        );

    \I__10237\ : InMux
    port map (
            O => \N__44491\,
            I => \N__44485\
        );

    \I__10236\ : Odrv4
    port map (
            O => \N__44488\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__44485\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__10234\ : CascadeMux
    port map (
            O => \N__44480\,
            I => \N__44477\
        );

    \I__10233\ : InMux
    port map (
            O => \N__44477\,
            I => \N__44473\
        );

    \I__10232\ : CascadeMux
    port map (
            O => \N__44476\,
            I => \N__44470\
        );

    \I__10231\ : LocalMux
    port map (
            O => \N__44473\,
            I => \N__44467\
        );

    \I__10230\ : InMux
    port map (
            O => \N__44470\,
            I => \N__44464\
        );

    \I__10229\ : Odrv4
    port map (
            O => \N__44467\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__44464\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__10227\ : InMux
    port map (
            O => \N__44459\,
            I => \N__44456\
        );

    \I__10226\ : LocalMux
    port map (
            O => \N__44456\,
            I => \N__44452\
        );

    \I__10225\ : InMux
    port map (
            O => \N__44455\,
            I => \N__44449\
        );

    \I__10224\ : Odrv4
    port map (
            O => \N__44452\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__10223\ : LocalMux
    port map (
            O => \N__44449\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__10222\ : InMux
    port map (
            O => \N__44444\,
            I => \N__44441\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__44441\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__10220\ : InMux
    port map (
            O => \N__44438\,
            I => \N__44435\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__44435\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__10218\ : CascadeMux
    port map (
            O => \N__44432\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_\
        );

    \I__10217\ : InMux
    port map (
            O => \N__44429\,
            I => \N__44426\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__44426\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__10215\ : InMux
    port map (
            O => \N__44423\,
            I => \N__44420\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__44420\,
            I => \N__44416\
        );

    \I__10213\ : InMux
    port map (
            O => \N__44419\,
            I => \N__44413\
        );

    \I__10212\ : Span12Mux_v
    port map (
            O => \N__44416\,
            I => \N__44408\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__44413\,
            I => \N__44408\
        );

    \I__10210\ : Span12Mux_h
    port map (
            O => \N__44408\,
            I => \N__44405\
        );

    \I__10209\ : Odrv12
    port map (
            O => \N__44405\,
            I => \pwm_generator_inst.O_10\
        );

    \I__10208\ : CascadeMux
    port map (
            O => \N__44402\,
            I => \N__44399\
        );

    \I__10207\ : InMux
    port map (
            O => \N__44399\,
            I => \N__44396\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__44396\,
            I => \N__44391\
        );

    \I__10205\ : InMux
    port map (
            O => \N__44395\,
            I => \N__44388\
        );

    \I__10204\ : InMux
    port map (
            O => \N__44394\,
            I => \N__44385\
        );

    \I__10203\ : Span4Mux_h
    port map (
            O => \N__44391\,
            I => \N__44382\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__44388\,
            I => \N__44379\
        );

    \I__10201\ : LocalMux
    port map (
            O => \N__44385\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__10200\ : Odrv4
    port map (
            O => \N__44382\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__10199\ : Odrv4
    port map (
            O => \N__44379\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__10198\ : InMux
    port map (
            O => \N__44372\,
            I => \N__44368\
        );

    \I__10197\ : InMux
    port map (
            O => \N__44371\,
            I => \N__44364\
        );

    \I__10196\ : LocalMux
    port map (
            O => \N__44368\,
            I => \N__44361\
        );

    \I__10195\ : InMux
    port map (
            O => \N__44367\,
            I => \N__44358\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__44364\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__10193\ : Odrv4
    port map (
            O => \N__44361\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__44358\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__10191\ : InMux
    port map (
            O => \N__44351\,
            I => \N__44346\
        );

    \I__10190\ : InMux
    port map (
            O => \N__44350\,
            I => \N__44342\
        );

    \I__10189\ : InMux
    port map (
            O => \N__44349\,
            I => \N__44339\
        );

    \I__10188\ : LocalMux
    port map (
            O => \N__44346\,
            I => \N__44336\
        );

    \I__10187\ : InMux
    port map (
            O => \N__44345\,
            I => \N__44333\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__44342\,
            I => \N__44330\
        );

    \I__10185\ : LocalMux
    port map (
            O => \N__44339\,
            I => \N__44327\
        );

    \I__10184\ : Span4Mux_h
    port map (
            O => \N__44336\,
            I => \N__44324\
        );

    \I__10183\ : LocalMux
    port map (
            O => \N__44333\,
            I => \N__44321\
        );

    \I__10182\ : Span12Mux_s7_v
    port map (
            O => \N__44330\,
            I => \N__44318\
        );

    \I__10181\ : Span12Mux_v
    port map (
            O => \N__44327\,
            I => \N__44315\
        );

    \I__10180\ : Span4Mux_v
    port map (
            O => \N__44324\,
            I => \N__44310\
        );

    \I__10179\ : Span4Mux_h
    port map (
            O => \N__44321\,
            I => \N__44310\
        );

    \I__10178\ : Odrv12
    port map (
            O => \N__44318\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__10177\ : Odrv12
    port map (
            O => \N__44315\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__10176\ : Odrv4
    port map (
            O => \N__44310\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__10175\ : InMux
    port map (
            O => \N__44303\,
            I => \N__44299\
        );

    \I__10174\ : InMux
    port map (
            O => \N__44302\,
            I => \N__44294\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__44299\,
            I => \N__44291\
        );

    \I__10172\ : InMux
    port map (
            O => \N__44298\,
            I => \N__44288\
        );

    \I__10171\ : InMux
    port map (
            O => \N__44297\,
            I => \N__44285\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__44294\,
            I => \N__44282\
        );

    \I__10169\ : Span4Mux_v
    port map (
            O => \N__44291\,
            I => \N__44279\
        );

    \I__10168\ : LocalMux
    port map (
            O => \N__44288\,
            I => \N__44276\
        );

    \I__10167\ : LocalMux
    port map (
            O => \N__44285\,
            I => \N__44273\
        );

    \I__10166\ : Span4Mux_v
    port map (
            O => \N__44282\,
            I => \N__44268\
        );

    \I__10165\ : Span4Mux_h
    port map (
            O => \N__44279\,
            I => \N__44268\
        );

    \I__10164\ : Span4Mux_v
    port map (
            O => \N__44276\,
            I => \N__44263\
        );

    \I__10163\ : Span4Mux_h
    port map (
            O => \N__44273\,
            I => \N__44263\
        );

    \I__10162\ : Odrv4
    port map (
            O => \N__44268\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__10161\ : Odrv4
    port map (
            O => \N__44263\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__10160\ : InMux
    port map (
            O => \N__44258\,
            I => \N__44254\
        );

    \I__10159\ : InMux
    port map (
            O => \N__44257\,
            I => \N__44250\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__44254\,
            I => \N__44247\
        );

    \I__10157\ : InMux
    port map (
            O => \N__44253\,
            I => \N__44244\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__44250\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__10155\ : Odrv4
    port map (
            O => \N__44247\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__44244\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__10153\ : CascadeMux
    port map (
            O => \N__44237\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\
        );

    \I__10152\ : InMux
    port map (
            O => \N__44234\,
            I => \N__44226\
        );

    \I__10151\ : InMux
    port map (
            O => \N__44233\,
            I => \N__44226\
        );

    \I__10150\ : InMux
    port map (
            O => \N__44232\,
            I => \N__44223\
        );

    \I__10149\ : InMux
    port map (
            O => \N__44231\,
            I => \N__44220\
        );

    \I__10148\ : LocalMux
    port map (
            O => \N__44226\,
            I => \N__44217\
        );

    \I__10147\ : LocalMux
    port map (
            O => \N__44223\,
            I => \N__44214\
        );

    \I__10146\ : LocalMux
    port map (
            O => \N__44220\,
            I => \N__44211\
        );

    \I__10145\ : Span4Mux_h
    port map (
            O => \N__44217\,
            I => \N__44208\
        );

    \I__10144\ : Span4Mux_h
    port map (
            O => \N__44214\,
            I => \N__44203\
        );

    \I__10143\ : Span4Mux_v
    port map (
            O => \N__44211\,
            I => \N__44203\
        );

    \I__10142\ : Odrv4
    port map (
            O => \N__44208\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__10141\ : Odrv4
    port map (
            O => \N__44203\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__10140\ : InMux
    port map (
            O => \N__44198\,
            I => \N__44193\
        );

    \I__10139\ : InMux
    port map (
            O => \N__44197\,
            I => \N__44188\
        );

    \I__10138\ : InMux
    port map (
            O => \N__44196\,
            I => \N__44188\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__44193\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__44188\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__10135\ : CascadeMux
    port map (
            O => \N__44183\,
            I => \N__44180\
        );

    \I__10134\ : InMux
    port map (
            O => \N__44180\,
            I => \N__44174\
        );

    \I__10133\ : InMux
    port map (
            O => \N__44179\,
            I => \N__44174\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__44174\,
            I => \N__44171\
        );

    \I__10131\ : Span4Mux_h
    port map (
            O => \N__44171\,
            I => \N__44168\
        );

    \I__10130\ : Odrv4
    port map (
            O => \N__44168\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\
        );

    \I__10129\ : CascadeMux
    port map (
            O => \N__44165\,
            I => \N__44160\
        );

    \I__10128\ : InMux
    port map (
            O => \N__44164\,
            I => \N__44157\
        );

    \I__10127\ : InMux
    port map (
            O => \N__44163\,
            I => \N__44152\
        );

    \I__10126\ : InMux
    port map (
            O => \N__44160\,
            I => \N__44152\
        );

    \I__10125\ : LocalMux
    port map (
            O => \N__44157\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__10124\ : LocalMux
    port map (
            O => \N__44152\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44147\,
            I => \N__44141\
        );

    \I__10122\ : InMux
    port map (
            O => \N__44146\,
            I => \N__44141\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__44141\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\
        );

    \I__10120\ : CascadeMux
    port map (
            O => \N__44138\,
            I => \N__44133\
        );

    \I__10119\ : InMux
    port map (
            O => \N__44137\,
            I => \N__44126\
        );

    \I__10118\ : InMux
    port map (
            O => \N__44136\,
            I => \N__44126\
        );

    \I__10117\ : InMux
    port map (
            O => \N__44133\,
            I => \N__44126\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__44126\,
            I => \N__44123\
        );

    \I__10115\ : Span4Mux_h
    port map (
            O => \N__44123\,
            I => \N__44120\
        );

    \I__10114\ : Odrv4
    port map (
            O => \N__44120\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\
        );

    \I__10113\ : CEMux
    port map (
            O => \N__44117\,
            I => \N__44113\
        );

    \I__10112\ : CEMux
    port map (
            O => \N__44116\,
            I => \N__44109\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__44113\,
            I => \N__44105\
        );

    \I__10110\ : CEMux
    port map (
            O => \N__44112\,
            I => \N__44102\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__44109\,
            I => \N__44099\
        );

    \I__10108\ : CEMux
    port map (
            O => \N__44108\,
            I => \N__44096\
        );

    \I__10107\ : Span4Mux_h
    port map (
            O => \N__44105\,
            I => \N__44092\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__44102\,
            I => \N__44089\
        );

    \I__10105\ : Span4Mux_v
    port map (
            O => \N__44099\,
            I => \N__44086\
        );

    \I__10104\ : LocalMux
    port map (
            O => \N__44096\,
            I => \N__44083\
        );

    \I__10103\ : CEMux
    port map (
            O => \N__44095\,
            I => \N__44080\
        );

    \I__10102\ : Span4Mux_v
    port map (
            O => \N__44092\,
            I => \N__44075\
        );

    \I__10101\ : Span4Mux_h
    port map (
            O => \N__44089\,
            I => \N__44075\
        );

    \I__10100\ : Span4Mux_h
    port map (
            O => \N__44086\,
            I => \N__44072\
        );

    \I__10099\ : Span4Mux_h
    port map (
            O => \N__44083\,
            I => \N__44069\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__44080\,
            I => \N__44066\
        );

    \I__10097\ : Odrv4
    port map (
            O => \N__44075\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__10096\ : Odrv4
    port map (
            O => \N__44072\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__10095\ : Odrv4
    port map (
            O => \N__44069\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__10094\ : Odrv12
    port map (
            O => \N__44066\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__10093\ : InMux
    port map (
            O => \N__44057\,
            I => \N__44052\
        );

    \I__10092\ : InMux
    port map (
            O => \N__44056\,
            I => \N__44049\
        );

    \I__10091\ : CascadeMux
    port map (
            O => \N__44055\,
            I => \N__44046\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__44052\,
            I => \N__44043\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__44049\,
            I => \N__44039\
        );

    \I__10088\ : InMux
    port map (
            O => \N__44046\,
            I => \N__44036\
        );

    \I__10087\ : Span12Mux_v
    port map (
            O => \N__44043\,
            I => \N__44033\
        );

    \I__10086\ : InMux
    port map (
            O => \N__44042\,
            I => \N__44030\
        );

    \I__10085\ : Span12Mux_s11_v
    port map (
            O => \N__44039\,
            I => \N__44027\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__44036\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__10083\ : Odrv12
    port map (
            O => \N__44033\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__10082\ : LocalMux
    port map (
            O => \N__44030\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__10081\ : Odrv12
    port map (
            O => \N__44027\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__10080\ : InMux
    port map (
            O => \N__44018\,
            I => \N__44013\
        );

    \I__10079\ : InMux
    port map (
            O => \N__44017\,
            I => \N__44010\
        );

    \I__10078\ : InMux
    port map (
            O => \N__44016\,
            I => \N__44007\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__44013\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__10076\ : LocalMux
    port map (
            O => \N__44010\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__44007\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__10074\ : InMux
    port map (
            O => \N__44000\,
            I => \N__43996\
        );

    \I__10073\ : InMux
    port map (
            O => \N__43999\,
            I => \N__43992\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__43996\,
            I => \N__43989\
        );

    \I__10071\ : InMux
    port map (
            O => \N__43995\,
            I => \N__43986\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__43992\,
            I => \N__43978\
        );

    \I__10069\ : Span4Mux_v
    port map (
            O => \N__43989\,
            I => \N__43978\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__43986\,
            I => \N__43978\
        );

    \I__10067\ : InMux
    port map (
            O => \N__43985\,
            I => \N__43975\
        );

    \I__10066\ : Odrv4
    port map (
            O => \N__43978\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__43975\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__10064\ : InMux
    port map (
            O => \N__43970\,
            I => \N__43967\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__43967\,
            I => \N__43961\
        );

    \I__10062\ : InMux
    port map (
            O => \N__43966\,
            I => \N__43958\
        );

    \I__10061\ : InMux
    port map (
            O => \N__43965\,
            I => \N__43955\
        );

    \I__10060\ : InMux
    port map (
            O => \N__43964\,
            I => \N__43952\
        );

    \I__10059\ : Span4Mux_v
    port map (
            O => \N__43961\,
            I => \N__43949\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__43958\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__43955\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__43952\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__10055\ : Odrv4
    port map (
            O => \N__43949\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__10054\ : CEMux
    port map (
            O => \N__43940\,
            I => \N__43935\
        );

    \I__10053\ : CEMux
    port map (
            O => \N__43939\,
            I => \N__43931\
        );

    \I__10052\ : CEMux
    port map (
            O => \N__43938\,
            I => \N__43928\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__43935\,
            I => \N__43925\
        );

    \I__10050\ : CEMux
    port map (
            O => \N__43934\,
            I => \N__43922\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__43931\,
            I => \N__43919\
        );

    \I__10048\ : LocalMux
    port map (
            O => \N__43928\,
            I => \N__43916\
        );

    \I__10047\ : Span4Mux_v
    port map (
            O => \N__43925\,
            I => \N__43911\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__43922\,
            I => \N__43911\
        );

    \I__10045\ : Span4Mux_h
    port map (
            O => \N__43919\,
            I => \N__43908\
        );

    \I__10044\ : Span4Mux_h
    port map (
            O => \N__43916\,
            I => \N__43905\
        );

    \I__10043\ : Span4Mux_h
    port map (
            O => \N__43911\,
            I => \N__43902\
        );

    \I__10042\ : Odrv4
    port map (
            O => \N__43908\,
            I => \delay_measurement_inst.delay_tr_timer.N_201_i\
        );

    \I__10041\ : Odrv4
    port map (
            O => \N__43905\,
            I => \delay_measurement_inst.delay_tr_timer.N_201_i\
        );

    \I__10040\ : Odrv4
    port map (
            O => \N__43902\,
            I => \delay_measurement_inst.delay_tr_timer.N_201_i\
        );

    \I__10039\ : InMux
    port map (
            O => \N__43895\,
            I => \bfn_17_14_0_\
        );

    \I__10038\ : InMux
    port map (
            O => \N__43892\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__10037\ : InMux
    port map (
            O => \N__43889\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__10036\ : InMux
    port map (
            O => \N__43886\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__10035\ : InMux
    port map (
            O => \N__43883\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__10034\ : InMux
    port map (
            O => \N__43880\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__10033\ : InMux
    port map (
            O => \N__43877\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__10032\ : InMux
    port map (
            O => \N__43874\,
            I => \N__43870\
        );

    \I__10031\ : InMux
    port map (
            O => \N__43873\,
            I => \N__43865\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__43870\,
            I => \N__43862\
        );

    \I__10029\ : InMux
    port map (
            O => \N__43869\,
            I => \N__43859\
        );

    \I__10028\ : InMux
    port map (
            O => \N__43868\,
            I => \N__43856\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__43865\,
            I => \N__43853\
        );

    \I__10026\ : Span4Mux_h
    port map (
            O => \N__43862\,
            I => \N__43848\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__43859\,
            I => \N__43848\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__43856\,
            I => \N__43845\
        );

    \I__10023\ : Span4Mux_h
    port map (
            O => \N__43853\,
            I => \N__43842\
        );

    \I__10022\ : Span4Mux_v
    port map (
            O => \N__43848\,
            I => \N__43839\
        );

    \I__10021\ : Odrv12
    port map (
            O => \N__43845\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__10020\ : Odrv4
    port map (
            O => \N__43842\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__10019\ : Odrv4
    port map (
            O => \N__43839\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__10018\ : InMux
    port map (
            O => \N__43832\,
            I => \N__43829\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__43829\,
            I => \N__43825\
        );

    \I__10016\ : InMux
    port map (
            O => \N__43828\,
            I => \N__43821\
        );

    \I__10015\ : Span4Mux_v
    port map (
            O => \N__43825\,
            I => \N__43818\
        );

    \I__10014\ : InMux
    port map (
            O => \N__43824\,
            I => \N__43815\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__43821\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__10012\ : Odrv4
    port map (
            O => \N__43818\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__43815\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__10010\ : InMux
    port map (
            O => \N__43808\,
            I => \N__43805\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__43805\,
            I => \N__43802\
        );

    \I__10008\ : Span4Mux_v
    port map (
            O => \N__43802\,
            I => \N__43798\
        );

    \I__10007\ : InMux
    port map (
            O => \N__43801\,
            I => \N__43795\
        );

    \I__10006\ : Odrv4
    port map (
            O => \N__43798\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__43795\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__10004\ : InMux
    port map (
            O => \N__43790\,
            I => \N__43785\
        );

    \I__10003\ : InMux
    port map (
            O => \N__43789\,
            I => \N__43780\
        );

    \I__10002\ : InMux
    port map (
            O => \N__43788\,
            I => \N__43780\
        );

    \I__10001\ : LocalMux
    port map (
            O => \N__43785\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__10000\ : LocalMux
    port map (
            O => \N__43780\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__9999\ : InMux
    port map (
            O => \N__43775\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__9998\ : CascadeMux
    port map (
            O => \N__43772\,
            I => \N__43767\
        );

    \I__9997\ : CascadeMux
    port map (
            O => \N__43771\,
            I => \N__43764\
        );

    \I__9996\ : InMux
    port map (
            O => \N__43770\,
            I => \N__43761\
        );

    \I__9995\ : InMux
    port map (
            O => \N__43767\,
            I => \N__43756\
        );

    \I__9994\ : InMux
    port map (
            O => \N__43764\,
            I => \N__43756\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__43761\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__43756\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9991\ : InMux
    port map (
            O => \N__43751\,
            I => \bfn_17_13_0_\
        );

    \I__9990\ : InMux
    port map (
            O => \N__43748\,
            I => \N__43741\
        );

    \I__9989\ : InMux
    port map (
            O => \N__43747\,
            I => \N__43741\
        );

    \I__9988\ : InMux
    port map (
            O => \N__43746\,
            I => \N__43738\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__43741\,
            I => \N__43735\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__43738\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9985\ : Odrv12
    port map (
            O => \N__43735\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9984\ : InMux
    port map (
            O => \N__43730\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__9983\ : CascadeMux
    port map (
            O => \N__43727\,
            I => \N__43724\
        );

    \I__9982\ : InMux
    port map (
            O => \N__43724\,
            I => \N__43717\
        );

    \I__9981\ : InMux
    port map (
            O => \N__43723\,
            I => \N__43717\
        );

    \I__9980\ : InMux
    port map (
            O => \N__43722\,
            I => \N__43714\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__43717\,
            I => \N__43711\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__43714\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9977\ : Odrv12
    port map (
            O => \N__43711\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9976\ : InMux
    port map (
            O => \N__43706\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__9975\ : InMux
    port map (
            O => \N__43703\,
            I => \N__43696\
        );

    \I__9974\ : InMux
    port map (
            O => \N__43702\,
            I => \N__43696\
        );

    \I__9973\ : InMux
    port map (
            O => \N__43701\,
            I => \N__43693\
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__43696\,
            I => \N__43690\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__43693\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__9970\ : Odrv4
    port map (
            O => \N__43690\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__9969\ : InMux
    port map (
            O => \N__43685\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__9968\ : CascadeMux
    port map (
            O => \N__43682\,
            I => \N__43678\
        );

    \I__9967\ : InMux
    port map (
            O => \N__43681\,
            I => \N__43672\
        );

    \I__9966\ : InMux
    port map (
            O => \N__43678\,
            I => \N__43672\
        );

    \I__9965\ : InMux
    port map (
            O => \N__43677\,
            I => \N__43669\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__43672\,
            I => \N__43666\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__43669\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__9962\ : Odrv4
    port map (
            O => \N__43666\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__9961\ : InMux
    port map (
            O => \N__43661\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__9960\ : InMux
    port map (
            O => \N__43658\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__9959\ : InMux
    port map (
            O => \N__43655\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__9958\ : InMux
    port map (
            O => \N__43652\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__9957\ : InMux
    port map (
            O => \N__43649\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__9956\ : InMux
    port map (
            O => \N__43646\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__9955\ : InMux
    port map (
            O => \N__43643\,
            I => \bfn_17_12_0_\
        );

    \I__9954\ : InMux
    port map (
            O => \N__43640\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__9953\ : InMux
    port map (
            O => \N__43637\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__9952\ : InMux
    port map (
            O => \N__43634\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__9951\ : InMux
    port map (
            O => \N__43631\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__9950\ : InMux
    port map (
            O => \N__43628\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__9949\ : InMux
    port map (
            O => \N__43625\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__9948\ : InMux
    port map (
            O => \N__43622\,
            I => \N__43619\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__43619\,
            I => \N__43614\
        );

    \I__9946\ : InMux
    port map (
            O => \N__43618\,
            I => \N__43611\
        );

    \I__9945\ : InMux
    port map (
            O => \N__43617\,
            I => \N__43608\
        );

    \I__9944\ : Span4Mux_v
    port map (
            O => \N__43614\,
            I => \N__43605\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__43611\,
            I => \N__43600\
        );

    \I__9942\ : LocalMux
    port map (
            O => \N__43608\,
            I => \N__43600\
        );

    \I__9941\ : Span4Mux_h
    port map (
            O => \N__43605\,
            I => \N__43597\
        );

    \I__9940\ : Odrv12
    port map (
            O => \N__43600\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__9939\ : Odrv4
    port map (
            O => \N__43597\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__9938\ : InMux
    port map (
            O => \N__43592\,
            I => \N__43589\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__43589\,
            I => \N__43585\
        );

    \I__9936\ : InMux
    port map (
            O => \N__43588\,
            I => \N__43582\
        );

    \I__9935\ : Span4Mux_v
    port map (
            O => \N__43585\,
            I => \N__43575\
        );

    \I__9934\ : LocalMux
    port map (
            O => \N__43582\,
            I => \N__43575\
        );

    \I__9933\ : InMux
    port map (
            O => \N__43581\,
            I => \N__43570\
        );

    \I__9932\ : InMux
    port map (
            O => \N__43580\,
            I => \N__43570\
        );

    \I__9931\ : Odrv4
    port map (
            O => \N__43575\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__43570\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__9929\ : InMux
    port map (
            O => \N__43565\,
            I => \N__43561\
        );

    \I__9928\ : InMux
    port map (
            O => \N__43564\,
            I => \N__43556\
        );

    \I__9927\ : LocalMux
    port map (
            O => \N__43561\,
            I => \N__43553\
        );

    \I__9926\ : InMux
    port map (
            O => \N__43560\,
            I => \N__43550\
        );

    \I__9925\ : CascadeMux
    port map (
            O => \N__43559\,
            I => \N__43547\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__43556\,
            I => \N__43544\
        );

    \I__9923\ : Span4Mux_v
    port map (
            O => \N__43553\,
            I => \N__43539\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__43550\,
            I => \N__43539\
        );

    \I__9921\ : InMux
    port map (
            O => \N__43547\,
            I => \N__43536\
        );

    \I__9920\ : Span4Mux_h
    port map (
            O => \N__43544\,
            I => \N__43533\
        );

    \I__9919\ : Span4Mux_v
    port map (
            O => \N__43539\,
            I => \N__43530\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__43536\,
            I => \N__43527\
        );

    \I__9917\ : Odrv4
    port map (
            O => \N__43533\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__9916\ : Odrv4
    port map (
            O => \N__43530\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__9915\ : Odrv12
    port map (
            O => \N__43527\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__9914\ : InMux
    port map (
            O => \N__43520\,
            I => \N__43515\
        );

    \I__9913\ : InMux
    port map (
            O => \N__43519\,
            I => \N__43512\
        );

    \I__9912\ : InMux
    port map (
            O => \N__43518\,
            I => \N__43509\
        );

    \I__9911\ : LocalMux
    port map (
            O => \N__43515\,
            I => \N__43506\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__43512\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__43509\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__9908\ : Odrv4
    port map (
            O => \N__43506\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__9907\ : InMux
    port map (
            O => \N__43499\,
            I => \N__43494\
        );

    \I__9906\ : InMux
    port map (
            O => \N__43498\,
            I => \N__43491\
        );

    \I__9905\ : InMux
    port map (
            O => \N__43497\,
            I => \N__43488\
        );

    \I__9904\ : LocalMux
    port map (
            O => \N__43494\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__9903\ : LocalMux
    port map (
            O => \N__43491\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__43488\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__9901\ : InMux
    port map (
            O => \N__43481\,
            I => \N__43477\
        );

    \I__9900\ : InMux
    port map (
            O => \N__43480\,
            I => \N__43474\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__43477\,
            I => \N__43469\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__43474\,
            I => \N__43466\
        );

    \I__9897\ : InMux
    port map (
            O => \N__43473\,
            I => \N__43463\
        );

    \I__9896\ : InMux
    port map (
            O => \N__43472\,
            I => \N__43460\
        );

    \I__9895\ : Span4Mux_h
    port map (
            O => \N__43469\,
            I => \N__43457\
        );

    \I__9894\ : Span4Mux_v
    port map (
            O => \N__43466\,
            I => \N__43454\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__43463\,
            I => \N__43449\
        );

    \I__9892\ : LocalMux
    port map (
            O => \N__43460\,
            I => \N__43449\
        );

    \I__9891\ : Odrv4
    port map (
            O => \N__43457\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__9890\ : Odrv4
    port map (
            O => \N__43454\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__9889\ : Odrv12
    port map (
            O => \N__43449\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__9888\ : InMux
    port map (
            O => \N__43442\,
            I => \N__43439\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__43439\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\
        );

    \I__9886\ : InMux
    port map (
            O => \N__43436\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__9885\ : CascadeMux
    port map (
            O => \N__43433\,
            I => \N__43430\
        );

    \I__9884\ : InMux
    port map (
            O => \N__43430\,
            I => \N__43427\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__43427\,
            I => \N__43424\
        );

    \I__9882\ : Odrv4
    port map (
            O => \N__43424\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28\
        );

    \I__9881\ : InMux
    port map (
            O => \N__43421\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__9880\ : InMux
    port map (
            O => \N__43418\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__9879\ : InMux
    port map (
            O => \N__43415\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__9878\ : InMux
    port map (
            O => \N__43412\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__9877\ : InMux
    port map (
            O => \N__43409\,
            I => \N__43406\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__43406\,
            I => \N__43402\
        );

    \I__9875\ : InMux
    port map (
            O => \N__43405\,
            I => \N__43398\
        );

    \I__9874\ : Span4Mux_h
    port map (
            O => \N__43402\,
            I => \N__43395\
        );

    \I__9873\ : InMux
    port map (
            O => \N__43401\,
            I => \N__43392\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__43398\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__9871\ : Odrv4
    port map (
            O => \N__43395\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__43392\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__9869\ : InMux
    port map (
            O => \N__43385\,
            I => \N__43380\
        );

    \I__9868\ : InMux
    port map (
            O => \N__43384\,
            I => \N__43377\
        );

    \I__9867\ : InMux
    port map (
            O => \N__43383\,
            I => \N__43374\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__43380\,
            I => \N__43371\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__43377\,
            I => \N__43368\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__43374\,
            I => \N__43365\
        );

    \I__9863\ : Span4Mux_h
    port map (
            O => \N__43371\,
            I => \N__43362\
        );

    \I__9862\ : Span4Mux_h
    port map (
            O => \N__43368\,
            I => \N__43359\
        );

    \I__9861\ : Span4Mux_v
    port map (
            O => \N__43365\,
            I => \N__43355\
        );

    \I__9860\ : Span4Mux_v
    port map (
            O => \N__43362\,
            I => \N__43352\
        );

    \I__9859\ : Span4Mux_v
    port map (
            O => \N__43359\,
            I => \N__43349\
        );

    \I__9858\ : InMux
    port map (
            O => \N__43358\,
            I => \N__43346\
        );

    \I__9857\ : Odrv4
    port map (
            O => \N__43355\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__9856\ : Odrv4
    port map (
            O => \N__43352\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__9855\ : Odrv4
    port map (
            O => \N__43349\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__9854\ : LocalMux
    port map (
            O => \N__43346\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__9853\ : InMux
    port map (
            O => \N__43337\,
            I => \N__43334\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__43334\,
            I => \N__43330\
        );

    \I__9851\ : InMux
    port map (
            O => \N__43333\,
            I => \N__43327\
        );

    \I__9850\ : Odrv4
    port map (
            O => \N__43330\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__9849\ : LocalMux
    port map (
            O => \N__43327\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__9848\ : CascadeMux
    port map (
            O => \N__43322\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\
        );

    \I__9847\ : InMux
    port map (
            O => \N__43319\,
            I => \N__43312\
        );

    \I__9846\ : InMux
    port map (
            O => \N__43318\,
            I => \N__43312\
        );

    \I__9845\ : InMux
    port map (
            O => \N__43317\,
            I => \N__43309\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__43312\,
            I => \N__43306\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__43309\,
            I => \N__43303\
        );

    \I__9842\ : Span4Mux_h
    port map (
            O => \N__43306\,
            I => \N__43300\
        );

    \I__9841\ : Span12Mux_v
    port map (
            O => \N__43303\,
            I => \N__43296\
        );

    \I__9840\ : Span4Mux_v
    port map (
            O => \N__43300\,
            I => \N__43293\
        );

    \I__9839\ : InMux
    port map (
            O => \N__43299\,
            I => \N__43290\
        );

    \I__9838\ : Odrv12
    port map (
            O => \N__43296\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__9837\ : Odrv4
    port map (
            O => \N__43293\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__9836\ : LocalMux
    port map (
            O => \N__43290\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__9835\ : InMux
    port map (
            O => \N__43283\,
            I => \N__43277\
        );

    \I__9834\ : InMux
    port map (
            O => \N__43282\,
            I => \N__43277\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__43277\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__9832\ : InMux
    port map (
            O => \N__43274\,
            I => \N__43269\
        );

    \I__9831\ : InMux
    port map (
            O => \N__43273\,
            I => \N__43266\
        );

    \I__9830\ : InMux
    port map (
            O => \N__43272\,
            I => \N__43263\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__43269\,
            I => \N__43260\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__43266\,
            I => \N__43257\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__43263\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__9826\ : Odrv4
    port map (
            O => \N__43260\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__9825\ : Odrv4
    port map (
            O => \N__43257\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__9824\ : InMux
    port map (
            O => \N__43250\,
            I => \N__43246\
        );

    \I__9823\ : InMux
    port map (
            O => \N__43249\,
            I => \N__43242\
        );

    \I__9822\ : LocalMux
    port map (
            O => \N__43246\,
            I => \N__43239\
        );

    \I__9821\ : InMux
    port map (
            O => \N__43245\,
            I => \N__43236\
        );

    \I__9820\ : LocalMux
    port map (
            O => \N__43242\,
            I => \N__43233\
        );

    \I__9819\ : Span4Mux_h
    port map (
            O => \N__43239\,
            I => \N__43229\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__43236\,
            I => \N__43224\
        );

    \I__9817\ : Span4Mux_h
    port map (
            O => \N__43233\,
            I => \N__43224\
        );

    \I__9816\ : CascadeMux
    port map (
            O => \N__43232\,
            I => \N__43221\
        );

    \I__9815\ : Span4Mux_v
    port map (
            O => \N__43229\,
            I => \N__43218\
        );

    \I__9814\ : Span4Mux_v
    port map (
            O => \N__43224\,
            I => \N__43215\
        );

    \I__9813\ : InMux
    port map (
            O => \N__43221\,
            I => \N__43212\
        );

    \I__9812\ : Odrv4
    port map (
            O => \N__43218\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__9811\ : Odrv4
    port map (
            O => \N__43215\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__43212\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__9809\ : InMux
    port map (
            O => \N__43205\,
            I => \N__43199\
        );

    \I__9808\ : InMux
    port map (
            O => \N__43204\,
            I => \N__43199\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__43199\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\
        );

    \I__9806\ : CascadeMux
    port map (
            O => \N__43196\,
            I => \N__43193\
        );

    \I__9805\ : InMux
    port map (
            O => \N__43193\,
            I => \N__43187\
        );

    \I__9804\ : InMux
    port map (
            O => \N__43192\,
            I => \N__43187\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__43187\,
            I => \N__43184\
        );

    \I__9802\ : Span4Mux_v
    port map (
            O => \N__43184\,
            I => \N__43181\
        );

    \I__9801\ : Odrv4
    port map (
            O => \N__43181\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\
        );

    \I__9800\ : InMux
    port map (
            O => \N__43178\,
            I => \N__43174\
        );

    \I__9799\ : InMux
    port map (
            O => \N__43177\,
            I => \N__43170\
        );

    \I__9798\ : LocalMux
    port map (
            O => \N__43174\,
            I => \N__43167\
        );

    \I__9797\ : InMux
    port map (
            O => \N__43173\,
            I => \N__43164\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__43170\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__9795\ : Odrv4
    port map (
            O => \N__43167\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__9794\ : LocalMux
    port map (
            O => \N__43164\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__9793\ : InMux
    port map (
            O => \N__43157\,
            I => \N__43152\
        );

    \I__9792\ : InMux
    port map (
            O => \N__43156\,
            I => \N__43149\
        );

    \I__9791\ : InMux
    port map (
            O => \N__43155\,
            I => \N__43146\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__43152\,
            I => \N__43142\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__43149\,
            I => \N__43139\
        );

    \I__9788\ : LocalMux
    port map (
            O => \N__43146\,
            I => \N__43136\
        );

    \I__9787\ : InMux
    port map (
            O => \N__43145\,
            I => \N__43133\
        );

    \I__9786\ : Odrv4
    port map (
            O => \N__43142\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__9785\ : Odrv4
    port map (
            O => \N__43139\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__9784\ : Odrv4
    port map (
            O => \N__43136\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__43133\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__9782\ : InMux
    port map (
            O => \N__43124\,
            I => \N__43118\
        );

    \I__9781\ : InMux
    port map (
            O => \N__43123\,
            I => \N__43118\
        );

    \I__9780\ : LocalMux
    port map (
            O => \N__43118\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__9779\ : CascadeMux
    port map (
            O => \N__43115\,
            I => \N__43112\
        );

    \I__9778\ : InMux
    port map (
            O => \N__43112\,
            I => \N__43106\
        );

    \I__9777\ : InMux
    port map (
            O => \N__43111\,
            I => \N__43106\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__43106\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__9775\ : CascadeMux
    port map (
            O => \N__43103\,
            I => \N__43100\
        );

    \I__9774\ : InMux
    port map (
            O => \N__43100\,
            I => \N__43097\
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__43097\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__9772\ : CascadeMux
    port map (
            O => \N__43094\,
            I => \N__43090\
        );

    \I__9771\ : InMux
    port map (
            O => \N__43093\,
            I => \N__43087\
        );

    \I__9770\ : InMux
    port map (
            O => \N__43090\,
            I => \N__43084\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__43087\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__43084\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__9767\ : InMux
    port map (
            O => \N__43079\,
            I => \N__43076\
        );

    \I__9766\ : LocalMux
    port map (
            O => \N__43076\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\
        );

    \I__9765\ : InMux
    port map (
            O => \N__43073\,
            I => \N__43070\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__43070\,
            I => \N__43064\
        );

    \I__9763\ : InMux
    port map (
            O => \N__43069\,
            I => \N__43061\
        );

    \I__9762\ : InMux
    port map (
            O => \N__43068\,
            I => \N__43058\
        );

    \I__9761\ : InMux
    port map (
            O => \N__43067\,
            I => \N__43054\
        );

    \I__9760\ : Span12Mux_s2_v
    port map (
            O => \N__43064\,
            I => \N__43047\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__43061\,
            I => \N__43047\
        );

    \I__9758\ : LocalMux
    port map (
            O => \N__43058\,
            I => \N__43047\
        );

    \I__9757\ : InMux
    port map (
            O => \N__43057\,
            I => \N__43044\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__43054\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__9755\ : Odrv12
    port map (
            O => \N__43047\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__9754\ : LocalMux
    port map (
            O => \N__43044\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__9753\ : IoInMux
    port map (
            O => \N__43037\,
            I => \N__43034\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__43034\,
            I => \N__43031\
        );

    \I__9751\ : IoSpan4Mux
    port map (
            O => \N__43031\,
            I => \N__43028\
        );

    \I__9750\ : Odrv4
    port map (
            O => \N__43028\,
            I => s2_phy_c
        );

    \I__9749\ : InMux
    port map (
            O => \N__43025\,
            I => \N__43021\
        );

    \I__9748\ : InMux
    port map (
            O => \N__43024\,
            I => \N__43018\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__43021\,
            I => \N__43013\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__43018\,
            I => \N__43013\
        );

    \I__9745\ : Span4Mux_s3_v
    port map (
            O => \N__43013\,
            I => \N__43010\
        );

    \I__9744\ : Sp12to4
    port map (
            O => \N__43010\,
            I => \N__43007\
        );

    \I__9743\ : Span12Mux_s6_h
    port map (
            O => \N__43007\,
            I => \N__43003\
        );

    \I__9742\ : InMux
    port map (
            O => \N__43006\,
            I => \N__43000\
        );

    \I__9741\ : Span12Mux_v
    port map (
            O => \N__43003\,
            I => \N__42996\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__43000\,
            I => \N__42993\
        );

    \I__9739\ : InMux
    port map (
            O => \N__42999\,
            I => \N__42990\
        );

    \I__9738\ : Span12Mux_v
    port map (
            O => \N__42996\,
            I => \N__42987\
        );

    \I__9737\ : Span4Mux_v
    port map (
            O => \N__42993\,
            I => \N__42984\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__42990\,
            I => \N__42981\
        );

    \I__9735\ : Span12Mux_h
    port map (
            O => \N__42987\,
            I => \N__42978\
        );

    \I__9734\ : Span4Mux_h
    port map (
            O => \N__42984\,
            I => \N__42973\
        );

    \I__9733\ : Span4Mux_v
    port map (
            O => \N__42981\,
            I => \N__42973\
        );

    \I__9732\ : Odrv12
    port map (
            O => \N__42978\,
            I => start_stop_c
        );

    \I__9731\ : Odrv4
    port map (
            O => \N__42973\,
            I => start_stop_c
        );

    \I__9730\ : CascadeMux
    port map (
            O => \N__42968\,
            I => \N__42963\
        );

    \I__9729\ : InMux
    port map (
            O => \N__42967\,
            I => \N__42959\
        );

    \I__9728\ : InMux
    port map (
            O => \N__42966\,
            I => \N__42956\
        );

    \I__9727\ : InMux
    port map (
            O => \N__42963\,
            I => \N__42953\
        );

    \I__9726\ : InMux
    port map (
            O => \N__42962\,
            I => \N__42950\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__42959\,
            I => \N__42947\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__42956\,
            I => \N__42942\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__42953\,
            I => \N__42942\
        );

    \I__9722\ : LocalMux
    port map (
            O => \N__42950\,
            I => \N__42936\
        );

    \I__9721\ : Span4Mux_h
    port map (
            O => \N__42947\,
            I => \N__42936\
        );

    \I__9720\ : Span4Mux_v
    port map (
            O => \N__42942\,
            I => \N__42933\
        );

    \I__9719\ : InMux
    port map (
            O => \N__42941\,
            I => \N__42930\
        );

    \I__9718\ : Span4Mux_v
    port map (
            O => \N__42936\,
            I => \N__42926\
        );

    \I__9717\ : Span4Mux_v
    port map (
            O => \N__42933\,
            I => \N__42921\
        );

    \I__9716\ : LocalMux
    port map (
            O => \N__42930\,
            I => \N__42921\
        );

    \I__9715\ : InMux
    port map (
            O => \N__42929\,
            I => \N__42918\
        );

    \I__9714\ : Span4Mux_v
    port map (
            O => \N__42926\,
            I => \N__42913\
        );

    \I__9713\ : Span4Mux_h
    port map (
            O => \N__42921\,
            I => \N__42913\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__42918\,
            I => phase_controller_inst1_state_4
        );

    \I__9711\ : Odrv4
    port map (
            O => \N__42913\,
            I => phase_controller_inst1_state_4
        );

    \I__9710\ : CascadeMux
    port map (
            O => \N__42908\,
            I => \N__42904\
        );

    \I__9709\ : InMux
    port map (
            O => \N__42907\,
            I => \N__42901\
        );

    \I__9708\ : InMux
    port map (
            O => \N__42904\,
            I => \N__42898\
        );

    \I__9707\ : LocalMux
    port map (
            O => \N__42901\,
            I => \N__42895\
        );

    \I__9706\ : LocalMux
    port map (
            O => \N__42898\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__9705\ : Odrv12
    port map (
            O => \N__42895\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__9704\ : InMux
    port map (
            O => \N__42890\,
            I => \N__42884\
        );

    \I__9703\ : InMux
    port map (
            O => \N__42889\,
            I => \N__42884\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__42884\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__9701\ : InMux
    port map (
            O => \N__42881\,
            I => \N__42875\
        );

    \I__9700\ : InMux
    port map (
            O => \N__42880\,
            I => \N__42875\
        );

    \I__9699\ : LocalMux
    port map (
            O => \N__42875\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__9698\ : CascadeMux
    port map (
            O => \N__42872\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__9697\ : InMux
    port map (
            O => \N__42869\,
            I => \N__42863\
        );

    \I__9696\ : InMux
    port map (
            O => \N__42868\,
            I => \N__42863\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__42863\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__9694\ : InMux
    port map (
            O => \N__42860\,
            I => \N__42854\
        );

    \I__9693\ : InMux
    port map (
            O => \N__42859\,
            I => \N__42854\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__42854\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__9691\ : InMux
    port map (
            O => \N__42851\,
            I => \N__42845\
        );

    \I__9690\ : InMux
    port map (
            O => \N__42850\,
            I => \N__42845\
        );

    \I__9689\ : LocalMux
    port map (
            O => \N__42845\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__9688\ : InMux
    port map (
            O => \N__42842\,
            I => \N__42836\
        );

    \I__9687\ : InMux
    port map (
            O => \N__42841\,
            I => \N__42836\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__42836\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__9685\ : InMux
    port map (
            O => \N__42833\,
            I => \N__42827\
        );

    \I__9684\ : InMux
    port map (
            O => \N__42832\,
            I => \N__42827\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__42827\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__9682\ : InMux
    port map (
            O => \N__42824\,
            I => \N__42820\
        );

    \I__9681\ : InMux
    port map (
            O => \N__42823\,
            I => \N__42817\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__42820\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__9679\ : LocalMux
    port map (
            O => \N__42817\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__9678\ : CascadeMux
    port map (
            O => \N__42812\,
            I => \N__42809\
        );

    \I__9677\ : InMux
    port map (
            O => \N__42809\,
            I => \N__42805\
        );

    \I__9676\ : InMux
    port map (
            O => \N__42808\,
            I => \N__42802\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__42805\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__42802\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__9673\ : CascadeMux
    port map (
            O => \N__42797\,
            I => \N__42794\
        );

    \I__9672\ : InMux
    port map (
            O => \N__42794\,
            I => \N__42791\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__42791\,
            I => \N__42787\
        );

    \I__9670\ : InMux
    port map (
            O => \N__42790\,
            I => \N__42784\
        );

    \I__9669\ : Odrv4
    port map (
            O => \N__42787\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__9668\ : LocalMux
    port map (
            O => \N__42784\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__9667\ : InMux
    port map (
            O => \N__42779\,
            I => \N__42776\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__42776\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__9665\ : InMux
    port map (
            O => \N__42773\,
            I => \N__42769\
        );

    \I__9664\ : InMux
    port map (
            O => \N__42772\,
            I => \N__42766\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__42769\,
            I => \N__42763\
        );

    \I__9662\ : LocalMux
    port map (
            O => \N__42766\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__9661\ : Odrv4
    port map (
            O => \N__42763\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__9660\ : CascadeMux
    port map (
            O => \N__42758\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\
        );

    \I__9659\ : CascadeMux
    port map (
            O => \N__42755\,
            I => \N__42751\
        );

    \I__9658\ : InMux
    port map (
            O => \N__42754\,
            I => \N__42748\
        );

    \I__9657\ : InMux
    port map (
            O => \N__42751\,
            I => \N__42745\
        );

    \I__9656\ : LocalMux
    port map (
            O => \N__42748\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__42745\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__9654\ : InMux
    port map (
            O => \N__42740\,
            I => \N__42734\
        );

    \I__9653\ : InMux
    port map (
            O => \N__42739\,
            I => \N__42734\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__42734\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__9651\ : InMux
    port map (
            O => \N__42731\,
            I => \N__42725\
        );

    \I__9650\ : InMux
    port map (
            O => \N__42730\,
            I => \N__42725\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__42725\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__9648\ : ClkMux
    port map (
            O => \N__42722\,
            I => \N__42716\
        );

    \I__9647\ : ClkMux
    port map (
            O => \N__42721\,
            I => \N__42716\
        );

    \I__9646\ : GlobalMux
    port map (
            O => \N__42716\,
            I => \N__42713\
        );

    \I__9645\ : gio2CtrlBuf
    port map (
            O => \N__42713\,
            I => delay_tr_input_c_g
        );

    \I__9644\ : CascadeMux
    port map (
            O => \N__42710\,
            I => \N__42705\
        );

    \I__9643\ : InMux
    port map (
            O => \N__42709\,
            I => \N__42700\
        );

    \I__9642\ : InMux
    port map (
            O => \N__42708\,
            I => \N__42700\
        );

    \I__9641\ : InMux
    port map (
            O => \N__42705\,
            I => \N__42696\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__42700\,
            I => \N__42693\
        );

    \I__9639\ : InMux
    port map (
            O => \N__42699\,
            I => \N__42690\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__42696\,
            I => \N__42687\
        );

    \I__9637\ : Span4Mux_v
    port map (
            O => \N__42693\,
            I => \N__42684\
        );

    \I__9636\ : LocalMux
    port map (
            O => \N__42690\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__9635\ : Odrv4
    port map (
            O => \N__42687\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__9634\ : Odrv4
    port map (
            O => \N__42684\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__9633\ : InMux
    port map (
            O => \N__42677\,
            I => \N__42674\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__42674\,
            I => \N__42671\
        );

    \I__9631\ : Odrv4
    port map (
            O => \N__42671\,
            I => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\
        );

    \I__9630\ : InMux
    port map (
            O => \N__42668\,
            I => \N__42664\
        );

    \I__9629\ : InMux
    port map (
            O => \N__42667\,
            I => \N__42661\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__42664\,
            I => \phase_controller_inst1.state_RNIE87FZ0Z_2\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__42661\,
            I => \phase_controller_inst1.state_RNIE87FZ0Z_2\
        );

    \I__9626\ : IoInMux
    port map (
            O => \N__42656\,
            I => \N__42653\
        );

    \I__9625\ : LocalMux
    port map (
            O => \N__42653\,
            I => \N__42649\
        );

    \I__9624\ : InMux
    port map (
            O => \N__42652\,
            I => \N__42646\
        );

    \I__9623\ : Odrv12
    port map (
            O => \N__42649\,
            I => \T45_c\
        );

    \I__9622\ : LocalMux
    port map (
            O => \N__42646\,
            I => \T45_c\
        );

    \I__9621\ : CascadeMux
    port map (
            O => \N__42641\,
            I => \N__42638\
        );

    \I__9620\ : InMux
    port map (
            O => \N__42638\,
            I => \N__42635\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__42635\,
            I => \N__42630\
        );

    \I__9618\ : InMux
    port map (
            O => \N__42634\,
            I => \N__42627\
        );

    \I__9617\ : InMux
    port map (
            O => \N__42633\,
            I => \N__42624\
        );

    \I__9616\ : Span4Mux_v
    port map (
            O => \N__42630\,
            I => \N__42619\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__42627\,
            I => \N__42619\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__42624\,
            I => \N__42616\
        );

    \I__9613\ : Span4Mux_v
    port map (
            O => \N__42619\,
            I => \N__42613\
        );

    \I__9612\ : Span4Mux_h
    port map (
            O => \N__42616\,
            I => \N__42610\
        );

    \I__9611\ : Span4Mux_h
    port map (
            O => \N__42613\,
            I => \N__42607\
        );

    \I__9610\ : Span4Mux_h
    port map (
            O => \N__42610\,
            I => \N__42604\
        );

    \I__9609\ : Span4Mux_v
    port map (
            O => \N__42607\,
            I => \N__42601\
        );

    \I__9608\ : Span4Mux_v
    port map (
            O => \N__42604\,
            I => \N__42598\
        );

    \I__9607\ : Odrv4
    port map (
            O => \N__42601\,
            I => \il_min_comp1_D2\
        );

    \I__9606\ : Odrv4
    port map (
            O => \N__42598\,
            I => \il_min_comp1_D2\
        );

    \I__9605\ : IoInMux
    port map (
            O => \N__42593\,
            I => \N__42590\
        );

    \I__9604\ : LocalMux
    port map (
            O => \N__42590\,
            I => \N__42587\
        );

    \I__9603\ : Span12Mux_s7_v
    port map (
            O => \N__42587\,
            I => \N__42583\
        );

    \I__9602\ : InMux
    port map (
            O => \N__42586\,
            I => \N__42580\
        );

    \I__9601\ : Odrv12
    port map (
            O => \N__42583\,
            I => \T23_c\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__42580\,
            I => \T23_c\
        );

    \I__9599\ : InMux
    port map (
            O => \N__42575\,
            I => \N__42572\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__42572\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__9597\ : CascadeMux
    port map (
            O => \N__42569\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18_cascade_\
        );

    \I__9596\ : InMux
    port map (
            O => \N__42566\,
            I => \N__42563\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__42563\,
            I => \N__42560\
        );

    \I__9594\ : Span4Mux_h
    port map (
            O => \N__42560\,
            I => \N__42557\
        );

    \I__9593\ : Odrv4
    port map (
            O => \N__42557\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\
        );

    \I__9592\ : InMux
    port map (
            O => \N__42554\,
            I => \N__42549\
        );

    \I__9591\ : InMux
    port map (
            O => \N__42553\,
            I => \N__42546\
        );

    \I__9590\ : InMux
    port map (
            O => \N__42552\,
            I => \N__42543\
        );

    \I__9589\ : LocalMux
    port map (
            O => \N__42549\,
            I => \N__42540\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__42546\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__9587\ : LocalMux
    port map (
            O => \N__42543\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__9586\ : Odrv12
    port map (
            O => \N__42540\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__9585\ : InMux
    port map (
            O => \N__42533\,
            I => \N__42530\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__42530\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\
        );

    \I__9583\ : InMux
    port map (
            O => \N__42527\,
            I => \N__42524\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__42524\,
            I => \N__42519\
        );

    \I__9581\ : InMux
    port map (
            O => \N__42523\,
            I => \N__42516\
        );

    \I__9580\ : InMux
    port map (
            O => \N__42522\,
            I => \N__42513\
        );

    \I__9579\ : Span4Mux_h
    port map (
            O => \N__42519\,
            I => \N__42507\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__42516\,
            I => \N__42507\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__42513\,
            I => \N__42504\
        );

    \I__9576\ : InMux
    port map (
            O => \N__42512\,
            I => \N__42501\
        );

    \I__9575\ : Odrv4
    port map (
            O => \N__42507\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__9574\ : Odrv4
    port map (
            O => \N__42504\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__9573\ : LocalMux
    port map (
            O => \N__42501\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__9572\ : InMux
    port map (
            O => \N__42494\,
            I => \N__42491\
        );

    \I__9571\ : LocalMux
    port map (
            O => \N__42491\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\
        );

    \I__9570\ : InMux
    port map (
            O => \N__42488\,
            I => \N__42483\
        );

    \I__9569\ : InMux
    port map (
            O => \N__42487\,
            I => \N__42480\
        );

    \I__9568\ : InMux
    port map (
            O => \N__42486\,
            I => \N__42477\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__42483\,
            I => \N__42474\
        );

    \I__9566\ : LocalMux
    port map (
            O => \N__42480\,
            I => \N__42470\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__42477\,
            I => \N__42465\
        );

    \I__9564\ : Span4Mux_h
    port map (
            O => \N__42474\,
            I => \N__42465\
        );

    \I__9563\ : InMux
    port map (
            O => \N__42473\,
            I => \N__42462\
        );

    \I__9562\ : Odrv12
    port map (
            O => \N__42470\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__9561\ : Odrv4
    port map (
            O => \N__42465\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__42462\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__9559\ : InMux
    port map (
            O => \N__42455\,
            I => \N__42452\
        );

    \I__9558\ : LocalMux
    port map (
            O => \N__42452\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\
        );

    \I__9557\ : InMux
    port map (
            O => \N__42449\,
            I => \N__42446\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__42446\,
            I => \N__42442\
        );

    \I__9555\ : InMux
    port map (
            O => \N__42445\,
            I => \N__42438\
        );

    \I__9554\ : Span4Mux_h
    port map (
            O => \N__42442\,
            I => \N__42435\
        );

    \I__9553\ : InMux
    port map (
            O => \N__42441\,
            I => \N__42432\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__42438\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__9551\ : Odrv4
    port map (
            O => \N__42435\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__42432\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__9549\ : InMux
    port map (
            O => \N__42425\,
            I => \N__42422\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__42422\,
            I => \N__42419\
        );

    \I__9547\ : Span4Mux_h
    port map (
            O => \N__42419\,
            I => \N__42414\
        );

    \I__9546\ : InMux
    port map (
            O => \N__42418\,
            I => \N__42408\
        );

    \I__9545\ : InMux
    port map (
            O => \N__42417\,
            I => \N__42408\
        );

    \I__9544\ : Span4Mux_v
    port map (
            O => \N__42414\,
            I => \N__42405\
        );

    \I__9543\ : InMux
    port map (
            O => \N__42413\,
            I => \N__42402\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__42408\,
            I => \N__42399\
        );

    \I__9541\ : Odrv4
    port map (
            O => \N__42405\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__42402\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__9539\ : Odrv4
    port map (
            O => \N__42399\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__9538\ : InMux
    port map (
            O => \N__42392\,
            I => \N__42389\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__42389\,
            I => \N__42385\
        );

    \I__9536\ : CascadeMux
    port map (
            O => \N__42388\,
            I => \N__42381\
        );

    \I__9535\ : Sp12to4
    port map (
            O => \N__42385\,
            I => \N__42377\
        );

    \I__9534\ : InMux
    port map (
            O => \N__42384\,
            I => \N__42374\
        );

    \I__9533\ : InMux
    port map (
            O => \N__42381\,
            I => \N__42371\
        );

    \I__9532\ : InMux
    port map (
            O => \N__42380\,
            I => \N__42368\
        );

    \I__9531\ : Span12Mux_s11_v
    port map (
            O => \N__42377\,
            I => \N__42365\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__42374\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__42371\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__42368\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__9527\ : Odrv12
    port map (
            O => \N__42365\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__9526\ : InMux
    port map (
            O => \N__42356\,
            I => \N__42352\
        );

    \I__9525\ : InMux
    port map (
            O => \N__42355\,
            I => \N__42349\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__42352\,
            I => \N__42345\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__42349\,
            I => \N__42341\
        );

    \I__9522\ : InMux
    port map (
            O => \N__42348\,
            I => \N__42337\
        );

    \I__9521\ : Span4Mux_h
    port map (
            O => \N__42345\,
            I => \N__42334\
        );

    \I__9520\ : InMux
    port map (
            O => \N__42344\,
            I => \N__42331\
        );

    \I__9519\ : Span4Mux_v
    port map (
            O => \N__42341\,
            I => \N__42328\
        );

    \I__9518\ : CascadeMux
    port map (
            O => \N__42340\,
            I => \N__42325\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__42337\,
            I => \N__42322\
        );

    \I__9516\ : Span4Mux_v
    port map (
            O => \N__42334\,
            I => \N__42319\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__42331\,
            I => \N__42316\
        );

    \I__9514\ : Span4Mux_v
    port map (
            O => \N__42328\,
            I => \N__42313\
        );

    \I__9513\ : InMux
    port map (
            O => \N__42325\,
            I => \N__42310\
        );

    \I__9512\ : Span12Mux_h
    port map (
            O => \N__42322\,
            I => \N__42307\
        );

    \I__9511\ : Span4Mux_v
    port map (
            O => \N__42319\,
            I => \N__42302\
        );

    \I__9510\ : Span4Mux_h
    port map (
            O => \N__42316\,
            I => \N__42302\
        );

    \I__9509\ : Span4Mux_h
    port map (
            O => \N__42313\,
            I => \N__42299\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__42310\,
            I => \N__42294\
        );

    \I__9507\ : Span12Mux_v
    port map (
            O => \N__42307\,
            I => \N__42294\
        );

    \I__9506\ : Odrv4
    port map (
            O => \N__42302\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__9505\ : Odrv4
    port map (
            O => \N__42299\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__9504\ : Odrv12
    port map (
            O => \N__42294\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__9503\ : CascadeMux
    port map (
            O => \N__42287\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__9502\ : InMux
    port map (
            O => \N__42284\,
            I => \N__42281\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__42281\,
            I => \N__42278\
        );

    \I__9500\ : Span4Mux_h
    port map (
            O => \N__42278\,
            I => \N__42274\
        );

    \I__9499\ : InMux
    port map (
            O => \N__42277\,
            I => \N__42271\
        );

    \I__9498\ : Odrv4
    port map (
            O => \N__42274\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__9497\ : LocalMux
    port map (
            O => \N__42271\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__9496\ : InMux
    port map (
            O => \N__42266\,
            I => \N__42263\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__42263\,
            I => \N__42259\
        );

    \I__9494\ : InMux
    port map (
            O => \N__42262\,
            I => \N__42255\
        );

    \I__9493\ : Span4Mux_h
    port map (
            O => \N__42259\,
            I => \N__42252\
        );

    \I__9492\ : InMux
    port map (
            O => \N__42258\,
            I => \N__42249\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__42255\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__9490\ : Odrv4
    port map (
            O => \N__42252\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__42249\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__9488\ : InMux
    port map (
            O => \N__42242\,
            I => \N__42236\
        );

    \I__9487\ : InMux
    port map (
            O => \N__42241\,
            I => \N__42236\
        );

    \I__9486\ : LocalMux
    port map (
            O => \N__42236\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__9485\ : InMux
    port map (
            O => \N__42233\,
            I => \N__42227\
        );

    \I__9484\ : InMux
    port map (
            O => \N__42232\,
            I => \N__42227\
        );

    \I__9483\ : LocalMux
    port map (
            O => \N__42227\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__9482\ : InMux
    port map (
            O => \N__42224\,
            I => \N__42221\
        );

    \I__9481\ : LocalMux
    port map (
            O => \N__42221\,
            I => \N__42217\
        );

    \I__9480\ : InMux
    port map (
            O => \N__42220\,
            I => \N__42213\
        );

    \I__9479\ : Span4Mux_h
    port map (
            O => \N__42217\,
            I => \N__42210\
        );

    \I__9478\ : InMux
    port map (
            O => \N__42216\,
            I => \N__42207\
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__42213\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__9476\ : Odrv4
    port map (
            O => \N__42210\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__42207\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__9474\ : InMux
    port map (
            O => \N__42200\,
            I => \N__42194\
        );

    \I__9473\ : InMux
    port map (
            O => \N__42199\,
            I => \N__42194\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__42194\,
            I => \N__42189\
        );

    \I__9471\ : InMux
    port map (
            O => \N__42193\,
            I => \N__42186\
        );

    \I__9470\ : InMux
    port map (
            O => \N__42192\,
            I => \N__42183\
        );

    \I__9469\ : Span4Mux_h
    port map (
            O => \N__42189\,
            I => \N__42180\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__42186\,
            I => \N__42175\
        );

    \I__9467\ : LocalMux
    port map (
            O => \N__42183\,
            I => \N__42175\
        );

    \I__9466\ : Odrv4
    port map (
            O => \N__42180\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__9465\ : Odrv4
    port map (
            O => \N__42175\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__9464\ : InMux
    port map (
            O => \N__42170\,
            I => \N__42166\
        );

    \I__9463\ : InMux
    port map (
            O => \N__42169\,
            I => \N__42161\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__42166\,
            I => \N__42158\
        );

    \I__9461\ : InMux
    port map (
            O => \N__42165\,
            I => \N__42155\
        );

    \I__9460\ : CascadeMux
    port map (
            O => \N__42164\,
            I => \N__42152\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__42161\,
            I => \N__42145\
        );

    \I__9458\ : Span4Mux_h
    port map (
            O => \N__42158\,
            I => \N__42145\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__42155\,
            I => \N__42145\
        );

    \I__9456\ : InMux
    port map (
            O => \N__42152\,
            I => \N__42142\
        );

    \I__9455\ : Odrv4
    port map (
            O => \N__42145\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__42142\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__9453\ : CascadeMux
    port map (
            O => \N__42137\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_\
        );

    \I__9452\ : CascadeMux
    port map (
            O => \N__42134\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\
        );

    \I__9451\ : InMux
    port map (
            O => \N__42131\,
            I => \N__42128\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__42128\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\
        );

    \I__9449\ : CascadeMux
    port map (
            O => \N__42125\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\
        );

    \I__9448\ : InMux
    port map (
            O => \N__42122\,
            I => \N__42119\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__42119\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\
        );

    \I__9446\ : InMux
    port map (
            O => \N__42116\,
            I => \N__42112\
        );

    \I__9445\ : InMux
    port map (
            O => \N__42115\,
            I => \N__42109\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__42112\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__9443\ : LocalMux
    port map (
            O => \N__42109\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__9442\ : InMux
    port map (
            O => \N__42104\,
            I => \N__42098\
        );

    \I__9441\ : InMux
    port map (
            O => \N__42103\,
            I => \N__42091\
        );

    \I__9440\ : InMux
    port map (
            O => \N__42102\,
            I => \N__42091\
        );

    \I__9439\ : InMux
    port map (
            O => \N__42101\,
            I => \N__42091\
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__42098\,
            I => \N__42086\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__42091\,
            I => \N__42086\
        );

    \I__9436\ : Span4Mux_h
    port map (
            O => \N__42086\,
            I => \N__42083\
        );

    \I__9435\ : Odrv4
    port map (
            O => \N__42083\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__9434\ : CascadeMux
    port map (
            O => \N__42080\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\
        );

    \I__9433\ : CascadeMux
    port map (
            O => \N__42077\,
            I => \N__42073\
        );

    \I__9432\ : InMux
    port map (
            O => \N__42076\,
            I => \N__42066\
        );

    \I__9431\ : InMux
    port map (
            O => \N__42073\,
            I => \N__42066\
        );

    \I__9430\ : InMux
    port map (
            O => \N__42072\,
            I => \N__42061\
        );

    \I__9429\ : InMux
    port map (
            O => \N__42071\,
            I => \N__42061\
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__42066\,
            I => \N__42058\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__42061\,
            I => \N__42053\
        );

    \I__9426\ : Span4Mux_h
    port map (
            O => \N__42058\,
            I => \N__42053\
        );

    \I__9425\ : Odrv4
    port map (
            O => \N__42053\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__9424\ : InMux
    port map (
            O => \N__42050\,
            I => \N__42046\
        );

    \I__9423\ : InMux
    port map (
            O => \N__42049\,
            I => \N__42043\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__42046\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__42043\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__9420\ : CascadeMux
    port map (
            O => \N__42038\,
            I => \N__42035\
        );

    \I__9419\ : InMux
    port map (
            O => \N__42035\,
            I => \N__42032\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__42032\,
            I => \N__42029\
        );

    \I__9417\ : Odrv4
    port map (
            O => \N__42029\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt26\
        );

    \I__9416\ : InMux
    port map (
            O => \N__42026\,
            I => \N__42020\
        );

    \I__9415\ : InMux
    port map (
            O => \N__42025\,
            I => \N__42020\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__42020\,
            I => \N__42016\
        );

    \I__9413\ : InMux
    port map (
            O => \N__42019\,
            I => \N__42013\
        );

    \I__9412\ : Span4Mux_h
    port map (
            O => \N__42016\,
            I => \N__42010\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__42013\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__9410\ : Odrv4
    port map (
            O => \N__42010\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__9409\ : CascadeMux
    port map (
            O => \N__42005\,
            I => \N__42001\
        );

    \I__9408\ : CascadeMux
    port map (
            O => \N__42004\,
            I => \N__41998\
        );

    \I__9407\ : InMux
    port map (
            O => \N__42001\,
            I => \N__41995\
        );

    \I__9406\ : InMux
    port map (
            O => \N__41998\,
            I => \N__41992\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__41995\,
            I => \N__41987\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__41992\,
            I => \N__41987\
        );

    \I__9403\ : Span4Mux_h
    port map (
            O => \N__41987\,
            I => \N__41983\
        );

    \I__9402\ : InMux
    port map (
            O => \N__41986\,
            I => \N__41980\
        );

    \I__9401\ : Span4Mux_h
    port map (
            O => \N__41983\,
            I => \N__41977\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__41980\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__9399\ : Odrv4
    port map (
            O => \N__41977\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__9398\ : InMux
    port map (
            O => \N__41972\,
            I => \N__41968\
        );

    \I__9397\ : InMux
    port map (
            O => \N__41971\,
            I => \N__41965\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__41968\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__41965\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\
        );

    \I__9394\ : InMux
    port map (
            O => \N__41960\,
            I => \N__41957\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__41957\,
            I => \N__41954\
        );

    \I__9392\ : Odrv4
    port map (
            O => \N__41954\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\
        );

    \I__9391\ : InMux
    port map (
            O => \N__41951\,
            I => \N__41948\
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__41948\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\
        );

    \I__9389\ : InMux
    port map (
            O => \N__41945\,
            I => \N__41939\
        );

    \I__9388\ : InMux
    port map (
            O => \N__41944\,
            I => \N__41936\
        );

    \I__9387\ : CascadeMux
    port map (
            O => \N__41943\,
            I => \N__41933\
        );

    \I__9386\ : InMux
    port map (
            O => \N__41942\,
            I => \N__41930\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__41939\,
            I => \N__41927\
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__41936\,
            I => \N__41924\
        );

    \I__9383\ : InMux
    port map (
            O => \N__41933\,
            I => \N__41921\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__41930\,
            I => \N__41914\
        );

    \I__9381\ : Span4Mux_v
    port map (
            O => \N__41927\,
            I => \N__41914\
        );

    \I__9380\ : Span4Mux_h
    port map (
            O => \N__41924\,
            I => \N__41914\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__41921\,
            I => \N__41911\
        );

    \I__9378\ : Span4Mux_h
    port map (
            O => \N__41914\,
            I => \N__41906\
        );

    \I__9377\ : Span4Mux_v
    port map (
            O => \N__41911\,
            I => \N__41906\
        );

    \I__9376\ : Odrv4
    port map (
            O => \N__41906\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__9375\ : InMux
    port map (
            O => \N__41903\,
            I => \N__41875\
        );

    \I__9374\ : InMux
    port map (
            O => \N__41902\,
            I => \N__41868\
        );

    \I__9373\ : InMux
    port map (
            O => \N__41901\,
            I => \N__41868\
        );

    \I__9372\ : InMux
    port map (
            O => \N__41900\,
            I => \N__41868\
        );

    \I__9371\ : InMux
    port map (
            O => \N__41899\,
            I => \N__41865\
        );

    \I__9370\ : InMux
    port map (
            O => \N__41898\,
            I => \N__41862\
        );

    \I__9369\ : InMux
    port map (
            O => \N__41897\,
            I => \N__41844\
        );

    \I__9368\ : InMux
    port map (
            O => \N__41896\,
            I => \N__41844\
        );

    \I__9367\ : InMux
    port map (
            O => \N__41895\,
            I => \N__41841\
        );

    \I__9366\ : InMux
    port map (
            O => \N__41894\,
            I => \N__41834\
        );

    \I__9365\ : InMux
    port map (
            O => \N__41893\,
            I => \N__41834\
        );

    \I__9364\ : InMux
    port map (
            O => \N__41892\,
            I => \N__41834\
        );

    \I__9363\ : InMux
    port map (
            O => \N__41891\,
            I => \N__41829\
        );

    \I__9362\ : InMux
    port map (
            O => \N__41890\,
            I => \N__41826\
        );

    \I__9361\ : InMux
    port map (
            O => \N__41889\,
            I => \N__41822\
        );

    \I__9360\ : InMux
    port map (
            O => \N__41888\,
            I => \N__41817\
        );

    \I__9359\ : InMux
    port map (
            O => \N__41887\,
            I => \N__41811\
        );

    \I__9358\ : InMux
    port map (
            O => \N__41886\,
            I => \N__41806\
        );

    \I__9357\ : InMux
    port map (
            O => \N__41885\,
            I => \N__41806\
        );

    \I__9356\ : InMux
    port map (
            O => \N__41884\,
            I => \N__41803\
        );

    \I__9355\ : InMux
    port map (
            O => \N__41883\,
            I => \N__41796\
        );

    \I__9354\ : InMux
    port map (
            O => \N__41882\,
            I => \N__41796\
        );

    \I__9353\ : InMux
    port map (
            O => \N__41881\,
            I => \N__41796\
        );

    \I__9352\ : InMux
    port map (
            O => \N__41880\,
            I => \N__41776\
        );

    \I__9351\ : InMux
    port map (
            O => \N__41879\,
            I => \N__41765\
        );

    \I__9350\ : InMux
    port map (
            O => \N__41878\,
            I => \N__41762\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__41875\,
            I => \N__41757\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__41868\,
            I => \N__41757\
        );

    \I__9347\ : LocalMux
    port map (
            O => \N__41865\,
            I => \N__41752\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__41862\,
            I => \N__41752\
        );

    \I__9345\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41749\
        );

    \I__9344\ : InMux
    port map (
            O => \N__41860\,
            I => \N__41744\
        );

    \I__9343\ : InMux
    port map (
            O => \N__41859\,
            I => \N__41744\
        );

    \I__9342\ : InMux
    port map (
            O => \N__41858\,
            I => \N__41733\
        );

    \I__9341\ : InMux
    port map (
            O => \N__41857\,
            I => \N__41733\
        );

    \I__9340\ : InMux
    port map (
            O => \N__41856\,
            I => \N__41733\
        );

    \I__9339\ : InMux
    port map (
            O => \N__41855\,
            I => \N__41733\
        );

    \I__9338\ : InMux
    port map (
            O => \N__41854\,
            I => \N__41728\
        );

    \I__9337\ : InMux
    port map (
            O => \N__41853\,
            I => \N__41728\
        );

    \I__9336\ : InMux
    port map (
            O => \N__41852\,
            I => \N__41723\
        );

    \I__9335\ : InMux
    port map (
            O => \N__41851\,
            I => \N__41723\
        );

    \I__9334\ : InMux
    port map (
            O => \N__41850\,
            I => \N__41718\
        );

    \I__9333\ : InMux
    port map (
            O => \N__41849\,
            I => \N__41718\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__41844\,
            I => \N__41711\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__41841\,
            I => \N__41711\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__41834\,
            I => \N__41711\
        );

    \I__9329\ : InMux
    port map (
            O => \N__41833\,
            I => \N__41706\
        );

    \I__9328\ : InMux
    port map (
            O => \N__41832\,
            I => \N__41706\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__41829\,
            I => \N__41701\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__41826\,
            I => \N__41701\
        );

    \I__9325\ : InMux
    port map (
            O => \N__41825\,
            I => \N__41698\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__41822\,
            I => \N__41695\
        );

    \I__9323\ : InMux
    port map (
            O => \N__41821\,
            I => \N__41690\
        );

    \I__9322\ : InMux
    port map (
            O => \N__41820\,
            I => \N__41690\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__41817\,
            I => \N__41687\
        );

    \I__9320\ : InMux
    port map (
            O => \N__41816\,
            I => \N__41684\
        );

    \I__9319\ : InMux
    port map (
            O => \N__41815\,
            I => \N__41679\
        );

    \I__9318\ : InMux
    port map (
            O => \N__41814\,
            I => \N__41679\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__41811\,
            I => \N__41676\
        );

    \I__9316\ : LocalMux
    port map (
            O => \N__41806\,
            I => \N__41669\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__41803\,
            I => \N__41669\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__41796\,
            I => \N__41669\
        );

    \I__9313\ : InMux
    port map (
            O => \N__41795\,
            I => \N__41648\
        );

    \I__9312\ : InMux
    port map (
            O => \N__41794\,
            I => \N__41635\
        );

    \I__9311\ : InMux
    port map (
            O => \N__41793\,
            I => \N__41635\
        );

    \I__9310\ : InMux
    port map (
            O => \N__41792\,
            I => \N__41635\
        );

    \I__9309\ : InMux
    port map (
            O => \N__41791\,
            I => \N__41635\
        );

    \I__9308\ : InMux
    port map (
            O => \N__41790\,
            I => \N__41635\
        );

    \I__9307\ : InMux
    port map (
            O => \N__41789\,
            I => \N__41635\
        );

    \I__9306\ : InMux
    port map (
            O => \N__41788\,
            I => \N__41628\
        );

    \I__9305\ : InMux
    port map (
            O => \N__41787\,
            I => \N__41628\
        );

    \I__9304\ : InMux
    port map (
            O => \N__41786\,
            I => \N__41628\
        );

    \I__9303\ : InMux
    port map (
            O => \N__41785\,
            I => \N__41623\
        );

    \I__9302\ : InMux
    port map (
            O => \N__41784\,
            I => \N__41623\
        );

    \I__9301\ : InMux
    port map (
            O => \N__41783\,
            I => \N__41620\
        );

    \I__9300\ : InMux
    port map (
            O => \N__41782\,
            I => \N__41613\
        );

    \I__9299\ : InMux
    port map (
            O => \N__41781\,
            I => \N__41613\
        );

    \I__9298\ : InMux
    port map (
            O => \N__41780\,
            I => \N__41613\
        );

    \I__9297\ : InMux
    port map (
            O => \N__41779\,
            I => \N__41610\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__41776\,
            I => \N__41607\
        );

    \I__9295\ : InMux
    port map (
            O => \N__41775\,
            I => \N__41596\
        );

    \I__9294\ : InMux
    port map (
            O => \N__41774\,
            I => \N__41596\
        );

    \I__9293\ : InMux
    port map (
            O => \N__41773\,
            I => \N__41596\
        );

    \I__9292\ : InMux
    port map (
            O => \N__41772\,
            I => \N__41596\
        );

    \I__9291\ : InMux
    port map (
            O => \N__41771\,
            I => \N__41596\
        );

    \I__9290\ : InMux
    port map (
            O => \N__41770\,
            I => \N__41589\
        );

    \I__9289\ : InMux
    port map (
            O => \N__41769\,
            I => \N__41589\
        );

    \I__9288\ : InMux
    port map (
            O => \N__41768\,
            I => \N__41589\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__41765\,
            I => \N__41584\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__41762\,
            I => \N__41584\
        );

    \I__9285\ : Span4Mux_v
    port map (
            O => \N__41757\,
            I => \N__41577\
        );

    \I__9284\ : Span4Mux_v
    port map (
            O => \N__41752\,
            I => \N__41577\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__41749\,
            I => \N__41577\
        );

    \I__9282\ : LocalMux
    port map (
            O => \N__41744\,
            I => \N__41574\
        );

    \I__9281\ : InMux
    port map (
            O => \N__41743\,
            I => \N__41569\
        );

    \I__9280\ : InMux
    port map (
            O => \N__41742\,
            I => \N__41569\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__41733\,
            I => \N__41562\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__41728\,
            I => \N__41562\
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__41723\,
            I => \N__41562\
        );

    \I__9276\ : LocalMux
    port map (
            O => \N__41718\,
            I => \N__41551\
        );

    \I__9275\ : Span4Mux_h
    port map (
            O => \N__41711\,
            I => \N__41551\
        );

    \I__9274\ : LocalMux
    port map (
            O => \N__41706\,
            I => \N__41551\
        );

    \I__9273\ : Span4Mux_s3_v
    port map (
            O => \N__41701\,
            I => \N__41551\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__41698\,
            I => \N__41551\
        );

    \I__9271\ : Span4Mux_h
    port map (
            O => \N__41695\,
            I => \N__41548\
        );

    \I__9270\ : LocalMux
    port map (
            O => \N__41690\,
            I => \N__41543\
        );

    \I__9269\ : Span4Mux_v
    port map (
            O => \N__41687\,
            I => \N__41543\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__41684\,
            I => \N__41534\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__41679\,
            I => \N__41534\
        );

    \I__9266\ : Span4Mux_v
    port map (
            O => \N__41676\,
            I => \N__41534\
        );

    \I__9265\ : Span4Mux_v
    port map (
            O => \N__41669\,
            I => \N__41534\
        );

    \I__9264\ : InMux
    port map (
            O => \N__41668\,
            I => \N__41531\
        );

    \I__9263\ : InMux
    port map (
            O => \N__41667\,
            I => \N__41524\
        );

    \I__9262\ : InMux
    port map (
            O => \N__41666\,
            I => \N__41524\
        );

    \I__9261\ : InMux
    port map (
            O => \N__41665\,
            I => \N__41524\
        );

    \I__9260\ : InMux
    port map (
            O => \N__41664\,
            I => \N__41513\
        );

    \I__9259\ : InMux
    port map (
            O => \N__41663\,
            I => \N__41513\
        );

    \I__9258\ : InMux
    port map (
            O => \N__41662\,
            I => \N__41513\
        );

    \I__9257\ : InMux
    port map (
            O => \N__41661\,
            I => \N__41513\
        );

    \I__9256\ : InMux
    port map (
            O => \N__41660\,
            I => \N__41513\
        );

    \I__9255\ : InMux
    port map (
            O => \N__41659\,
            I => \N__41500\
        );

    \I__9254\ : InMux
    port map (
            O => \N__41658\,
            I => \N__41500\
        );

    \I__9253\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41500\
        );

    \I__9252\ : InMux
    port map (
            O => \N__41656\,
            I => \N__41500\
        );

    \I__9251\ : InMux
    port map (
            O => \N__41655\,
            I => \N__41500\
        );

    \I__9250\ : InMux
    port map (
            O => \N__41654\,
            I => \N__41500\
        );

    \I__9249\ : InMux
    port map (
            O => \N__41653\,
            I => \N__41497\
        );

    \I__9248\ : InMux
    port map (
            O => \N__41652\,
            I => \N__41492\
        );

    \I__9247\ : InMux
    port map (
            O => \N__41651\,
            I => \N__41492\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__41648\,
            I => \N__41485\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__41635\,
            I => \N__41485\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__41628\,
            I => \N__41485\
        );

    \I__9243\ : LocalMux
    port map (
            O => \N__41623\,
            I => \N__41482\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__41620\,
            I => \N__41477\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__41613\,
            I => \N__41477\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__41610\,
            I => \N__41474\
        );

    \I__9239\ : Span12Mux_s7_v
    port map (
            O => \N__41607\,
            I => \N__41471\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__41596\,
            I => \N__41462\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__41589\,
            I => \N__41462\
        );

    \I__9236\ : Span4Mux_h
    port map (
            O => \N__41584\,
            I => \N__41462\
        );

    \I__9235\ : Span4Mux_h
    port map (
            O => \N__41577\,
            I => \N__41462\
        );

    \I__9234\ : Span4Mux_v
    port map (
            O => \N__41574\,
            I => \N__41447\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__41569\,
            I => \N__41447\
        );

    \I__9232\ : Span4Mux_v
    port map (
            O => \N__41562\,
            I => \N__41447\
        );

    \I__9231\ : Span4Mux_v
    port map (
            O => \N__41551\,
            I => \N__41447\
        );

    \I__9230\ : Span4Mux_v
    port map (
            O => \N__41548\,
            I => \N__41447\
        );

    \I__9229\ : Span4Mux_h
    port map (
            O => \N__41543\,
            I => \N__41447\
        );

    \I__9228\ : Span4Mux_h
    port map (
            O => \N__41534\,
            I => \N__41447\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__41531\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__41524\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__9225\ : LocalMux
    port map (
            O => \N__41513\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__9224\ : LocalMux
    port map (
            O => \N__41500\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__41497\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__41492\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__9221\ : Odrv4
    port map (
            O => \N__41485\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__9220\ : Odrv4
    port map (
            O => \N__41482\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__9219\ : Odrv4
    port map (
            O => \N__41477\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__9218\ : Odrv12
    port map (
            O => \N__41474\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__9217\ : Odrv12
    port map (
            O => \N__41471\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__9216\ : Odrv4
    port map (
            O => \N__41462\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__9215\ : Odrv4
    port map (
            O => \N__41447\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__9214\ : InMux
    port map (
            O => \N__41420\,
            I => \N__41416\
        );

    \I__9213\ : InMux
    port map (
            O => \N__41419\,
            I => \N__41412\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__41416\,
            I => \N__41409\
        );

    \I__9211\ : InMux
    port map (
            O => \N__41415\,
            I => \N__41406\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__41412\,
            I => \N__41403\
        );

    \I__9209\ : Span12Mux_h
    port map (
            O => \N__41409\,
            I => \N__41400\
        );

    \I__9208\ : LocalMux
    port map (
            O => \N__41406\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__9207\ : Odrv12
    port map (
            O => \N__41403\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__9206\ : Odrv12
    port map (
            O => \N__41400\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__9205\ : InMux
    port map (
            O => \N__41393\,
            I => \N__41390\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__41390\,
            I => \N__41387\
        );

    \I__9203\ : Span4Mux_h
    port map (
            O => \N__41387\,
            I => \N__41383\
        );

    \I__9202\ : InMux
    port map (
            O => \N__41386\,
            I => \N__41380\
        );

    \I__9201\ : Odrv4
    port map (
            O => \N__41383\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__41380\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__9199\ : InMux
    port map (
            O => \N__41375\,
            I => \N__41372\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__41372\,
            I => \N__41368\
        );

    \I__9197\ : InMux
    port map (
            O => \N__41371\,
            I => \N__41364\
        );

    \I__9196\ : Span4Mux_h
    port map (
            O => \N__41368\,
            I => \N__41361\
        );

    \I__9195\ : InMux
    port map (
            O => \N__41367\,
            I => \N__41358\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__41364\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__9193\ : Odrv4
    port map (
            O => \N__41361\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__41358\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__9191\ : InMux
    port map (
            O => \N__41351\,
            I => \N__41345\
        );

    \I__9190\ : InMux
    port map (
            O => \N__41350\,
            I => \N__41345\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__41345\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__9188\ : CascadeMux
    port map (
            O => \N__41342\,
            I => \N__41339\
        );

    \I__9187\ : InMux
    port map (
            O => \N__41339\,
            I => \N__41333\
        );

    \I__9186\ : InMux
    port map (
            O => \N__41338\,
            I => \N__41333\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__41333\,
            I => \N__41330\
        );

    \I__9184\ : Odrv4
    port map (
            O => \N__41330\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\
        );

    \I__9183\ : CascadeMux
    port map (
            O => \N__41327\,
            I => \N__41324\
        );

    \I__9182\ : InMux
    port map (
            O => \N__41324\,
            I => \N__41321\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__41321\,
            I => \N__41318\
        );

    \I__9180\ : Odrv4
    port map (
            O => \N__41318\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__9179\ : CascadeMux
    port map (
            O => \N__41315\,
            I => \N__41311\
        );

    \I__9178\ : CascadeMux
    port map (
            O => \N__41314\,
            I => \N__41308\
        );

    \I__9177\ : InMux
    port map (
            O => \N__41311\,
            I => \N__41305\
        );

    \I__9176\ : InMux
    port map (
            O => \N__41308\,
            I => \N__41301\
        );

    \I__9175\ : LocalMux
    port map (
            O => \N__41305\,
            I => \N__41298\
        );

    \I__9174\ : InMux
    port map (
            O => \N__41304\,
            I => \N__41294\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__41301\,
            I => \N__41291\
        );

    \I__9172\ : Span12Mux_v
    port map (
            O => \N__41298\,
            I => \N__41288\
        );

    \I__9171\ : InMux
    port map (
            O => \N__41297\,
            I => \N__41285\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__41294\,
            I => \N__41280\
        );

    \I__9169\ : Span4Mux_v
    port map (
            O => \N__41291\,
            I => \N__41280\
        );

    \I__9168\ : Odrv12
    port map (
            O => \N__41288\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__41285\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__9166\ : Odrv4
    port map (
            O => \N__41280\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__9165\ : InMux
    port map (
            O => \N__41273\,
            I => \bfn_15_26_0_\
        );

    \I__9164\ : CascadeMux
    port map (
            O => \N__41270\,
            I => \N__41266\
        );

    \I__9163\ : InMux
    port map (
            O => \N__41269\,
            I => \N__41263\
        );

    \I__9162\ : InMux
    port map (
            O => \N__41266\,
            I => \N__41260\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__41263\,
            I => \N__41255\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__41260\,
            I => \N__41252\
        );

    \I__9159\ : InMux
    port map (
            O => \N__41259\,
            I => \N__41249\
        );

    \I__9158\ : InMux
    port map (
            O => \N__41258\,
            I => \N__41246\
        );

    \I__9157\ : Span12Mux_h
    port map (
            O => \N__41255\,
            I => \N__41239\
        );

    \I__9156\ : Sp12to4
    port map (
            O => \N__41252\,
            I => \N__41239\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__41249\,
            I => \N__41239\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__41246\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__9153\ : Odrv12
    port map (
            O => \N__41239\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__9152\ : InMux
    port map (
            O => \N__41234\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__9151\ : CascadeMux
    port map (
            O => \N__41231\,
            I => \N__41228\
        );

    \I__9150\ : InMux
    port map (
            O => \N__41228\,
            I => \N__41225\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__41225\,
            I => \N__41221\
        );

    \I__9148\ : InMux
    port map (
            O => \N__41224\,
            I => \N__41218\
        );

    \I__9147\ : Span4Mux_v
    port map (
            O => \N__41221\,
            I => \N__41215\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__41218\,
            I => \N__41212\
        );

    \I__9145\ : Sp12to4
    port map (
            O => \N__41215\,
            I => \N__41208\
        );

    \I__9144\ : Span4Mux_h
    port map (
            O => \N__41212\,
            I => \N__41204\
        );

    \I__9143\ : InMux
    port map (
            O => \N__41211\,
            I => \N__41201\
        );

    \I__9142\ : Span12Mux_h
    port map (
            O => \N__41208\,
            I => \N__41198\
        );

    \I__9141\ : InMux
    port map (
            O => \N__41207\,
            I => \N__41195\
        );

    \I__9140\ : Span4Mux_v
    port map (
            O => \N__41204\,
            I => \N__41192\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__41201\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__9138\ : Odrv12
    port map (
            O => \N__41198\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__41195\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__9136\ : Odrv4
    port map (
            O => \N__41192\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__9135\ : InMux
    port map (
            O => \N__41183\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__9134\ : InMux
    port map (
            O => \N__41180\,
            I => \N__41176\
        );

    \I__9133\ : InMux
    port map (
            O => \N__41179\,
            I => \N__41173\
        );

    \I__9132\ : LocalMux
    port map (
            O => \N__41176\,
            I => \N__41170\
        );

    \I__9131\ : LocalMux
    port map (
            O => \N__41173\,
            I => \N__41165\
        );

    \I__9130\ : Span12Mux_v
    port map (
            O => \N__41170\,
            I => \N__41162\
        );

    \I__9129\ : InMux
    port map (
            O => \N__41169\,
            I => \N__41159\
        );

    \I__9128\ : InMux
    port map (
            O => \N__41168\,
            I => \N__41156\
        );

    \I__9127\ : Span4Mux_v
    port map (
            O => \N__41165\,
            I => \N__41153\
        );

    \I__9126\ : Odrv12
    port map (
            O => \N__41162\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__41159\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__9124\ : LocalMux
    port map (
            O => \N__41156\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__9123\ : Odrv4
    port map (
            O => \N__41153\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__9122\ : InMux
    port map (
            O => \N__41144\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__9121\ : CascadeMux
    port map (
            O => \N__41141\,
            I => \N__41137\
        );

    \I__9120\ : InMux
    port map (
            O => \N__41140\,
            I => \N__41133\
        );

    \I__9119\ : InMux
    port map (
            O => \N__41137\,
            I => \N__41130\
        );

    \I__9118\ : InMux
    port map (
            O => \N__41136\,
            I => \N__41127\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__41133\,
            I => \N__41124\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__41130\,
            I => \N__41121\
        );

    \I__9115\ : LocalMux
    port map (
            O => \N__41127\,
            I => \N__41115\
        );

    \I__9114\ : Span4Mux_v
    port map (
            O => \N__41124\,
            I => \N__41115\
        );

    \I__9113\ : Span12Mux_v
    port map (
            O => \N__41121\,
            I => \N__41112\
        );

    \I__9112\ : InMux
    port map (
            O => \N__41120\,
            I => \N__41109\
        );

    \I__9111\ : Span4Mux_v
    port map (
            O => \N__41115\,
            I => \N__41106\
        );

    \I__9110\ : Odrv12
    port map (
            O => \N__41112\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__41109\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__9108\ : Odrv4
    port map (
            O => \N__41106\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__9107\ : InMux
    port map (
            O => \N__41099\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__9106\ : InMux
    port map (
            O => \N__41096\,
            I => \N__41093\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__41093\,
            I => \N__41089\
        );

    \I__9104\ : InMux
    port map (
            O => \N__41092\,
            I => \N__41085\
        );

    \I__9103\ : Span12Mux_s10_h
    port map (
            O => \N__41089\,
            I => \N__41082\
        );

    \I__9102\ : CascadeMux
    port map (
            O => \N__41088\,
            I => \N__41079\
        );

    \I__9101\ : LocalMux
    port map (
            O => \N__41085\,
            I => \N__41075\
        );

    \I__9100\ : Span12Mux_h
    port map (
            O => \N__41082\,
            I => \N__41072\
        );

    \I__9099\ : InMux
    port map (
            O => \N__41079\,
            I => \N__41069\
        );

    \I__9098\ : InMux
    port map (
            O => \N__41078\,
            I => \N__41066\
        );

    \I__9097\ : Span4Mux_v
    port map (
            O => \N__41075\,
            I => \N__41063\
        );

    \I__9096\ : Odrv12
    port map (
            O => \N__41072\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__41069\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__41066\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__9093\ : Odrv4
    port map (
            O => \N__41063\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__9092\ : InMux
    port map (
            O => \N__41054\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__9091\ : InMux
    port map (
            O => \N__41051\,
            I => \N__41047\
        );

    \I__9090\ : CascadeMux
    port map (
            O => \N__41050\,
            I => \N__41043\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__41047\,
            I => \N__41037\
        );

    \I__9088\ : InMux
    port map (
            O => \N__41046\,
            I => \N__41028\
        );

    \I__9087\ : InMux
    port map (
            O => \N__41043\,
            I => \N__41025\
        );

    \I__9086\ : InMux
    port map (
            O => \N__41042\,
            I => \N__41022\
        );

    \I__9085\ : InMux
    port map (
            O => \N__41041\,
            I => \N__41017\
        );

    \I__9084\ : InMux
    port map (
            O => \N__41040\,
            I => \N__41017\
        );

    \I__9083\ : Sp12to4
    port map (
            O => \N__41037\,
            I => \N__41014\
        );

    \I__9082\ : InMux
    port map (
            O => \N__41036\,
            I => \N__40992\
        );

    \I__9081\ : InMux
    port map (
            O => \N__41035\,
            I => \N__40989\
        );

    \I__9080\ : InMux
    port map (
            O => \N__41034\,
            I => \N__40980\
        );

    \I__9079\ : InMux
    port map (
            O => \N__41033\,
            I => \N__40980\
        );

    \I__9078\ : InMux
    port map (
            O => \N__41032\,
            I => \N__40980\
        );

    \I__9077\ : InMux
    port map (
            O => \N__41031\,
            I => \N__40980\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__41028\,
            I => \N__40977\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__41025\,
            I => \N__40972\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__41022\,
            I => \N__40972\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__41017\,
            I => \N__40968\
        );

    \I__9072\ : Span12Mux_v
    port map (
            O => \N__41014\,
            I => \N__40965\
        );

    \I__9071\ : InMux
    port map (
            O => \N__41013\,
            I => \N__40962\
        );

    \I__9070\ : InMux
    port map (
            O => \N__41012\,
            I => \N__40959\
        );

    \I__9069\ : InMux
    port map (
            O => \N__41011\,
            I => \N__40956\
        );

    \I__9068\ : InMux
    port map (
            O => \N__41010\,
            I => \N__40949\
        );

    \I__9067\ : InMux
    port map (
            O => \N__41009\,
            I => \N__40949\
        );

    \I__9066\ : InMux
    port map (
            O => \N__41008\,
            I => \N__40949\
        );

    \I__9065\ : InMux
    port map (
            O => \N__41007\,
            I => \N__40946\
        );

    \I__9064\ : InMux
    port map (
            O => \N__41006\,
            I => \N__40931\
        );

    \I__9063\ : InMux
    port map (
            O => \N__41005\,
            I => \N__40931\
        );

    \I__9062\ : InMux
    port map (
            O => \N__41004\,
            I => \N__40931\
        );

    \I__9061\ : InMux
    port map (
            O => \N__41003\,
            I => \N__40931\
        );

    \I__9060\ : InMux
    port map (
            O => \N__41002\,
            I => \N__40931\
        );

    \I__9059\ : InMux
    port map (
            O => \N__41001\,
            I => \N__40931\
        );

    \I__9058\ : InMux
    port map (
            O => \N__41000\,
            I => \N__40931\
        );

    \I__9057\ : InMux
    port map (
            O => \N__40999\,
            I => \N__40920\
        );

    \I__9056\ : InMux
    port map (
            O => \N__40998\,
            I => \N__40920\
        );

    \I__9055\ : InMux
    port map (
            O => \N__40997\,
            I => \N__40920\
        );

    \I__9054\ : InMux
    port map (
            O => \N__40996\,
            I => \N__40920\
        );

    \I__9053\ : InMux
    port map (
            O => \N__40995\,
            I => \N__40920\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__40992\,
            I => \N__40917\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__40989\,
            I => \N__40908\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__40980\,
            I => \N__40908\
        );

    \I__9049\ : Span4Mux_h
    port map (
            O => \N__40977\,
            I => \N__40908\
        );

    \I__9048\ : Span4Mux_h
    port map (
            O => \N__40972\,
            I => \N__40908\
        );

    \I__9047\ : InMux
    port map (
            O => \N__40971\,
            I => \N__40905\
        );

    \I__9046\ : Span12Mux_s4_h
    port map (
            O => \N__40968\,
            I => \N__40898\
        );

    \I__9045\ : Span12Mux_h
    port map (
            O => \N__40965\,
            I => \N__40898\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__40962\,
            I => \N__40898\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__40959\,
            I => \N__40895\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__40956\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__40949\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__40946\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__40931\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__40920\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9037\ : Odrv4
    port map (
            O => \N__40917\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9036\ : Odrv4
    port map (
            O => \N__40908\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__40905\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9034\ : Odrv12
    port map (
            O => \N__40898\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9033\ : Odrv4
    port map (
            O => \N__40895\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__9032\ : CascadeMux
    port map (
            O => \N__40874\,
            I => \N__40863\
        );

    \I__9031\ : CascadeMux
    port map (
            O => \N__40873\,
            I => \N__40859\
        );

    \I__9030\ : CascadeMux
    port map (
            O => \N__40872\,
            I => \N__40855\
        );

    \I__9029\ : CascadeMux
    port map (
            O => \N__40871\,
            I => \N__40851\
        );

    \I__9028\ : CascadeMux
    port map (
            O => \N__40870\,
            I => \N__40847\
        );

    \I__9027\ : CascadeMux
    port map (
            O => \N__40869\,
            I => \N__40843\
        );

    \I__9026\ : CascadeMux
    port map (
            O => \N__40868\,
            I => \N__40839\
        );

    \I__9025\ : CascadeMux
    port map (
            O => \N__40867\,
            I => \N__40834\
        );

    \I__9024\ : InMux
    port map (
            O => \N__40866\,
            I => \N__40818\
        );

    \I__9023\ : InMux
    port map (
            O => \N__40863\,
            I => \N__40818\
        );

    \I__9022\ : InMux
    port map (
            O => \N__40862\,
            I => \N__40818\
        );

    \I__9021\ : InMux
    port map (
            O => \N__40859\,
            I => \N__40818\
        );

    \I__9020\ : InMux
    port map (
            O => \N__40858\,
            I => \N__40818\
        );

    \I__9019\ : InMux
    port map (
            O => \N__40855\,
            I => \N__40818\
        );

    \I__9018\ : InMux
    port map (
            O => \N__40854\,
            I => \N__40818\
        );

    \I__9017\ : InMux
    port map (
            O => \N__40851\,
            I => \N__40801\
        );

    \I__9016\ : InMux
    port map (
            O => \N__40850\,
            I => \N__40801\
        );

    \I__9015\ : InMux
    port map (
            O => \N__40847\,
            I => \N__40801\
        );

    \I__9014\ : InMux
    port map (
            O => \N__40846\,
            I => \N__40801\
        );

    \I__9013\ : InMux
    port map (
            O => \N__40843\,
            I => \N__40801\
        );

    \I__9012\ : InMux
    port map (
            O => \N__40842\,
            I => \N__40801\
        );

    \I__9011\ : InMux
    port map (
            O => \N__40839\,
            I => \N__40801\
        );

    \I__9010\ : InMux
    port map (
            O => \N__40838\,
            I => \N__40801\
        );

    \I__9009\ : InMux
    port map (
            O => \N__40837\,
            I => \N__40794\
        );

    \I__9008\ : InMux
    port map (
            O => \N__40834\,
            I => \N__40794\
        );

    \I__9007\ : InMux
    port map (
            O => \N__40833\,
            I => \N__40794\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__40818\,
            I => \N__40787\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__40801\,
            I => \N__40787\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__40794\,
            I => \N__40787\
        );

    \I__9003\ : Span4Mux_v
    port map (
            O => \N__40787\,
            I => \N__40784\
        );

    \I__9002\ : Odrv4
    port map (
            O => \N__40784\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__9001\ : InMux
    port map (
            O => \N__40781\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__9000\ : InMux
    port map (
            O => \N__40778\,
            I => \N__40775\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__40775\,
            I => \N__40771\
        );

    \I__8998\ : InMux
    port map (
            O => \N__40774\,
            I => \N__40768\
        );

    \I__8997\ : Odrv4
    port map (
            O => \N__40771\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__40768\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__8995\ : CascadeMux
    port map (
            O => \N__40763\,
            I => \N__40760\
        );

    \I__8994\ : InMux
    port map (
            O => \N__40760\,
            I => \N__40756\
        );

    \I__8993\ : InMux
    port map (
            O => \N__40759\,
            I => \N__40753\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__40756\,
            I => \N__40750\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__40753\,
            I => \N__40744\
        );

    \I__8990\ : Span4Mux_v
    port map (
            O => \N__40750\,
            I => \N__40744\
        );

    \I__8989\ : InMux
    port map (
            O => \N__40749\,
            I => \N__40741\
        );

    \I__8988\ : Odrv4
    port map (
            O => \N__40744\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__40741\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__8986\ : CascadeMux
    port map (
            O => \N__40736\,
            I => \N__40732\
        );

    \I__8985\ : CascadeMux
    port map (
            O => \N__40735\,
            I => \N__40729\
        );

    \I__8984\ : InMux
    port map (
            O => \N__40732\,
            I => \N__40726\
        );

    \I__8983\ : InMux
    port map (
            O => \N__40729\,
            I => \N__40722\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__40726\,
            I => \N__40719\
        );

    \I__8981\ : CascadeMux
    port map (
            O => \N__40725\,
            I => \N__40716\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__40722\,
            I => \N__40713\
        );

    \I__8979\ : Span4Mux_h
    port map (
            O => \N__40719\,
            I => \N__40710\
        );

    \I__8978\ : InMux
    port map (
            O => \N__40716\,
            I => \N__40706\
        );

    \I__8977\ : Span4Mux_v
    port map (
            O => \N__40713\,
            I => \N__40703\
        );

    \I__8976\ : Sp12to4
    port map (
            O => \N__40710\,
            I => \N__40700\
        );

    \I__8975\ : InMux
    port map (
            O => \N__40709\,
            I => \N__40697\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__40706\,
            I => \N__40694\
        );

    \I__8973\ : Span4Mux_v
    port map (
            O => \N__40703\,
            I => \N__40691\
        );

    \I__8972\ : Span12Mux_v
    port map (
            O => \N__40700\,
            I => \N__40688\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__40697\,
            I => \N__40683\
        );

    \I__8970\ : Span4Mux_v
    port map (
            O => \N__40694\,
            I => \N__40683\
        );

    \I__8969\ : Odrv4
    port map (
            O => \N__40691\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__8968\ : Odrv12
    port map (
            O => \N__40688\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__8967\ : Odrv4
    port map (
            O => \N__40683\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__8966\ : InMux
    port map (
            O => \N__40676\,
            I => \bfn_15_25_0_\
        );

    \I__8965\ : InMux
    port map (
            O => \N__40673\,
            I => \N__40670\
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__40670\,
            I => \N__40666\
        );

    \I__8963\ : InMux
    port map (
            O => \N__40669\,
            I => \N__40662\
        );

    \I__8962\ : Span12Mux_s7_v
    port map (
            O => \N__40666\,
            I => \N__40658\
        );

    \I__8961\ : InMux
    port map (
            O => \N__40665\,
            I => \N__40655\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__40662\,
            I => \N__40652\
        );

    \I__8959\ : InMux
    port map (
            O => \N__40661\,
            I => \N__40649\
        );

    \I__8958\ : Span12Mux_h
    port map (
            O => \N__40658\,
            I => \N__40646\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__40655\,
            I => \N__40643\
        );

    \I__8956\ : Span4Mux_v
    port map (
            O => \N__40652\,
            I => \N__40640\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__40649\,
            I => \N__40637\
        );

    \I__8954\ : Odrv12
    port map (
            O => \N__40646\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__8953\ : Odrv4
    port map (
            O => \N__40643\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__8952\ : Odrv4
    port map (
            O => \N__40640\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__8951\ : Odrv4
    port map (
            O => \N__40637\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__8950\ : InMux
    port map (
            O => \N__40628\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__8949\ : CascadeMux
    port map (
            O => \N__40625\,
            I => \N__40622\
        );

    \I__8948\ : InMux
    port map (
            O => \N__40622\,
            I => \N__40619\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__40619\,
            I => \N__40616\
        );

    \I__8946\ : Span4Mux_v
    port map (
            O => \N__40616\,
            I => \N__40611\
        );

    \I__8945\ : InMux
    port map (
            O => \N__40615\,
            I => \N__40608\
        );

    \I__8944\ : InMux
    port map (
            O => \N__40614\,
            I => \N__40605\
        );

    \I__8943\ : Sp12to4
    port map (
            O => \N__40611\,
            I => \N__40599\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__40608\,
            I => \N__40599\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__40605\,
            I => \N__40596\
        );

    \I__8940\ : InMux
    port map (
            O => \N__40604\,
            I => \N__40593\
        );

    \I__8939\ : Span12Mux_h
    port map (
            O => \N__40599\,
            I => \N__40590\
        );

    \I__8938\ : Span4Mux_v
    port map (
            O => \N__40596\,
            I => \N__40587\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__40593\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__8936\ : Odrv12
    port map (
            O => \N__40590\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__8935\ : Odrv4
    port map (
            O => \N__40587\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__8934\ : InMux
    port map (
            O => \N__40580\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__8933\ : InMux
    port map (
            O => \N__40577\,
            I => \N__40574\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__40574\,
            I => \N__40570\
        );

    \I__8931\ : InMux
    port map (
            O => \N__40573\,
            I => \N__40567\
        );

    \I__8930\ : Span4Mux_v
    port map (
            O => \N__40570\,
            I => \N__40564\
        );

    \I__8929\ : LocalMux
    port map (
            O => \N__40567\,
            I => \N__40561\
        );

    \I__8928\ : Sp12to4
    port map (
            O => \N__40564\,
            I => \N__40557\
        );

    \I__8927\ : Span4Mux_h
    port map (
            O => \N__40561\,
            I => \N__40554\
        );

    \I__8926\ : InMux
    port map (
            O => \N__40560\,
            I => \N__40551\
        );

    \I__8925\ : Span12Mux_h
    port map (
            O => \N__40557\,
            I => \N__40543\
        );

    \I__8924\ : Sp12to4
    port map (
            O => \N__40554\,
            I => \N__40543\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__40551\,
            I => \N__40543\
        );

    \I__8922\ : InMux
    port map (
            O => \N__40550\,
            I => \N__40540\
        );

    \I__8921\ : Span12Mux_v
    port map (
            O => \N__40543\,
            I => \N__40537\
        );

    \I__8920\ : LocalMux
    port map (
            O => \N__40540\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__8919\ : Odrv12
    port map (
            O => \N__40537\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__8918\ : InMux
    port map (
            O => \N__40532\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__8917\ : CascadeMux
    port map (
            O => \N__40529\,
            I => \N__40525\
        );

    \I__8916\ : CascadeMux
    port map (
            O => \N__40528\,
            I => \N__40522\
        );

    \I__8915\ : InMux
    port map (
            O => \N__40525\,
            I => \N__40519\
        );

    \I__8914\ : InMux
    port map (
            O => \N__40522\,
            I => \N__40516\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__40519\,
            I => \N__40511\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__40516\,
            I => \N__40508\
        );

    \I__8911\ : InMux
    port map (
            O => \N__40515\,
            I => \N__40505\
        );

    \I__8910\ : InMux
    port map (
            O => \N__40514\,
            I => \N__40502\
        );

    \I__8909\ : Span4Mux_v
    port map (
            O => \N__40511\,
            I => \N__40499\
        );

    \I__8908\ : Span12Mux_h
    port map (
            O => \N__40508\,
            I => \N__40494\
        );

    \I__8907\ : LocalMux
    port map (
            O => \N__40505\,
            I => \N__40494\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__40502\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__8905\ : Odrv4
    port map (
            O => \N__40499\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__8904\ : Odrv12
    port map (
            O => \N__40494\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__8903\ : InMux
    port map (
            O => \N__40487\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__8902\ : InMux
    port map (
            O => \N__40484\,
            I => \N__40481\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__40481\,
            I => \N__40478\
        );

    \I__8900\ : Sp12to4
    port map (
            O => \N__40478\,
            I => \N__40474\
        );

    \I__8899\ : InMux
    port map (
            O => \N__40477\,
            I => \N__40470\
        );

    \I__8898\ : Span12Mux_v
    port map (
            O => \N__40474\,
            I => \N__40466\
        );

    \I__8897\ : InMux
    port map (
            O => \N__40473\,
            I => \N__40463\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__40470\,
            I => \N__40460\
        );

    \I__8895\ : InMux
    port map (
            O => \N__40469\,
            I => \N__40457\
        );

    \I__8894\ : Span12Mux_h
    port map (
            O => \N__40466\,
            I => \N__40454\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__40463\,
            I => \N__40451\
        );

    \I__8892\ : Span4Mux_v
    port map (
            O => \N__40460\,
            I => \N__40448\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__40457\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__8890\ : Odrv12
    port map (
            O => \N__40454\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__8889\ : Odrv12
    port map (
            O => \N__40451\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__8888\ : Odrv4
    port map (
            O => \N__40448\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__8887\ : InMux
    port map (
            O => \N__40439\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__8886\ : CascadeMux
    port map (
            O => \N__40436\,
            I => \N__40433\
        );

    \I__8885\ : InMux
    port map (
            O => \N__40433\,
            I => \N__40430\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__40430\,
            I => \N__40427\
        );

    \I__8883\ : Span4Mux_v
    port map (
            O => \N__40427\,
            I => \N__40424\
        );

    \I__8882\ : Span4Mux_h
    port map (
            O => \N__40424\,
            I => \N__40421\
        );

    \I__8881\ : Span4Mux_h
    port map (
            O => \N__40421\,
            I => \N__40417\
        );

    \I__8880\ : InMux
    port map (
            O => \N__40420\,
            I => \N__40414\
        );

    \I__8879\ : Span4Mux_h
    port map (
            O => \N__40417\,
            I => \N__40407\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__40414\,
            I => \N__40407\
        );

    \I__8877\ : InMux
    port map (
            O => \N__40413\,
            I => \N__40404\
        );

    \I__8876\ : InMux
    port map (
            O => \N__40412\,
            I => \N__40401\
        );

    \I__8875\ : Span4Mux_v
    port map (
            O => \N__40407\,
            I => \N__40396\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__40404\,
            I => \N__40396\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__40401\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__8872\ : Odrv4
    port map (
            O => \N__40396\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__8871\ : InMux
    port map (
            O => \N__40391\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__8870\ : InMux
    port map (
            O => \N__40388\,
            I => \N__40385\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__40385\,
            I => \N__40380\
        );

    \I__8868\ : InMux
    port map (
            O => \N__40384\,
            I => \N__40376\
        );

    \I__8867\ : InMux
    port map (
            O => \N__40383\,
            I => \N__40373\
        );

    \I__8866\ : Sp12to4
    port map (
            O => \N__40380\,
            I => \N__40370\
        );

    \I__8865\ : CascadeMux
    port map (
            O => \N__40379\,
            I => \N__40367\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__40376\,
            I => \N__40362\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__40373\,
            I => \N__40362\
        );

    \I__8862\ : Span12Mux_v
    port map (
            O => \N__40370\,
            I => \N__40359\
        );

    \I__8861\ : InMux
    port map (
            O => \N__40367\,
            I => \N__40356\
        );

    \I__8860\ : Span4Mux_v
    port map (
            O => \N__40362\,
            I => \N__40353\
        );

    \I__8859\ : Odrv12
    port map (
            O => \N__40359\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__40356\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__8857\ : Odrv4
    port map (
            O => \N__40353\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__8856\ : InMux
    port map (
            O => \N__40346\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\
        );

    \I__8855\ : InMux
    port map (
            O => \N__40343\,
            I => \N__40340\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__40340\,
            I => \N__40337\
        );

    \I__8853\ : Odrv4
    port map (
            O => \N__40337\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__8852\ : CascadeMux
    port map (
            O => \N__40334\,
            I => \N__40331\
        );

    \I__8851\ : InMux
    port map (
            O => \N__40331\,
            I => \N__40328\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__40328\,
            I => \N__40324\
        );

    \I__8849\ : InMux
    port map (
            O => \N__40327\,
            I => \N__40320\
        );

    \I__8848\ : Span4Mux_v
    port map (
            O => \N__40324\,
            I => \N__40317\
        );

    \I__8847\ : InMux
    port map (
            O => \N__40323\,
            I => \N__40314\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__40320\,
            I => \N__40311\
        );

    \I__8845\ : Span4Mux_h
    port map (
            O => \N__40317\,
            I => \N__40308\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__40314\,
            I => \N__40303\
        );

    \I__8843\ : Span4Mux_v
    port map (
            O => \N__40311\,
            I => \N__40303\
        );

    \I__8842\ : Sp12to4
    port map (
            O => \N__40308\,
            I => \N__40299\
        );

    \I__8841\ : Span4Mux_v
    port map (
            O => \N__40303\,
            I => \N__40296\
        );

    \I__8840\ : InMux
    port map (
            O => \N__40302\,
            I => \N__40293\
        );

    \I__8839\ : Span12Mux_h
    port map (
            O => \N__40299\,
            I => \N__40290\
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__40296\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__40293\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__8836\ : Odrv12
    port map (
            O => \N__40290\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__8835\ : InMux
    port map (
            O => \N__40283\,
            I => \bfn_15_24_0_\
        );

    \I__8834\ : InMux
    port map (
            O => \N__40280\,
            I => \N__40277\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__40277\,
            I => \N__40274\
        );

    \I__8832\ : Odrv12
    port map (
            O => \N__40274\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__8831\ : CascadeMux
    port map (
            O => \N__40271\,
            I => \N__40268\
        );

    \I__8830\ : InMux
    port map (
            O => \N__40268\,
            I => \N__40265\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__40265\,
            I => \N__40262\
        );

    \I__8828\ : Span4Mux_v
    port map (
            O => \N__40262\,
            I => \N__40258\
        );

    \I__8827\ : CascadeMux
    port map (
            O => \N__40261\,
            I => \N__40255\
        );

    \I__8826\ : Span4Mux_v
    port map (
            O => \N__40258\,
            I => \N__40251\
        );

    \I__8825\ : InMux
    port map (
            O => \N__40255\,
            I => \N__40247\
        );

    \I__8824\ : InMux
    port map (
            O => \N__40254\,
            I => \N__40244\
        );

    \I__8823\ : Span4Mux_v
    port map (
            O => \N__40251\,
            I => \N__40241\
        );

    \I__8822\ : InMux
    port map (
            O => \N__40250\,
            I => \N__40238\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__40247\,
            I => \N__40235\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__40244\,
            I => \N__40232\
        );

    \I__8819\ : Sp12to4
    port map (
            O => \N__40241\,
            I => \N__40229\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__40238\,
            I => \N__40222\
        );

    \I__8817\ : Span4Mux_v
    port map (
            O => \N__40235\,
            I => \N__40222\
        );

    \I__8816\ : Span4Mux_h
    port map (
            O => \N__40232\,
            I => \N__40222\
        );

    \I__8815\ : Odrv12
    port map (
            O => \N__40229\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__8814\ : Odrv4
    port map (
            O => \N__40222\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__8813\ : InMux
    port map (
            O => \N__40217\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__8812\ : InMux
    port map (
            O => \N__40214\,
            I => \N__40211\
        );

    \I__8811\ : LocalMux
    port map (
            O => \N__40211\,
            I => \N__40208\
        );

    \I__8810\ : Span12Mux_h
    port map (
            O => \N__40208\,
            I => \N__40205\
        );

    \I__8809\ : Odrv12
    port map (
            O => \N__40205\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__8808\ : CascadeMux
    port map (
            O => \N__40202\,
            I => \N__40199\
        );

    \I__8807\ : InMux
    port map (
            O => \N__40199\,
            I => \N__40195\
        );

    \I__8806\ : CascadeMux
    port map (
            O => \N__40198\,
            I => \N__40191\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__40195\,
            I => \N__40188\
        );

    \I__8804\ : InMux
    port map (
            O => \N__40194\,
            I => \N__40185\
        );

    \I__8803\ : InMux
    port map (
            O => \N__40191\,
            I => \N__40182\
        );

    \I__8802\ : Sp12to4
    port map (
            O => \N__40188\,
            I => \N__40178\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__40185\,
            I => \N__40175\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__40182\,
            I => \N__40172\
        );

    \I__8799\ : InMux
    port map (
            O => \N__40181\,
            I => \N__40169\
        );

    \I__8798\ : Span12Mux_h
    port map (
            O => \N__40178\,
            I => \N__40166\
        );

    \I__8797\ : Span4Mux_v
    port map (
            O => \N__40175\,
            I => \N__40161\
        );

    \I__8796\ : Span4Mux_v
    port map (
            O => \N__40172\,
            I => \N__40161\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__40169\,
            I => \N__40158\
        );

    \I__8794\ : Odrv12
    port map (
            O => \N__40166\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__8793\ : Odrv4
    port map (
            O => \N__40161\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__8792\ : Odrv4
    port map (
            O => \N__40158\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__8791\ : InMux
    port map (
            O => \N__40151\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__8790\ : InMux
    port map (
            O => \N__40148\,
            I => \N__40145\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__40145\,
            I => \N__40142\
        );

    \I__8788\ : Sp12to4
    port map (
            O => \N__40142\,
            I => \N__40139\
        );

    \I__8787\ : Odrv12
    port map (
            O => \N__40139\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__8786\ : CascadeMux
    port map (
            O => \N__40136\,
            I => \N__40133\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40133\,
            I => \N__40130\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__40130\,
            I => \N__40125\
        );

    \I__8783\ : InMux
    port map (
            O => \N__40129\,
            I => \N__40122\
        );

    \I__8782\ : InMux
    port map (
            O => \N__40128\,
            I => \N__40119\
        );

    \I__8781\ : Span4Mux_v
    port map (
            O => \N__40125\,
            I => \N__40115\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__40122\,
            I => \N__40112\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__40119\,
            I => \N__40109\
        );

    \I__8778\ : CascadeMux
    port map (
            O => \N__40118\,
            I => \N__40106\
        );

    \I__8777\ : Sp12to4
    port map (
            O => \N__40115\,
            I => \N__40103\
        );

    \I__8776\ : Span4Mux_v
    port map (
            O => \N__40112\,
            I => \N__40098\
        );

    \I__8775\ : Span4Mux_v
    port map (
            O => \N__40109\,
            I => \N__40098\
        );

    \I__8774\ : InMux
    port map (
            O => \N__40106\,
            I => \N__40095\
        );

    \I__8773\ : Span12Mux_h
    port map (
            O => \N__40103\,
            I => \N__40092\
        );

    \I__8772\ : Odrv4
    port map (
            O => \N__40098\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__40095\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__8770\ : Odrv12
    port map (
            O => \N__40092\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__8769\ : InMux
    port map (
            O => \N__40085\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__8768\ : InMux
    port map (
            O => \N__40082\,
            I => \N__40077\
        );

    \I__8767\ : CascadeMux
    port map (
            O => \N__40081\,
            I => \N__40074\
        );

    \I__8766\ : InMux
    port map (
            O => \N__40080\,
            I => \N__40071\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__40077\,
            I => \N__40068\
        );

    \I__8764\ : InMux
    port map (
            O => \N__40074\,
            I => \N__40064\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__40071\,
            I => \N__40061\
        );

    \I__8762\ : Span12Mux_v
    port map (
            O => \N__40068\,
            I => \N__40058\
        );

    \I__8761\ : InMux
    port map (
            O => \N__40067\,
            I => \N__40055\
        );

    \I__8760\ : LocalMux
    port map (
            O => \N__40064\,
            I => \N__40050\
        );

    \I__8759\ : Span4Mux_v
    port map (
            O => \N__40061\,
            I => \N__40050\
        );

    \I__8758\ : Odrv12
    port map (
            O => \N__40058\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__40055\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__8756\ : Odrv4
    port map (
            O => \N__40050\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__8755\ : CascadeMux
    port map (
            O => \N__40043\,
            I => \N__40040\
        );

    \I__8754\ : InMux
    port map (
            O => \N__40040\,
            I => \N__40037\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__40037\,
            I => \N__40034\
        );

    \I__8752\ : Odrv12
    port map (
            O => \N__40034\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__8751\ : InMux
    port map (
            O => \N__40031\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__8750\ : CascadeMux
    port map (
            O => \N__40028\,
            I => \N__40025\
        );

    \I__8749\ : InMux
    port map (
            O => \N__40025\,
            I => \N__40022\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__40022\,
            I => \N__40017\
        );

    \I__8747\ : InMux
    port map (
            O => \N__40021\,
            I => \N__40013\
        );

    \I__8746\ : InMux
    port map (
            O => \N__40020\,
            I => \N__40010\
        );

    \I__8745\ : Sp12to4
    port map (
            O => \N__40017\,
            I => \N__40007\
        );

    \I__8744\ : InMux
    port map (
            O => \N__40016\,
            I => \N__40004\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__40013\,
            I => \N__40001\
        );

    \I__8742\ : LocalMux
    port map (
            O => \N__40010\,
            I => \N__39994\
        );

    \I__8741\ : Span12Mux_h
    port map (
            O => \N__40007\,
            I => \N__39994\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__40004\,
            I => \N__39994\
        );

    \I__8739\ : Span4Mux_v
    port map (
            O => \N__40001\,
            I => \N__39991\
        );

    \I__8738\ : Odrv12
    port map (
            O => \N__39994\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__8737\ : Odrv4
    port map (
            O => \N__39991\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__8736\ : InMux
    port map (
            O => \N__39986\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__8735\ : InMux
    port map (
            O => \N__39983\,
            I => \N__39980\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__39980\,
            I => \N__39976\
        );

    \I__8733\ : InMux
    port map (
            O => \N__39979\,
            I => \N__39973\
        );

    \I__8732\ : Sp12to4
    port map (
            O => \N__39976\,
            I => \N__39970\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__39973\,
            I => \N__39967\
        );

    \I__8730\ : Span12Mux_v
    port map (
            O => \N__39970\,
            I => \N__39962\
        );

    \I__8729\ : Span4Mux_h
    port map (
            O => \N__39967\,
            I => \N__39959\
        );

    \I__8728\ : InMux
    port map (
            O => \N__39966\,
            I => \N__39956\
        );

    \I__8727\ : InMux
    port map (
            O => \N__39965\,
            I => \N__39953\
        );

    \I__8726\ : Span12Mux_h
    port map (
            O => \N__39962\,
            I => \N__39946\
        );

    \I__8725\ : Sp12to4
    port map (
            O => \N__39959\,
            I => \N__39946\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__39956\,
            I => \N__39946\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__39953\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__8722\ : Odrv12
    port map (
            O => \N__39946\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__8721\ : InMux
    port map (
            O => \N__39941\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__8720\ : CascadeMux
    port map (
            O => \N__39938\,
            I => \N__39935\
        );

    \I__8719\ : InMux
    port map (
            O => \N__39935\,
            I => \N__39932\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__39932\,
            I => \N__39929\
        );

    \I__8717\ : Span4Mux_v
    port map (
            O => \N__39929\,
            I => \N__39926\
        );

    \I__8716\ : Span4Mux_h
    port map (
            O => \N__39926\,
            I => \N__39922\
        );

    \I__8715\ : InMux
    port map (
            O => \N__39925\,
            I => \N__39917\
        );

    \I__8714\ : Sp12to4
    port map (
            O => \N__39922\,
            I => \N__39914\
        );

    \I__8713\ : InMux
    port map (
            O => \N__39921\,
            I => \N__39911\
        );

    \I__8712\ : InMux
    port map (
            O => \N__39920\,
            I => \N__39908\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__39917\,
            I => \N__39901\
        );

    \I__8710\ : Span12Mux_h
    port map (
            O => \N__39914\,
            I => \N__39901\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__39911\,
            I => \N__39901\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__39908\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__8707\ : Odrv12
    port map (
            O => \N__39901\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__8706\ : InMux
    port map (
            O => \N__39896\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\
        );

    \I__8705\ : InMux
    port map (
            O => \N__39893\,
            I => \N__39889\
        );

    \I__8704\ : InMux
    port map (
            O => \N__39892\,
            I => \N__39886\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__39889\,
            I => \N__39881\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__39886\,
            I => \N__39881\
        );

    \I__8701\ : Odrv12
    port map (
            O => \N__39881\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__8700\ : CascadeMux
    port map (
            O => \N__39878\,
            I => \N__39874\
        );

    \I__8699\ : CascadeMux
    port map (
            O => \N__39877\,
            I => \N__39870\
        );

    \I__8698\ : InMux
    port map (
            O => \N__39874\,
            I => \N__39867\
        );

    \I__8697\ : InMux
    port map (
            O => \N__39873\,
            I => \N__39864\
        );

    \I__8696\ : InMux
    port map (
            O => \N__39870\,
            I => \N__39861\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__39867\,
            I => \N__39858\
        );

    \I__8694\ : LocalMux
    port map (
            O => \N__39864\,
            I => \N__39854\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__39861\,
            I => \N__39851\
        );

    \I__8692\ : Span4Mux_v
    port map (
            O => \N__39858\,
            I => \N__39848\
        );

    \I__8691\ : CascadeMux
    port map (
            O => \N__39857\,
            I => \N__39845\
        );

    \I__8690\ : Span4Mux_v
    port map (
            O => \N__39854\,
            I => \N__39842\
        );

    \I__8689\ : Span4Mux_v
    port map (
            O => \N__39851\,
            I => \N__39839\
        );

    \I__8688\ : Span4Mux_h
    port map (
            O => \N__39848\,
            I => \N__39836\
        );

    \I__8687\ : InMux
    port map (
            O => \N__39845\,
            I => \N__39832\
        );

    \I__8686\ : Sp12to4
    port map (
            O => \N__39842\,
            I => \N__39825\
        );

    \I__8685\ : Sp12to4
    port map (
            O => \N__39839\,
            I => \N__39825\
        );

    \I__8684\ : Sp12to4
    port map (
            O => \N__39836\,
            I => \N__39825\
        );

    \I__8683\ : InMux
    port map (
            O => \N__39835\,
            I => \N__39822\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__39832\,
            I => \N__39819\
        );

    \I__8681\ : Span12Mux_h
    port map (
            O => \N__39825\,
            I => \N__39816\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__39822\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__8679\ : Odrv4
    port map (
            O => \N__39819\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__8678\ : Odrv12
    port map (
            O => \N__39816\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__8677\ : InMux
    port map (
            O => \N__39809\,
            I => \N__39806\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__39806\,
            I => \N__39803\
        );

    \I__8675\ : Odrv12
    port map (
            O => \N__39803\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__8674\ : CascadeMux
    port map (
            O => \N__39800\,
            I => \N__39797\
        );

    \I__8673\ : InMux
    port map (
            O => \N__39797\,
            I => \N__39793\
        );

    \I__8672\ : InMux
    port map (
            O => \N__39796\,
            I => \N__39790\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__39793\,
            I => \N__39787\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__39790\,
            I => \N__39781\
        );

    \I__8669\ : Span12Mux_h
    port map (
            O => \N__39787\,
            I => \N__39781\
        );

    \I__8668\ : InMux
    port map (
            O => \N__39786\,
            I => \N__39778\
        );

    \I__8667\ : Odrv12
    port map (
            O => \N__39781\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__39778\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__8665\ : InMux
    port map (
            O => \N__39773\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__8664\ : InMux
    port map (
            O => \N__39770\,
            I => \N__39767\
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__39767\,
            I => \N__39764\
        );

    \I__8662\ : Span4Mux_v
    port map (
            O => \N__39764\,
            I => \N__39761\
        );

    \I__8661\ : Odrv4
    port map (
            O => \N__39761\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__8660\ : CascadeMux
    port map (
            O => \N__39758\,
            I => \N__39755\
        );

    \I__8659\ : InMux
    port map (
            O => \N__39755\,
            I => \N__39752\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__39752\,
            I => \N__39749\
        );

    \I__8657\ : Span4Mux_v
    port map (
            O => \N__39749\,
            I => \N__39744\
        );

    \I__8656\ : InMux
    port map (
            O => \N__39748\,
            I => \N__39741\
        );

    \I__8655\ : InMux
    port map (
            O => \N__39747\,
            I => \N__39738\
        );

    \I__8654\ : Span4Mux_h
    port map (
            O => \N__39744\,
            I => \N__39735\
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__39741\,
            I => \N__39730\
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__39738\,
            I => \N__39730\
        );

    \I__8651\ : Sp12to4
    port map (
            O => \N__39735\,
            I => \N__39726\
        );

    \I__8650\ : Span12Mux_v
    port map (
            O => \N__39730\,
            I => \N__39723\
        );

    \I__8649\ : InMux
    port map (
            O => \N__39729\,
            I => \N__39720\
        );

    \I__8648\ : Span12Mux_v
    port map (
            O => \N__39726\,
            I => \N__39717\
        );

    \I__8647\ : Odrv12
    port map (
            O => \N__39723\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__39720\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__8645\ : Odrv12
    port map (
            O => \N__39717\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__8644\ : InMux
    port map (
            O => \N__39710\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__8643\ : InMux
    port map (
            O => \N__39707\,
            I => \N__39704\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__39704\,
            I => \N__39701\
        );

    \I__8641\ : Span4Mux_h
    port map (
            O => \N__39701\,
            I => \N__39698\
        );

    \I__8640\ : Odrv4
    port map (
            O => \N__39698\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__8639\ : CascadeMux
    port map (
            O => \N__39695\,
            I => \N__39691\
        );

    \I__8638\ : InMux
    port map (
            O => \N__39694\,
            I => \N__39687\
        );

    \I__8637\ : InMux
    port map (
            O => \N__39691\,
            I => \N__39684\
        );

    \I__8636\ : InMux
    port map (
            O => \N__39690\,
            I => \N__39681\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__39687\,
            I => \N__39678\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__39684\,
            I => \N__39675\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__39681\,
            I => \N__39670\
        );

    \I__8632\ : Span4Mux_v
    port map (
            O => \N__39678\,
            I => \N__39670\
        );

    \I__8631\ : Span4Mux_v
    port map (
            O => \N__39675\,
            I => \N__39667\
        );

    \I__8630\ : Sp12to4
    port map (
            O => \N__39670\,
            I => \N__39661\
        );

    \I__8629\ : Sp12to4
    port map (
            O => \N__39667\,
            I => \N__39661\
        );

    \I__8628\ : InMux
    port map (
            O => \N__39666\,
            I => \N__39658\
        );

    \I__8627\ : Span12Mux_h
    port map (
            O => \N__39661\,
            I => \N__39655\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__39658\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__8625\ : Odrv12
    port map (
            O => \N__39655\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__8624\ : InMux
    port map (
            O => \N__39650\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__8623\ : InMux
    port map (
            O => \N__39647\,
            I => \N__39642\
        );

    \I__8622\ : InMux
    port map (
            O => \N__39646\,
            I => \N__39639\
        );

    \I__8621\ : InMux
    port map (
            O => \N__39645\,
            I => \N__39635\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__39642\,
            I => \N__39632\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__39639\,
            I => \N__39629\
        );

    \I__8618\ : InMux
    port map (
            O => \N__39638\,
            I => \N__39626\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__39635\,
            I => \N__39621\
        );

    \I__8616\ : Span4Mux_v
    port map (
            O => \N__39632\,
            I => \N__39621\
        );

    \I__8615\ : Span12Mux_v
    port map (
            O => \N__39629\,
            I => \N__39618\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__39626\,
            I => \N__39615\
        );

    \I__8613\ : Span4Mux_v
    port map (
            O => \N__39621\,
            I => \N__39612\
        );

    \I__8612\ : Odrv12
    port map (
            O => \N__39618\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__8611\ : Odrv4
    port map (
            O => \N__39615\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__8610\ : Odrv4
    port map (
            O => \N__39612\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__8609\ : CascadeMux
    port map (
            O => \N__39605\,
            I => \N__39602\
        );

    \I__8608\ : InMux
    port map (
            O => \N__39602\,
            I => \N__39599\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__39599\,
            I => \N__39596\
        );

    \I__8606\ : Odrv4
    port map (
            O => \N__39596\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__8605\ : InMux
    port map (
            O => \N__39593\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__8604\ : InMux
    port map (
            O => \N__39590\,
            I => \N__39587\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__39587\,
            I => \N__39584\
        );

    \I__8602\ : Odrv4
    port map (
            O => \N__39584\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__8601\ : CascadeMux
    port map (
            O => \N__39581\,
            I => \N__39577\
        );

    \I__8600\ : CascadeMux
    port map (
            O => \N__39580\,
            I => \N__39574\
        );

    \I__8599\ : InMux
    port map (
            O => \N__39577\,
            I => \N__39570\
        );

    \I__8598\ : InMux
    port map (
            O => \N__39574\,
            I => \N__39567\
        );

    \I__8597\ : InMux
    port map (
            O => \N__39573\,
            I => \N__39564\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__39570\,
            I => \N__39561\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__39567\,
            I => \N__39558\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__39564\,
            I => \N__39550\
        );

    \I__8593\ : Sp12to4
    port map (
            O => \N__39561\,
            I => \N__39550\
        );

    \I__8592\ : Span12Mux_h
    port map (
            O => \N__39558\,
            I => \N__39550\
        );

    \I__8591\ : InMux
    port map (
            O => \N__39557\,
            I => \N__39547\
        );

    \I__8590\ : Odrv12
    port map (
            O => \N__39550\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__39547\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__8588\ : InMux
    port map (
            O => \N__39542\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__8587\ : InMux
    port map (
            O => \N__39539\,
            I => \N__39536\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__39536\,
            I => \N__39533\
        );

    \I__8585\ : Odrv12
    port map (
            O => \N__39533\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__8584\ : CascadeMux
    port map (
            O => \N__39530\,
            I => \N__39527\
        );

    \I__8583\ : InMux
    port map (
            O => \N__39527\,
            I => \N__39524\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__39524\,
            I => \N__39520\
        );

    \I__8581\ : InMux
    port map (
            O => \N__39523\,
            I => \N__39516\
        );

    \I__8580\ : Sp12to4
    port map (
            O => \N__39520\,
            I => \N__39513\
        );

    \I__8579\ : InMux
    port map (
            O => \N__39519\,
            I => \N__39509\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__39516\,
            I => \N__39506\
        );

    \I__8577\ : Span12Mux_v
    port map (
            O => \N__39513\,
            I => \N__39503\
        );

    \I__8576\ : InMux
    port map (
            O => \N__39512\,
            I => \N__39500\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__39509\,
            I => \N__39495\
        );

    \I__8574\ : Span12Mux_s11_v
    port map (
            O => \N__39506\,
            I => \N__39495\
        );

    \I__8573\ : Odrv12
    port map (
            O => \N__39503\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__39500\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__8571\ : Odrv12
    port map (
            O => \N__39495\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__8570\ : InMux
    port map (
            O => \N__39488\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__8569\ : InMux
    port map (
            O => \N__39485\,
            I => \N__39482\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__39482\,
            I => \N__39479\
        );

    \I__8567\ : Odrv4
    port map (
            O => \N__39479\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__8566\ : CascadeMux
    port map (
            O => \N__39476\,
            I => \N__39473\
        );

    \I__8565\ : InMux
    port map (
            O => \N__39473\,
            I => \N__39468\
        );

    \I__8564\ : InMux
    port map (
            O => \N__39472\,
            I => \N__39465\
        );

    \I__8563\ : InMux
    port map (
            O => \N__39471\,
            I => \N__39462\
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__39468\,
            I => \N__39459\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__39465\,
            I => \N__39453\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__39462\,
            I => \N__39453\
        );

    \I__8559\ : Span12Mux_v
    port map (
            O => \N__39459\,
            I => \N__39450\
        );

    \I__8558\ : InMux
    port map (
            O => \N__39458\,
            I => \N__39447\
        );

    \I__8557\ : Span12Mux_v
    port map (
            O => \N__39453\,
            I => \N__39444\
        );

    \I__8556\ : Odrv12
    port map (
            O => \N__39450\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__39447\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__8554\ : Odrv12
    port map (
            O => \N__39444\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__8553\ : InMux
    port map (
            O => \N__39437\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\
        );

    \I__8552\ : InMux
    port map (
            O => \N__39434\,
            I => \N__39430\
        );

    \I__8551\ : InMux
    port map (
            O => \N__39433\,
            I => \N__39427\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__39430\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__39427\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__8548\ : CascadeMux
    port map (
            O => \N__39422\,
            I => \N__39419\
        );

    \I__8547\ : InMux
    port map (
            O => \N__39419\,
            I => \N__39414\
        );

    \I__8546\ : InMux
    port map (
            O => \N__39418\,
            I => \N__39411\
        );

    \I__8545\ : InMux
    port map (
            O => \N__39417\,
            I => \N__39408\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__39414\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__39411\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__39408\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__8541\ : InMux
    port map (
            O => \N__39401\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__8540\ : InMux
    port map (
            O => \N__39398\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__8539\ : InMux
    port map (
            O => \N__39395\,
            I => \N__39392\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__39392\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__8537\ : InMux
    port map (
            O => \N__39389\,
            I => \N__39385\
        );

    \I__8536\ : InMux
    port map (
            O => \N__39388\,
            I => \N__39382\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__39385\,
            I => \N__39379\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__39382\,
            I => \N__39376\
        );

    \I__8533\ : Span4Mux_s3_h
    port map (
            O => \N__39379\,
            I => \N__39373\
        );

    \I__8532\ : Span12Mux_h
    port map (
            O => \N__39376\,
            I => \N__39370\
        );

    \I__8531\ : Span4Mux_h
    port map (
            O => \N__39373\,
            I => \N__39367\
        );

    \I__8530\ : Odrv12
    port map (
            O => \N__39370\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__8529\ : Odrv4
    port map (
            O => \N__39367\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__8528\ : IoInMux
    port map (
            O => \N__39362\,
            I => \N__39359\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__39359\,
            I => \N__39356\
        );

    \I__8526\ : IoSpan4Mux
    port map (
            O => \N__39356\,
            I => \N__39353\
        );

    \I__8525\ : Sp12to4
    port map (
            O => \N__39353\,
            I => \N__39348\
        );

    \I__8524\ : InMux
    port map (
            O => \N__39352\,
            I => \N__39345\
        );

    \I__8523\ : InMux
    port map (
            O => \N__39351\,
            I => \N__39342\
        );

    \I__8522\ : Odrv12
    port map (
            O => \N__39348\,
            I => s1_phy_c
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__39345\,
            I => s1_phy_c
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__39342\,
            I => s1_phy_c
        );

    \I__8519\ : InMux
    port map (
            O => \N__39335\,
            I => \N__39329\
        );

    \I__8518\ : InMux
    port map (
            O => \N__39334\,
            I => \N__39324\
        );

    \I__8517\ : InMux
    port map (
            O => \N__39333\,
            I => \N__39324\
        );

    \I__8516\ : InMux
    port map (
            O => \N__39332\,
            I => \N__39321\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__39329\,
            I => \N__39318\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__39324\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__39321\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__8512\ : Odrv4
    port map (
            O => \N__39318\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__8511\ : InMux
    port map (
            O => \N__39311\,
            I => \N__39303\
        );

    \I__8510\ : InMux
    port map (
            O => \N__39310\,
            I => \N__39300\
        );

    \I__8509\ : InMux
    port map (
            O => \N__39309\,
            I => \N__39295\
        );

    \I__8508\ : InMux
    port map (
            O => \N__39308\,
            I => \N__39295\
        );

    \I__8507\ : InMux
    port map (
            O => \N__39307\,
            I => \N__39289\
        );

    \I__8506\ : InMux
    port map (
            O => \N__39306\,
            I => \N__39289\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__39303\,
            I => \N__39282\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__39300\,
            I => \N__39282\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__39295\,
            I => \N__39282\
        );

    \I__8502\ : InMux
    port map (
            O => \N__39294\,
            I => \N__39279\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__39289\,
            I => state_3
        );

    \I__8500\ : Odrv4
    port map (
            O => \N__39282\,
            I => state_3
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__39279\,
            I => state_3
        );

    \I__8498\ : IoInMux
    port map (
            O => \N__39272\,
            I => \N__39269\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__39269\,
            I => \N__39266\
        );

    \I__8496\ : Span4Mux_s1_v
    port map (
            O => \N__39266\,
            I => \N__39263\
        );

    \I__8495\ : Span4Mux_h
    port map (
            O => \N__39263\,
            I => \N__39260\
        );

    \I__8494\ : Span4Mux_v
    port map (
            O => \N__39260\,
            I => \N__39256\
        );

    \I__8493\ : InMux
    port map (
            O => \N__39259\,
            I => \N__39253\
        );

    \I__8492\ : Odrv4
    port map (
            O => \N__39256\,
            I => \T01_c\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__39253\,
            I => \T01_c\
        );

    \I__8490\ : CascadeMux
    port map (
            O => \N__39248\,
            I => \N__39245\
        );

    \I__8489\ : InMux
    port map (
            O => \N__39245\,
            I => \N__39240\
        );

    \I__8488\ : InMux
    port map (
            O => \N__39244\,
            I => \N__39237\
        );

    \I__8487\ : InMux
    port map (
            O => \N__39243\,
            I => \N__39234\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__39240\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__39237\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__39234\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__8483\ : InMux
    port map (
            O => \N__39227\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__8482\ : CascadeMux
    port map (
            O => \N__39224\,
            I => \N__39221\
        );

    \I__8481\ : InMux
    port map (
            O => \N__39221\,
            I => \N__39216\
        );

    \I__8480\ : InMux
    port map (
            O => \N__39220\,
            I => \N__39213\
        );

    \I__8479\ : InMux
    port map (
            O => \N__39219\,
            I => \N__39210\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__39216\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__39213\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__39210\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__8475\ : InMux
    port map (
            O => \N__39203\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__8474\ : CascadeMux
    port map (
            O => \N__39200\,
            I => \N__39197\
        );

    \I__8473\ : InMux
    port map (
            O => \N__39197\,
            I => \N__39192\
        );

    \I__8472\ : InMux
    port map (
            O => \N__39196\,
            I => \N__39189\
        );

    \I__8471\ : InMux
    port map (
            O => \N__39195\,
            I => \N__39186\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__39192\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__39189\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__39186\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39179\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__8466\ : CascadeMux
    port map (
            O => \N__39176\,
            I => \N__39173\
        );

    \I__8465\ : InMux
    port map (
            O => \N__39173\,
            I => \N__39168\
        );

    \I__8464\ : InMux
    port map (
            O => \N__39172\,
            I => \N__39165\
        );

    \I__8463\ : InMux
    port map (
            O => \N__39171\,
            I => \N__39162\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__39168\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__39165\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__39162\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__8459\ : InMux
    port map (
            O => \N__39155\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__8458\ : CascadeMux
    port map (
            O => \N__39152\,
            I => \N__39149\
        );

    \I__8457\ : InMux
    port map (
            O => \N__39149\,
            I => \N__39144\
        );

    \I__8456\ : InMux
    port map (
            O => \N__39148\,
            I => \N__39141\
        );

    \I__8455\ : InMux
    port map (
            O => \N__39147\,
            I => \N__39138\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__39144\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__39141\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__39138\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__8451\ : InMux
    port map (
            O => \N__39131\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__8450\ : CascadeMux
    port map (
            O => \N__39128\,
            I => \N__39125\
        );

    \I__8449\ : InMux
    port map (
            O => \N__39125\,
            I => \N__39120\
        );

    \I__8448\ : InMux
    port map (
            O => \N__39124\,
            I => \N__39117\
        );

    \I__8447\ : InMux
    port map (
            O => \N__39123\,
            I => \N__39114\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__39120\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__39117\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__39114\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__8443\ : InMux
    port map (
            O => \N__39107\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__8442\ : CascadeMux
    port map (
            O => \N__39104\,
            I => \N__39101\
        );

    \I__8441\ : InMux
    port map (
            O => \N__39101\,
            I => \N__39096\
        );

    \I__8440\ : InMux
    port map (
            O => \N__39100\,
            I => \N__39093\
        );

    \I__8439\ : InMux
    port map (
            O => \N__39099\,
            I => \N__39090\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__39096\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__39093\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__39090\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__8435\ : InMux
    port map (
            O => \N__39083\,
            I => \bfn_15_17_0_\
        );

    \I__8434\ : CascadeMux
    port map (
            O => \N__39080\,
            I => \N__39077\
        );

    \I__8433\ : InMux
    port map (
            O => \N__39077\,
            I => \N__39072\
        );

    \I__8432\ : InMux
    port map (
            O => \N__39076\,
            I => \N__39069\
        );

    \I__8431\ : InMux
    port map (
            O => \N__39075\,
            I => \N__39066\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__39072\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__39069\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__39066\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__8427\ : InMux
    port map (
            O => \N__39059\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__8426\ : InMux
    port map (
            O => \N__39056\,
            I => \N__39051\
        );

    \I__8425\ : InMux
    port map (
            O => \N__39055\,
            I => \N__39046\
        );

    \I__8424\ : InMux
    port map (
            O => \N__39054\,
            I => \N__39046\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__39051\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__39046\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__8421\ : CascadeMux
    port map (
            O => \N__39041\,
            I => \N__39037\
        );

    \I__8420\ : InMux
    port map (
            O => \N__39040\,
            I => \N__39034\
        );

    \I__8419\ : InMux
    port map (
            O => \N__39037\,
            I => \N__39031\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__39034\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__39031\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__8416\ : InMux
    port map (
            O => \N__39026\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__8415\ : InMux
    port map (
            O => \N__39023\,
            I => \N__39018\
        );

    \I__8414\ : InMux
    port map (
            O => \N__39022\,
            I => \N__39013\
        );

    \I__8413\ : InMux
    port map (
            O => \N__39021\,
            I => \N__39013\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__39018\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__39013\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__8410\ : InMux
    port map (
            O => \N__39008\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__8409\ : CascadeMux
    port map (
            O => \N__39005\,
            I => \N__39002\
        );

    \I__8408\ : InMux
    port map (
            O => \N__39002\,
            I => \N__38997\
        );

    \I__8407\ : InMux
    port map (
            O => \N__39001\,
            I => \N__38994\
        );

    \I__8406\ : InMux
    port map (
            O => \N__39000\,
            I => \N__38991\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__38997\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__38994\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__38991\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__8402\ : InMux
    port map (
            O => \N__38984\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__8401\ : CascadeMux
    port map (
            O => \N__38981\,
            I => \N__38976\
        );

    \I__8400\ : CascadeMux
    port map (
            O => \N__38980\,
            I => \N__38973\
        );

    \I__8399\ : InMux
    port map (
            O => \N__38979\,
            I => \N__38970\
        );

    \I__8398\ : InMux
    port map (
            O => \N__38976\,
            I => \N__38965\
        );

    \I__8397\ : InMux
    port map (
            O => \N__38973\,
            I => \N__38965\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__38970\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__38965\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__8394\ : InMux
    port map (
            O => \N__38960\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__8393\ : CascadeMux
    port map (
            O => \N__38957\,
            I => \N__38954\
        );

    \I__8392\ : InMux
    port map (
            O => \N__38954\,
            I => \N__38949\
        );

    \I__8391\ : InMux
    port map (
            O => \N__38953\,
            I => \N__38946\
        );

    \I__8390\ : InMux
    port map (
            O => \N__38952\,
            I => \N__38943\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__38949\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__38946\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__38943\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__8386\ : InMux
    port map (
            O => \N__38936\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__8385\ : CascadeMux
    port map (
            O => \N__38933\,
            I => \N__38930\
        );

    \I__8384\ : InMux
    port map (
            O => \N__38930\,
            I => \N__38925\
        );

    \I__8383\ : InMux
    port map (
            O => \N__38929\,
            I => \N__38922\
        );

    \I__8382\ : InMux
    port map (
            O => \N__38928\,
            I => \N__38919\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__38925\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__38922\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__38919\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__8378\ : InMux
    port map (
            O => \N__38912\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__8377\ : CascadeMux
    port map (
            O => \N__38909\,
            I => \N__38906\
        );

    \I__8376\ : InMux
    port map (
            O => \N__38906\,
            I => \N__38901\
        );

    \I__8375\ : InMux
    port map (
            O => \N__38905\,
            I => \N__38898\
        );

    \I__8374\ : InMux
    port map (
            O => \N__38904\,
            I => \N__38895\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__38901\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__38898\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__38895\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__8370\ : InMux
    port map (
            O => \N__38888\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__8369\ : CascadeMux
    port map (
            O => \N__38885\,
            I => \N__38882\
        );

    \I__8368\ : InMux
    port map (
            O => \N__38882\,
            I => \N__38877\
        );

    \I__8367\ : InMux
    port map (
            O => \N__38881\,
            I => \N__38874\
        );

    \I__8366\ : InMux
    port map (
            O => \N__38880\,
            I => \N__38871\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__38877\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__38874\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__38871\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__8362\ : InMux
    port map (
            O => \N__38864\,
            I => \bfn_15_16_0_\
        );

    \I__8361\ : CascadeMux
    port map (
            O => \N__38861\,
            I => \N__38858\
        );

    \I__8360\ : InMux
    port map (
            O => \N__38858\,
            I => \N__38853\
        );

    \I__8359\ : InMux
    port map (
            O => \N__38857\,
            I => \N__38850\
        );

    \I__8358\ : InMux
    port map (
            O => \N__38856\,
            I => \N__38847\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__38853\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__38850\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__38847\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__8354\ : InMux
    port map (
            O => \N__38840\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__8353\ : CascadeMux
    port map (
            O => \N__38837\,
            I => \N__38834\
        );

    \I__8352\ : InMux
    port map (
            O => \N__38834\,
            I => \N__38829\
        );

    \I__8351\ : InMux
    port map (
            O => \N__38833\,
            I => \N__38826\
        );

    \I__8350\ : InMux
    port map (
            O => \N__38832\,
            I => \N__38823\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__38829\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__38826\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__38823\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__8346\ : InMux
    port map (
            O => \N__38816\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__8345\ : CascadeMux
    port map (
            O => \N__38813\,
            I => \N__38810\
        );

    \I__8344\ : InMux
    port map (
            O => \N__38810\,
            I => \N__38805\
        );

    \I__8343\ : InMux
    port map (
            O => \N__38809\,
            I => \N__38802\
        );

    \I__8342\ : InMux
    port map (
            O => \N__38808\,
            I => \N__38799\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__38805\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__38802\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__38799\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__8338\ : InMux
    port map (
            O => \N__38792\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__8337\ : CascadeMux
    port map (
            O => \N__38789\,
            I => \N__38786\
        );

    \I__8336\ : InMux
    port map (
            O => \N__38786\,
            I => \N__38781\
        );

    \I__8335\ : InMux
    port map (
            O => \N__38785\,
            I => \N__38778\
        );

    \I__8334\ : InMux
    port map (
            O => \N__38784\,
            I => \N__38775\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__38781\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__38778\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__38775\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__8330\ : InMux
    port map (
            O => \N__38768\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__8329\ : CascadeMux
    port map (
            O => \N__38765\,
            I => \N__38762\
        );

    \I__8328\ : InMux
    port map (
            O => \N__38762\,
            I => \N__38757\
        );

    \I__8327\ : InMux
    port map (
            O => \N__38761\,
            I => \N__38754\
        );

    \I__8326\ : InMux
    port map (
            O => \N__38760\,
            I => \N__38751\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__38757\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__38754\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__38751\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__8322\ : InMux
    port map (
            O => \N__38744\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__8321\ : CascadeMux
    port map (
            O => \N__38741\,
            I => \N__38738\
        );

    \I__8320\ : InMux
    port map (
            O => \N__38738\,
            I => \N__38733\
        );

    \I__8319\ : InMux
    port map (
            O => \N__38737\,
            I => \N__38730\
        );

    \I__8318\ : InMux
    port map (
            O => \N__38736\,
            I => \N__38727\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__38733\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__38730\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__38727\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__8314\ : InMux
    port map (
            O => \N__38720\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__8313\ : CascadeMux
    port map (
            O => \N__38717\,
            I => \N__38714\
        );

    \I__8312\ : InMux
    port map (
            O => \N__38714\,
            I => \N__38709\
        );

    \I__8311\ : InMux
    port map (
            O => \N__38713\,
            I => \N__38706\
        );

    \I__8310\ : InMux
    port map (
            O => \N__38712\,
            I => \N__38703\
        );

    \I__8309\ : LocalMux
    port map (
            O => \N__38709\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__38706\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__38703\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__8306\ : InMux
    port map (
            O => \N__38696\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__8305\ : CascadeMux
    port map (
            O => \N__38693\,
            I => \N__38690\
        );

    \I__8304\ : InMux
    port map (
            O => \N__38690\,
            I => \N__38685\
        );

    \I__8303\ : InMux
    port map (
            O => \N__38689\,
            I => \N__38682\
        );

    \I__8302\ : InMux
    port map (
            O => \N__38688\,
            I => \N__38679\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__38685\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__38682\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__38679\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__8298\ : InMux
    port map (
            O => \N__38672\,
            I => \bfn_15_15_0_\
        );

    \I__8297\ : CascadeMux
    port map (
            O => \N__38669\,
            I => \N__38666\
        );

    \I__8296\ : InMux
    port map (
            O => \N__38666\,
            I => \N__38661\
        );

    \I__8295\ : InMux
    port map (
            O => \N__38665\,
            I => \N__38658\
        );

    \I__8294\ : InMux
    port map (
            O => \N__38664\,
            I => \N__38655\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__38661\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__38658\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__38655\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__8290\ : InMux
    port map (
            O => \N__38648\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__8289\ : CascadeMux
    port map (
            O => \N__38645\,
            I => \N__38642\
        );

    \I__8288\ : InMux
    port map (
            O => \N__38642\,
            I => \N__38636\
        );

    \I__8287\ : InMux
    port map (
            O => \N__38641\,
            I => \N__38636\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__38636\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\
        );

    \I__8285\ : CascadeMux
    port map (
            O => \N__38633\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12_cascade_\
        );

    \I__8284\ : InMux
    port map (
            O => \N__38630\,
            I => \N__38627\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__38627\,
            I => \N__38624\
        );

    \I__8282\ : Span4Mux_v
    port map (
            O => \N__38624\,
            I => \N__38621\
        );

    \I__8281\ : Odrv4
    port map (
            O => \N__38621\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__8280\ : InMux
    port map (
            O => \N__38618\,
            I => \N__38615\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__38615\,
            I => \N__38612\
        );

    \I__8278\ : Span4Mux_v
    port map (
            O => \N__38612\,
            I => \N__38609\
        );

    \I__8277\ : Odrv4
    port map (
            O => \N__38609\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__8276\ : InMux
    port map (
            O => \N__38606\,
            I => \N__38600\
        );

    \I__8275\ : InMux
    port map (
            O => \N__38605\,
            I => \N__38600\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__38600\,
            I => \N__38597\
        );

    \I__8273\ : Span4Mux_h
    port map (
            O => \N__38597\,
            I => \N__38594\
        );

    \I__8272\ : Odrv4
    port map (
            O => \N__38594\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\
        );

    \I__8271\ : InMux
    port map (
            O => \N__38591\,
            I => \N__38588\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__38588\,
            I => \N__38585\
        );

    \I__8269\ : Span4Mux_h
    port map (
            O => \N__38585\,
            I => \N__38581\
        );

    \I__8268\ : InMux
    port map (
            O => \N__38584\,
            I => \N__38578\
        );

    \I__8267\ : Odrv4
    port map (
            O => \N__38581\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__38578\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__8265\ : InMux
    port map (
            O => \N__38573\,
            I => \N__38570\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__38570\,
            I => \N__38566\
        );

    \I__8263\ : CascadeMux
    port map (
            O => \N__38569\,
            I => \N__38563\
        );

    \I__8262\ : Span4Mux_h
    port map (
            O => \N__38566\,
            I => \N__38559\
        );

    \I__8261\ : InMux
    port map (
            O => \N__38563\,
            I => \N__38556\
        );

    \I__8260\ : InMux
    port map (
            O => \N__38562\,
            I => \N__38553\
        );

    \I__8259\ : Odrv4
    port map (
            O => \N__38559\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__38556\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__38553\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__8256\ : InMux
    port map (
            O => \N__38546\,
            I => \N__38543\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__38543\,
            I => \N__38539\
        );

    \I__8254\ : CascadeMux
    port map (
            O => \N__38542\,
            I => \N__38536\
        );

    \I__8253\ : Span4Mux_v
    port map (
            O => \N__38539\,
            I => \N__38532\
        );

    \I__8252\ : InMux
    port map (
            O => \N__38536\,
            I => \N__38529\
        );

    \I__8251\ : InMux
    port map (
            O => \N__38535\,
            I => \N__38526\
        );

    \I__8250\ : Odrv4
    port map (
            O => \N__38532\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__38529\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__38526\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__8247\ : InMux
    port map (
            O => \N__38519\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__8246\ : InMux
    port map (
            O => \N__38516\,
            I => \N__38513\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__38513\,
            I => \N__38510\
        );

    \I__8244\ : Span4Mux_h
    port map (
            O => \N__38510\,
            I => \N__38507\
        );

    \I__8243\ : Odrv4
    port map (
            O => \N__38507\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt20\
        );

    \I__8242\ : CascadeMux
    port map (
            O => \N__38504\,
            I => \N__38499\
        );

    \I__8241\ : InMux
    port map (
            O => \N__38503\,
            I => \N__38496\
        );

    \I__8240\ : InMux
    port map (
            O => \N__38502\,
            I => \N__38491\
        );

    \I__8239\ : InMux
    port map (
            O => \N__38499\,
            I => \N__38491\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__38496\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__38491\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__8236\ : CascadeMux
    port map (
            O => \N__38486\,
            I => \N__38481\
        );

    \I__8235\ : InMux
    port map (
            O => \N__38485\,
            I => \N__38478\
        );

    \I__8234\ : InMux
    port map (
            O => \N__38484\,
            I => \N__38473\
        );

    \I__8233\ : InMux
    port map (
            O => \N__38481\,
            I => \N__38473\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__38478\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__38473\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__8230\ : CascadeMux
    port map (
            O => \N__38468\,
            I => \N__38465\
        );

    \I__8229\ : InMux
    port map (
            O => \N__38465\,
            I => \N__38462\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__38462\,
            I => \N__38459\
        );

    \I__8227\ : Span4Mux_h
    port map (
            O => \N__38459\,
            I => \N__38456\
        );

    \I__8226\ : Odrv4
    port map (
            O => \N__38456\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\
        );

    \I__8225\ : InMux
    port map (
            O => \N__38453\,
            I => \N__38447\
        );

    \I__8224\ : InMux
    port map (
            O => \N__38452\,
            I => \N__38447\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__38447\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\
        );

    \I__8222\ : InMux
    port map (
            O => \N__38444\,
            I => \N__38438\
        );

    \I__8221\ : InMux
    port map (
            O => \N__38443\,
            I => \N__38438\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__38438\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\
        );

    \I__8219\ : InMux
    port map (
            O => \N__38435\,
            I => \N__38432\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__38432\,
            I => \N__38429\
        );

    \I__8217\ : Span4Mux_h
    port map (
            O => \N__38429\,
            I => \N__38426\
        );

    \I__8216\ : Odrv4
    port map (
            O => \N__38426\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__8215\ : CascadeMux
    port map (
            O => \N__38423\,
            I => \N__38420\
        );

    \I__8214\ : InMux
    port map (
            O => \N__38420\,
            I => \N__38417\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__38417\,
            I => \N__38414\
        );

    \I__8212\ : Span4Mux_h
    port map (
            O => \N__38414\,
            I => \N__38411\
        );

    \I__8211\ : Odrv4
    port map (
            O => \N__38411\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt22\
        );

    \I__8210\ : InMux
    port map (
            O => \N__38408\,
            I => \N__38403\
        );

    \I__8209\ : InMux
    port map (
            O => \N__38407\,
            I => \N__38400\
        );

    \I__8208\ : InMux
    port map (
            O => \N__38406\,
            I => \N__38397\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__38403\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__38400\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__38397\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__8204\ : CascadeMux
    port map (
            O => \N__38390\,
            I => \N__38386\
        );

    \I__8203\ : InMux
    port map (
            O => \N__38389\,
            I => \N__38382\
        );

    \I__8202\ : InMux
    port map (
            O => \N__38386\,
            I => \N__38379\
        );

    \I__8201\ : InMux
    port map (
            O => \N__38385\,
            I => \N__38376\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__38382\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__38379\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__38376\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__8197\ : InMux
    port map (
            O => \N__38369\,
            I => \N__38366\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__38366\,
            I => \N__38363\
        );

    \I__8195\ : Odrv4
    port map (
            O => \N__38363\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\
        );

    \I__8194\ : InMux
    port map (
            O => \N__38360\,
            I => \N__38354\
        );

    \I__8193\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38354\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__38354\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\
        );

    \I__8191\ : InMux
    port map (
            O => \N__38351\,
            I => \N__38348\
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__38348\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__8189\ : InMux
    port map (
            O => \N__38345\,
            I => \N__38342\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__38342\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__8187\ : CascadeMux
    port map (
            O => \N__38339\,
            I => \N__38336\
        );

    \I__8186\ : InMux
    port map (
            O => \N__38336\,
            I => \N__38333\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__38333\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__8184\ : CascadeMux
    port map (
            O => \N__38330\,
            I => \N__38327\
        );

    \I__8183\ : InMux
    port map (
            O => \N__38327\,
            I => \N__38324\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__38324\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt24\
        );

    \I__8181\ : InMux
    port map (
            O => \N__38321\,
            I => \N__38315\
        );

    \I__8180\ : InMux
    port map (
            O => \N__38320\,
            I => \N__38315\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__38315\,
            I => \N__38311\
        );

    \I__8178\ : InMux
    port map (
            O => \N__38314\,
            I => \N__38308\
        );

    \I__8177\ : Span4Mux_h
    port map (
            O => \N__38311\,
            I => \N__38305\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__38308\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__8175\ : Odrv4
    port map (
            O => \N__38305\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__8174\ : CascadeMux
    port map (
            O => \N__38300\,
            I => \N__38297\
        );

    \I__8173\ : InMux
    port map (
            O => \N__38297\,
            I => \N__38291\
        );

    \I__8172\ : InMux
    port map (
            O => \N__38296\,
            I => \N__38291\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__38291\,
            I => \N__38287\
        );

    \I__8170\ : InMux
    port map (
            O => \N__38290\,
            I => \N__38284\
        );

    \I__8169\ : Span4Mux_h
    port map (
            O => \N__38287\,
            I => \N__38281\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__38284\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__8167\ : Odrv4
    port map (
            O => \N__38281\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__8166\ : InMux
    port map (
            O => \N__38276\,
            I => \N__38273\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__38273\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\
        );

    \I__8164\ : InMux
    port map (
            O => \N__38270\,
            I => \pwm_generator_inst.un3_threshold_cry_19\
        );

    \I__8163\ : InMux
    port map (
            O => \N__38267\,
            I => \N__38264\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__38264\,
            I => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\
        );

    \I__8161\ : InMux
    port map (
            O => \N__38261\,
            I => \N__38257\
        );

    \I__8160\ : InMux
    port map (
            O => \N__38260\,
            I => \N__38253\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__38257\,
            I => \N__38250\
        );

    \I__8158\ : InMux
    port map (
            O => \N__38256\,
            I => \N__38246\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__38253\,
            I => \N__38243\
        );

    \I__8156\ : Span4Mux_v
    port map (
            O => \N__38250\,
            I => \N__38240\
        );

    \I__8155\ : InMux
    port map (
            O => \N__38249\,
            I => \N__38237\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__38246\,
            I => \N__38234\
        );

    \I__8153\ : Span4Mux_v
    port map (
            O => \N__38243\,
            I => \N__38231\
        );

    \I__8152\ : Span4Mux_h
    port map (
            O => \N__38240\,
            I => \N__38228\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__38237\,
            I => \N__38225\
        );

    \I__8150\ : Span4Mux_h
    port map (
            O => \N__38234\,
            I => \N__38222\
        );

    \I__8149\ : Span4Mux_v
    port map (
            O => \N__38231\,
            I => \N__38219\
        );

    \I__8148\ : Span4Mux_h
    port map (
            O => \N__38228\,
            I => \N__38216\
        );

    \I__8147\ : Span4Mux_v
    port map (
            O => \N__38225\,
            I => \N__38213\
        );

    \I__8146\ : Odrv4
    port map (
            O => \N__38222\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__8145\ : Odrv4
    port map (
            O => \N__38219\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__8144\ : Odrv4
    port map (
            O => \N__38216\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__8143\ : Odrv4
    port map (
            O => \N__38213\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__8142\ : InMux
    port map (
            O => \N__38204\,
            I => \N__38201\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__38201\,
            I => \N__38197\
        );

    \I__8140\ : InMux
    port map (
            O => \N__38200\,
            I => \N__38193\
        );

    \I__8139\ : Span4Mux_h
    port map (
            O => \N__38197\,
            I => \N__38190\
        );

    \I__8138\ : InMux
    port map (
            O => \N__38196\,
            I => \N__38187\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__38193\,
            I => \N__38184\
        );

    \I__8136\ : Span4Mux_v
    port map (
            O => \N__38190\,
            I => \N__38181\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__38187\,
            I => \N__38176\
        );

    \I__8134\ : Span4Mux_h
    port map (
            O => \N__38184\,
            I => \N__38176\
        );

    \I__8133\ : Odrv4
    port map (
            O => \N__38181\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__8132\ : Odrv4
    port map (
            O => \N__38176\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__8131\ : CascadeMux
    port map (
            O => \N__38171\,
            I => \N__38168\
        );

    \I__8130\ : InMux
    port map (
            O => \N__38168\,
            I => \N__38165\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__38165\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38162\,
            I => \N__38159\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__38159\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__8126\ : InMux
    port map (
            O => \N__38156\,
            I => \N__38153\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__38153\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__8124\ : InMux
    port map (
            O => \N__38150\,
            I => \N__38147\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__38147\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__8122\ : CascadeMux
    port map (
            O => \N__38144\,
            I => \N__38141\
        );

    \I__8121\ : InMux
    port map (
            O => \N__38141\,
            I => \N__38138\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__38138\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt18\
        );

    \I__8119\ : InMux
    port map (
            O => \N__38135\,
            I => \N__38129\
        );

    \I__8118\ : InMux
    port map (
            O => \N__38134\,
            I => \N__38129\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__38129\,
            I => \N__38125\
        );

    \I__8116\ : InMux
    port map (
            O => \N__38128\,
            I => \N__38122\
        );

    \I__8115\ : Span4Mux_h
    port map (
            O => \N__38125\,
            I => \N__38119\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__38122\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8113\ : Odrv4
    port map (
            O => \N__38119\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8112\ : CascadeMux
    port map (
            O => \N__38114\,
            I => \N__38110\
        );

    \I__8111\ : InMux
    port map (
            O => \N__38113\,
            I => \N__38105\
        );

    \I__8110\ : InMux
    port map (
            O => \N__38110\,
            I => \N__38105\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__38105\,
            I => \N__38102\
        );

    \I__8108\ : Span4Mux_h
    port map (
            O => \N__38102\,
            I => \N__38099\
        );

    \I__8107\ : Span4Mux_v
    port map (
            O => \N__38099\,
            I => \N__38096\
        );

    \I__8106\ : Odrv4
    port map (
            O => \N__38096\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__8105\ : CascadeMux
    port map (
            O => \N__38093\,
            I => \N__38089\
        );

    \I__8104\ : InMux
    port map (
            O => \N__38092\,
            I => \N__38084\
        );

    \I__8103\ : InMux
    port map (
            O => \N__38089\,
            I => \N__38084\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__38084\,
            I => \N__38080\
        );

    \I__8101\ : InMux
    port map (
            O => \N__38083\,
            I => \N__38077\
        );

    \I__8100\ : Span4Mux_h
    port map (
            O => \N__38080\,
            I => \N__38074\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__38077\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8098\ : Odrv4
    port map (
            O => \N__38074\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8097\ : InMux
    port map (
            O => \N__38069\,
            I => \N__38066\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__38066\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\
        );

    \I__8095\ : InMux
    port map (
            O => \N__38063\,
            I => \N__38060\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__38060\,
            I => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\
        );

    \I__8093\ : InMux
    port map (
            O => \N__38057\,
            I => \N__38054\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__38054\,
            I => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\
        );

    \I__8091\ : InMux
    port map (
            O => \N__38051\,
            I => \N__38048\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__38048\,
            I => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\
        );

    \I__8089\ : InMux
    port map (
            O => \N__38045\,
            I => \N__38042\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__38042\,
            I => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\
        );

    \I__8087\ : InMux
    port map (
            O => \N__38039\,
            I => \N__38036\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__38036\,
            I => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\
        );

    \I__8085\ : InMux
    port map (
            O => \N__38033\,
            I => \N__38030\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__38030\,
            I => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\
        );

    \I__8083\ : InMux
    port map (
            O => \N__38027\,
            I => \N__38024\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__38024\,
            I => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\
        );

    \I__8081\ : InMux
    port map (
            O => \N__38021\,
            I => \N__38018\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__38018\,
            I => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\
        );

    \I__8079\ : InMux
    port map (
            O => \N__38015\,
            I => \N__38012\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__38012\,
            I => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\
        );

    \I__8077\ : InMux
    port map (
            O => \N__38009\,
            I => \N__38006\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__38006\,
            I => \N__38003\
        );

    \I__8075\ : Sp12to4
    port map (
            O => \N__38003\,
            I => \N__38000\
        );

    \I__8074\ : Span12Mux_s6_v
    port map (
            O => \N__38000\,
            I => \N__37997\
        );

    \I__8073\ : Odrv12
    port map (
            O => \N__37997\,
            I => \pwm_generator_inst.O_14\
        );

    \I__8072\ : InMux
    port map (
            O => \N__37994\,
            I => \pwm_generator_inst.un3_threshold_cry_2\
        );

    \I__8071\ : InMux
    port map (
            O => \N__37991\,
            I => \N__37988\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__37988\,
            I => \pwm_generator_inst.un3_threshold_axbZ0Z_4\
        );

    \I__8069\ : CascadeMux
    port map (
            O => \N__37985\,
            I => \N__37982\
        );

    \I__8068\ : InMux
    port map (
            O => \N__37982\,
            I => \N__37979\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__37979\,
            I => \N__37975\
        );

    \I__8066\ : InMux
    port map (
            O => \N__37978\,
            I => \N__37972\
        );

    \I__8065\ : Odrv4
    port map (
            O => \N__37975\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__37972\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__8063\ : InMux
    port map (
            O => \N__37967\,
            I => \pwm_generator_inst.un3_threshold_cry_3\
        );

    \I__8062\ : CascadeMux
    port map (
            O => \N__37964\,
            I => \N__37961\
        );

    \I__8061\ : InMux
    port map (
            O => \N__37961\,
            I => \N__37958\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__37958\,
            I => \N__37955\
        );

    \I__8059\ : Odrv4
    port map (
            O => \N__37955\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\
        );

    \I__8058\ : InMux
    port map (
            O => \N__37952\,
            I => \N__37949\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__37949\,
            I => \N__37945\
        );

    \I__8056\ : InMux
    port map (
            O => \N__37948\,
            I => \N__37942\
        );

    \I__8055\ : Odrv4
    port map (
            O => \N__37945\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__37942\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__8053\ : InMux
    port map (
            O => \N__37937\,
            I => \pwm_generator_inst.un3_threshold_cry_4\
        );

    \I__8052\ : InMux
    port map (
            O => \N__37934\,
            I => \N__37931\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__37931\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\
        );

    \I__8050\ : InMux
    port map (
            O => \N__37928\,
            I => \N__37924\
        );

    \I__8049\ : InMux
    port map (
            O => \N__37927\,
            I => \N__37921\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__37924\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__37921\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__8046\ : InMux
    port map (
            O => \N__37916\,
            I => \pwm_generator_inst.un3_threshold_cry_5\
        );

    \I__8045\ : InMux
    port map (
            O => \N__37913\,
            I => \N__37910\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__37910\,
            I => \N__37895\
        );

    \I__8043\ : InMux
    port map (
            O => \N__37909\,
            I => \N__37892\
        );

    \I__8042\ : CascadeMux
    port map (
            O => \N__37908\,
            I => \N__37875\
        );

    \I__8041\ : CascadeMux
    port map (
            O => \N__37907\,
            I => \N__37871\
        );

    \I__8040\ : CascadeMux
    port map (
            O => \N__37906\,
            I => \N__37867\
        );

    \I__8039\ : CascadeMux
    port map (
            O => \N__37905\,
            I => \N__37862\
        );

    \I__8038\ : CascadeMux
    port map (
            O => \N__37904\,
            I => \N__37858\
        );

    \I__8037\ : CascadeMux
    port map (
            O => \N__37903\,
            I => \N__37854\
        );

    \I__8036\ : CascadeMux
    port map (
            O => \N__37902\,
            I => \N__37850\
        );

    \I__8035\ : CascadeMux
    port map (
            O => \N__37901\,
            I => \N__37847\
        );

    \I__8034\ : CascadeMux
    port map (
            O => \N__37900\,
            I => \N__37843\
        );

    \I__8033\ : CascadeMux
    port map (
            O => \N__37899\,
            I => \N__37839\
        );

    \I__8032\ : CascadeMux
    port map (
            O => \N__37898\,
            I => \N__37835\
        );

    \I__8031\ : Span4Mux_s2_v
    port map (
            O => \N__37895\,
            I => \N__37826\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__37892\,
            I => \N__37826\
        );

    \I__8029\ : InMux
    port map (
            O => \N__37891\,
            I => \N__37819\
        );

    \I__8028\ : InMux
    port map (
            O => \N__37890\,
            I => \N__37819\
        );

    \I__8027\ : InMux
    port map (
            O => \N__37889\,
            I => \N__37819\
        );

    \I__8026\ : InMux
    port map (
            O => \N__37888\,
            I => \N__37810\
        );

    \I__8025\ : InMux
    port map (
            O => \N__37887\,
            I => \N__37810\
        );

    \I__8024\ : InMux
    port map (
            O => \N__37886\,
            I => \N__37810\
        );

    \I__8023\ : InMux
    port map (
            O => \N__37885\,
            I => \N__37810\
        );

    \I__8022\ : InMux
    port map (
            O => \N__37884\,
            I => \N__37807\
        );

    \I__8021\ : InMux
    port map (
            O => \N__37883\,
            I => \N__37802\
        );

    \I__8020\ : InMux
    port map (
            O => \N__37882\,
            I => \N__37802\
        );

    \I__8019\ : InMux
    port map (
            O => \N__37881\,
            I => \N__37799\
        );

    \I__8018\ : InMux
    port map (
            O => \N__37880\,
            I => \N__37779\
        );

    \I__8017\ : InMux
    port map (
            O => \N__37879\,
            I => \N__37779\
        );

    \I__8016\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37764\
        );

    \I__8015\ : InMux
    port map (
            O => \N__37875\,
            I => \N__37764\
        );

    \I__8014\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37764\
        );

    \I__8013\ : InMux
    port map (
            O => \N__37871\,
            I => \N__37764\
        );

    \I__8012\ : InMux
    port map (
            O => \N__37870\,
            I => \N__37764\
        );

    \I__8011\ : InMux
    port map (
            O => \N__37867\,
            I => \N__37764\
        );

    \I__8010\ : InMux
    port map (
            O => \N__37866\,
            I => \N__37764\
        );

    \I__8009\ : InMux
    port map (
            O => \N__37865\,
            I => \N__37747\
        );

    \I__8008\ : InMux
    port map (
            O => \N__37862\,
            I => \N__37747\
        );

    \I__8007\ : InMux
    port map (
            O => \N__37861\,
            I => \N__37747\
        );

    \I__8006\ : InMux
    port map (
            O => \N__37858\,
            I => \N__37747\
        );

    \I__8005\ : InMux
    port map (
            O => \N__37857\,
            I => \N__37747\
        );

    \I__8004\ : InMux
    port map (
            O => \N__37854\,
            I => \N__37747\
        );

    \I__8003\ : InMux
    port map (
            O => \N__37853\,
            I => \N__37747\
        );

    \I__8002\ : InMux
    port map (
            O => \N__37850\,
            I => \N__37747\
        );

    \I__8001\ : InMux
    port map (
            O => \N__37847\,
            I => \N__37730\
        );

    \I__8000\ : InMux
    port map (
            O => \N__37846\,
            I => \N__37730\
        );

    \I__7999\ : InMux
    port map (
            O => \N__37843\,
            I => \N__37730\
        );

    \I__7998\ : InMux
    port map (
            O => \N__37842\,
            I => \N__37730\
        );

    \I__7997\ : InMux
    port map (
            O => \N__37839\,
            I => \N__37730\
        );

    \I__7996\ : InMux
    port map (
            O => \N__37838\,
            I => \N__37730\
        );

    \I__7995\ : InMux
    port map (
            O => \N__37835\,
            I => \N__37730\
        );

    \I__7994\ : InMux
    port map (
            O => \N__37834\,
            I => \N__37730\
        );

    \I__7993\ : CascadeMux
    port map (
            O => \N__37833\,
            I => \N__37726\
        );

    \I__7992\ : CascadeMux
    port map (
            O => \N__37832\,
            I => \N__37722\
        );

    \I__7991\ : CascadeMux
    port map (
            O => \N__37831\,
            I => \N__37718\
        );

    \I__7990\ : Span4Mux_v
    port map (
            O => \N__37826\,
            I => \N__37709\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__37819\,
            I => \N__37709\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__37810\,
            I => \N__37709\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__37807\,
            I => \N__37702\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__37802\,
            I => \N__37702\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__37799\,
            I => \N__37702\
        );

    \I__7984\ : InMux
    port map (
            O => \N__37798\,
            I => \N__37699\
        );

    \I__7983\ : InMux
    port map (
            O => \N__37797\,
            I => \N__37694\
        );

    \I__7982\ : InMux
    port map (
            O => \N__37796\,
            I => \N__37694\
        );

    \I__7981\ : InMux
    port map (
            O => \N__37795\,
            I => \N__37691\
        );

    \I__7980\ : InMux
    port map (
            O => \N__37794\,
            I => \N__37688\
        );

    \I__7979\ : InMux
    port map (
            O => \N__37793\,
            I => \N__37685\
        );

    \I__7978\ : InMux
    port map (
            O => \N__37792\,
            I => \N__37682\
        );

    \I__7977\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37679\
        );

    \I__7976\ : InMux
    port map (
            O => \N__37790\,
            I => \N__37672\
        );

    \I__7975\ : InMux
    port map (
            O => \N__37789\,
            I => \N__37672\
        );

    \I__7974\ : InMux
    port map (
            O => \N__37788\,
            I => \N__37672\
        );

    \I__7973\ : InMux
    port map (
            O => \N__37787\,
            I => \N__37663\
        );

    \I__7972\ : InMux
    port map (
            O => \N__37786\,
            I => \N__37663\
        );

    \I__7971\ : InMux
    port map (
            O => \N__37785\,
            I => \N__37663\
        );

    \I__7970\ : InMux
    port map (
            O => \N__37784\,
            I => \N__37663\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__37779\,
            I => \N__37660\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__37764\,
            I => \N__37655\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__37747\,
            I => \N__37655\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__37730\,
            I => \N__37652\
        );

    \I__7965\ : InMux
    port map (
            O => \N__37729\,
            I => \N__37637\
        );

    \I__7964\ : InMux
    port map (
            O => \N__37726\,
            I => \N__37637\
        );

    \I__7963\ : InMux
    port map (
            O => \N__37725\,
            I => \N__37637\
        );

    \I__7962\ : InMux
    port map (
            O => \N__37722\,
            I => \N__37637\
        );

    \I__7961\ : InMux
    port map (
            O => \N__37721\,
            I => \N__37637\
        );

    \I__7960\ : InMux
    port map (
            O => \N__37718\,
            I => \N__37637\
        );

    \I__7959\ : InMux
    port map (
            O => \N__37717\,
            I => \N__37637\
        );

    \I__7958\ : CascadeMux
    port map (
            O => \N__37716\,
            I => \N__37633\
        );

    \I__7957\ : Span4Mux_v
    port map (
            O => \N__37709\,
            I => \N__37629\
        );

    \I__7956\ : Span12Mux_s7_v
    port map (
            O => \N__37702\,
            I => \N__37620\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__37699\,
            I => \N__37620\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__37694\,
            I => \N__37620\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__37691\,
            I => \N__37620\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__37688\,
            I => \N__37607\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__37685\,
            I => \N__37607\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__37682\,
            I => \N__37607\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__37679\,
            I => \N__37607\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__37672\,
            I => \N__37607\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__37663\,
            I => \N__37607\
        );

    \I__7946\ : Span4Mux_h
    port map (
            O => \N__37660\,
            I => \N__37604\
        );

    \I__7945\ : Span4Mux_v
    port map (
            O => \N__37655\,
            I => \N__37601\
        );

    \I__7944\ : Span4Mux_h
    port map (
            O => \N__37652\,
            I => \N__37596\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__37637\,
            I => \N__37596\
        );

    \I__7942\ : InMux
    port map (
            O => \N__37636\,
            I => \N__37589\
        );

    \I__7941\ : InMux
    port map (
            O => \N__37633\,
            I => \N__37589\
        );

    \I__7940\ : InMux
    port map (
            O => \N__37632\,
            I => \N__37589\
        );

    \I__7939\ : Sp12to4
    port map (
            O => \N__37629\,
            I => \N__37586\
        );

    \I__7938\ : Span12Mux_v
    port map (
            O => \N__37620\,
            I => \N__37581\
        );

    \I__7937\ : Span12Mux_s10_v
    port map (
            O => \N__37607\,
            I => \N__37581\
        );

    \I__7936\ : Span4Mux_v
    port map (
            O => \N__37604\,
            I => \N__37578\
        );

    \I__7935\ : Span4Mux_v
    port map (
            O => \N__37601\,
            I => \N__37573\
        );

    \I__7934\ : Span4Mux_v
    port map (
            O => \N__37596\,
            I => \N__37573\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__37589\,
            I => \N__37570\
        );

    \I__7932\ : Span12Mux_h
    port map (
            O => \N__37586\,
            I => \N__37565\
        );

    \I__7931\ : Span12Mux_h
    port map (
            O => \N__37581\,
            I => \N__37565\
        );

    \I__7930\ : Span4Mux_v
    port map (
            O => \N__37578\,
            I => \N__37562\
        );

    \I__7929\ : Span4Mux_v
    port map (
            O => \N__37573\,
            I => \N__37559\
        );

    \I__7928\ : Span4Mux_v
    port map (
            O => \N__37570\,
            I => \N__37556\
        );

    \I__7927\ : Odrv12
    port map (
            O => \N__37565\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7926\ : Odrv4
    port map (
            O => \N__37562\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7925\ : Odrv4
    port map (
            O => \N__37559\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7924\ : Odrv4
    port map (
            O => \N__37556\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7923\ : CascadeMux
    port map (
            O => \N__37547\,
            I => \N__37544\
        );

    \I__7922\ : InMux
    port map (
            O => \N__37544\,
            I => \N__37541\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__37541\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\
        );

    \I__7920\ : InMux
    port map (
            O => \N__37538\,
            I => \N__37535\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__37535\,
            I => \N__37531\
        );

    \I__7918\ : InMux
    port map (
            O => \N__37534\,
            I => \N__37528\
        );

    \I__7917\ : Odrv4
    port map (
            O => \N__37531\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__37528\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__7915\ : InMux
    port map (
            O => \N__37523\,
            I => \pwm_generator_inst.un3_threshold_cry_6\
        );

    \I__7914\ : InMux
    port map (
            O => \N__37520\,
            I => \N__37517\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__37517\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\
        );

    \I__7912\ : InMux
    port map (
            O => \N__37514\,
            I => \N__37511\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__37511\,
            I => \N__37508\
        );

    \I__7910\ : Span4Mux_v
    port map (
            O => \N__37508\,
            I => \N__37505\
        );

    \I__7909\ : Odrv4
    port map (
            O => \N__37505\,
            I => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\
        );

    \I__7908\ : InMux
    port map (
            O => \N__37502\,
            I => \bfn_14_29_0_\
        );

    \I__7907\ : InMux
    port map (
            O => \N__37499\,
            I => \N__37496\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__37496\,
            I => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\
        );

    \I__7905\ : InMux
    port map (
            O => \N__37493\,
            I => \N__37490\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__37490\,
            I => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\
        );

    \I__7903\ : InMux
    port map (
            O => \N__37487\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17\
        );

    \I__7902\ : InMux
    port map (
            O => \N__37484\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18\
        );

    \I__7901\ : InMux
    port map (
            O => \N__37481\,
            I => \N__37478\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__37478\,
            I => \N__37475\
        );

    \I__7899\ : Odrv4
    port map (
            O => \N__37475\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\
        );

    \I__7898\ : CascadeMux
    port map (
            O => \N__37472\,
            I => \N__37469\
        );

    \I__7897\ : InMux
    port map (
            O => \N__37469\,
            I => \N__37464\
        );

    \I__7896\ : InMux
    port map (
            O => \N__37468\,
            I => \N__37459\
        );

    \I__7895\ : InMux
    port map (
            O => \N__37467\,
            I => \N__37459\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__37464\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__37459\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__7892\ : InMux
    port map (
            O => \N__37454\,
            I => \N__37449\
        );

    \I__7891\ : InMux
    port map (
            O => \N__37453\,
            I => \N__37444\
        );

    \I__7890\ : InMux
    port map (
            O => \N__37452\,
            I => \N__37444\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__37449\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__37444\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__7887\ : InMux
    port map (
            O => \N__37439\,
            I => \N__37435\
        );

    \I__7886\ : InMux
    port map (
            O => \N__37438\,
            I => \N__37431\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__37435\,
            I => \N__37428\
        );

    \I__7884\ : InMux
    port map (
            O => \N__37434\,
            I => \N__37425\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__37431\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__7882\ : Odrv4
    port map (
            O => \N__37428\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__37425\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__7880\ : CascadeMux
    port map (
            O => \N__37418\,
            I => \N__37414\
        );

    \I__7879\ : InMux
    port map (
            O => \N__37417\,
            I => \N__37410\
        );

    \I__7878\ : InMux
    port map (
            O => \N__37414\,
            I => \N__37407\
        );

    \I__7877\ : InMux
    port map (
            O => \N__37413\,
            I => \N__37404\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__37410\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__37407\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__37404\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__7873\ : InMux
    port map (
            O => \N__37397\,
            I => \N__37394\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__37394\,
            I => \N__37390\
        );

    \I__7871\ : InMux
    port map (
            O => \N__37393\,
            I => \N__37387\
        );

    \I__7870\ : Span4Mux_v
    port map (
            O => \N__37390\,
            I => \N__37382\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__37387\,
            I => \N__37382\
        );

    \I__7868\ : Span4Mux_h
    port map (
            O => \N__37382\,
            I => \N__37379\
        );

    \I__7867\ : Span4Mux_h
    port map (
            O => \N__37379\,
            I => \N__37376\
        );

    \I__7866\ : Span4Mux_v
    port map (
            O => \N__37376\,
            I => \N__37373\
        );

    \I__7865\ : Odrv4
    port map (
            O => \N__37373\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__7864\ : InMux
    port map (
            O => \N__37370\,
            I => \N__37367\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__37367\,
            I => \N__37364\
        );

    \I__7862\ : Span12Mux_h
    port map (
            O => \N__37364\,
            I => \N__37361\
        );

    \I__7861\ : Odrv12
    port map (
            O => \N__37361\,
            I => \pwm_generator_inst.O_12\
        );

    \I__7860\ : InMux
    port map (
            O => \N__37358\,
            I => \N__37355\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__37355\,
            I => \N__37351\
        );

    \I__7858\ : InMux
    port map (
            O => \N__37354\,
            I => \N__37348\
        );

    \I__7857\ : Odrv4
    port map (
            O => \N__37351\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__37348\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__7855\ : InMux
    port map (
            O => \N__37343\,
            I => \pwm_generator_inst.un3_threshold_cry_0\
        );

    \I__7854\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37337\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__37337\,
            I => \N__37334\
        );

    \I__7852\ : Span4Mux_v
    port map (
            O => \N__37334\,
            I => \N__37331\
        );

    \I__7851\ : Span4Mux_h
    port map (
            O => \N__37331\,
            I => \N__37328\
        );

    \I__7850\ : Span4Mux_h
    port map (
            O => \N__37328\,
            I => \N__37325\
        );

    \I__7849\ : Odrv4
    port map (
            O => \N__37325\,
            I => \pwm_generator_inst.O_13\
        );

    \I__7848\ : InMux
    port map (
            O => \N__37322\,
            I => \pwm_generator_inst.un3_threshold_cry_1\
        );

    \I__7847\ : InMux
    port map (
            O => \N__37319\,
            I => \N__37316\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__37316\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\
        );

    \I__7845\ : InMux
    port map (
            O => \N__37313\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9\
        );

    \I__7844\ : CascadeMux
    port map (
            O => \N__37310\,
            I => \N__37302\
        );

    \I__7843\ : CascadeMux
    port map (
            O => \N__37309\,
            I => \N__37299\
        );

    \I__7842\ : CascadeMux
    port map (
            O => \N__37308\,
            I => \N__37292\
        );

    \I__7841\ : CascadeMux
    port map (
            O => \N__37307\,
            I => \N__37289\
        );

    \I__7840\ : CascadeMux
    port map (
            O => \N__37306\,
            I => \N__37285\
        );

    \I__7839\ : InMux
    port map (
            O => \N__37305\,
            I => \N__37281\
        );

    \I__7838\ : InMux
    port map (
            O => \N__37302\,
            I => \N__37278\
        );

    \I__7837\ : InMux
    port map (
            O => \N__37299\,
            I => \N__37273\
        );

    \I__7836\ : InMux
    port map (
            O => \N__37298\,
            I => \N__37273\
        );

    \I__7835\ : InMux
    port map (
            O => \N__37297\,
            I => \N__37268\
        );

    \I__7834\ : InMux
    port map (
            O => \N__37296\,
            I => \N__37268\
        );

    \I__7833\ : InMux
    port map (
            O => \N__37295\,
            I => \N__37265\
        );

    \I__7832\ : InMux
    port map (
            O => \N__37292\,
            I => \N__37262\
        );

    \I__7831\ : InMux
    port map (
            O => \N__37289\,
            I => \N__37253\
        );

    \I__7830\ : InMux
    port map (
            O => \N__37288\,
            I => \N__37253\
        );

    \I__7829\ : InMux
    port map (
            O => \N__37285\,
            I => \N__37253\
        );

    \I__7828\ : InMux
    port map (
            O => \N__37284\,
            I => \N__37253\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__37281\,
            I => \N__37246\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__37278\,
            I => \N__37246\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__37273\,
            I => \N__37246\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__37268\,
            I => \N__37241\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__37265\,
            I => \N__37241\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__37262\,
            I => \N__37238\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__37253\,
            I => \N__37235\
        );

    \I__7820\ : Span4Mux_v
    port map (
            O => \N__37246\,
            I => \N__37230\
        );

    \I__7819\ : Span4Mux_h
    port map (
            O => \N__37241\,
            I => \N__37230\
        );

    \I__7818\ : Odrv12
    port map (
            O => \N__37238\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__7817\ : Odrv12
    port map (
            O => \N__37235\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__7816\ : Odrv4
    port map (
            O => \N__37230\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__7815\ : InMux
    port map (
            O => \N__37223\,
            I => \N__37220\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__37220\,
            I => \N__37217\
        );

    \I__7813\ : Odrv4
    port map (
            O => \N__37217\,
            I => \pwm_generator_inst.un19_threshold_axb_1\
        );

    \I__7812\ : InMux
    port map (
            O => \N__37214\,
            I => \pwm_generator_inst.un15_threshold_1_cry_10\
        );

    \I__7811\ : InMux
    port map (
            O => \N__37211\,
            I => \N__37208\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__37208\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\
        );

    \I__7809\ : InMux
    port map (
            O => \N__37205\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11\
        );

    \I__7808\ : InMux
    port map (
            O => \N__37202\,
            I => \N__37199\
        );

    \I__7807\ : LocalMux
    port map (
            O => \N__37199\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\
        );

    \I__7806\ : InMux
    port map (
            O => \N__37196\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12\
        );

    \I__7805\ : InMux
    port map (
            O => \N__37193\,
            I => \N__37190\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__37190\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\
        );

    \I__7803\ : InMux
    port map (
            O => \N__37187\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13\
        );

    \I__7802\ : InMux
    port map (
            O => \N__37184\,
            I => \N__37181\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__37181\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\
        );

    \I__7800\ : InMux
    port map (
            O => \N__37178\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14\
        );

    \I__7799\ : InMux
    port map (
            O => \N__37175\,
            I => \N__37171\
        );

    \I__7798\ : InMux
    port map (
            O => \N__37174\,
            I => \N__37167\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__37171\,
            I => \N__37164\
        );

    \I__7796\ : InMux
    port map (
            O => \N__37170\,
            I => \N__37161\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__37167\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__7794\ : Odrv4
    port map (
            O => \N__37164\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__37161\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__7792\ : InMux
    port map (
            O => \N__37154\,
            I => \N__37151\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__37151\,
            I => \N__37148\
        );

    \I__7790\ : Odrv4
    port map (
            O => \N__37148\,
            I => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\
        );

    \I__7789\ : InMux
    port map (
            O => \N__37145\,
            I => \bfn_14_27_0_\
        );

    \I__7788\ : InMux
    port map (
            O => \N__37142\,
            I => \N__37139\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__37139\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\
        );

    \I__7786\ : InMux
    port map (
            O => \N__37136\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16\
        );

    \I__7785\ : InMux
    port map (
            O => \N__37133\,
            I => \N__37130\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__37130\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\
        );

    \I__7783\ : InMux
    port map (
            O => \N__37127\,
            I => \N__37124\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__37124\,
            I => \pwm_generator_inst.un15_threshold_1_axb_2\
        );

    \I__7781\ : InMux
    port map (
            O => \N__37121\,
            I => \N__37118\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__37118\,
            I => \N__37115\
        );

    \I__7779\ : Span4Mux_v
    port map (
            O => \N__37115\,
            I => \N__37112\
        );

    \I__7778\ : Span4Mux_h
    port map (
            O => \N__37112\,
            I => \N__37109\
        );

    \I__7777\ : Span4Mux_h
    port map (
            O => \N__37109\,
            I => \N__37106\
        );

    \I__7776\ : Odrv4
    port map (
            O => \N__37106\,
            I => \pwm_generator_inst.O_3\
        );

    \I__7775\ : InMux
    port map (
            O => \N__37103\,
            I => \N__37100\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__37100\,
            I => \pwm_generator_inst.un15_threshold_1_axb_3\
        );

    \I__7773\ : InMux
    port map (
            O => \N__37097\,
            I => \N__37094\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__37094\,
            I => \N__37091\
        );

    \I__7771\ : Span4Mux_v
    port map (
            O => \N__37091\,
            I => \N__37088\
        );

    \I__7770\ : Span4Mux_h
    port map (
            O => \N__37088\,
            I => \N__37085\
        );

    \I__7769\ : Span4Mux_h
    port map (
            O => \N__37085\,
            I => \N__37082\
        );

    \I__7768\ : Odrv4
    port map (
            O => \N__37082\,
            I => \pwm_generator_inst.O_4\
        );

    \I__7767\ : InMux
    port map (
            O => \N__37079\,
            I => \N__37076\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__37076\,
            I => \pwm_generator_inst.un15_threshold_1_axb_4\
        );

    \I__7765\ : InMux
    port map (
            O => \N__37073\,
            I => \N__37070\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__37070\,
            I => \N__37067\
        );

    \I__7763\ : Span4Mux_h
    port map (
            O => \N__37067\,
            I => \N__37064\
        );

    \I__7762\ : Span4Mux_h
    port map (
            O => \N__37064\,
            I => \N__37061\
        );

    \I__7761\ : Span4Mux_h
    port map (
            O => \N__37061\,
            I => \N__37058\
        );

    \I__7760\ : Odrv4
    port map (
            O => \N__37058\,
            I => \pwm_generator_inst.O_5\
        );

    \I__7759\ : InMux
    port map (
            O => \N__37055\,
            I => \N__37052\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__37052\,
            I => \pwm_generator_inst.un15_threshold_1_axb_5\
        );

    \I__7757\ : InMux
    port map (
            O => \N__37049\,
            I => \N__37046\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__37046\,
            I => \N__37043\
        );

    \I__7755\ : Span4Mux_h
    port map (
            O => \N__37043\,
            I => \N__37040\
        );

    \I__7754\ : Span4Mux_h
    port map (
            O => \N__37040\,
            I => \N__37037\
        );

    \I__7753\ : Span4Mux_h
    port map (
            O => \N__37037\,
            I => \N__37034\
        );

    \I__7752\ : Odrv4
    port map (
            O => \N__37034\,
            I => \pwm_generator_inst.O_6\
        );

    \I__7751\ : InMux
    port map (
            O => \N__37031\,
            I => \N__37028\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__37028\,
            I => \pwm_generator_inst.un15_threshold_1_axb_6\
        );

    \I__7749\ : InMux
    port map (
            O => \N__37025\,
            I => \N__37022\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__37022\,
            I => \N__37019\
        );

    \I__7747\ : Span12Mux_s7_v
    port map (
            O => \N__37019\,
            I => \N__37016\
        );

    \I__7746\ : Odrv12
    port map (
            O => \N__37016\,
            I => \pwm_generator_inst.O_7\
        );

    \I__7745\ : InMux
    port map (
            O => \N__37013\,
            I => \N__37010\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__37010\,
            I => \pwm_generator_inst.un15_threshold_1_axb_7\
        );

    \I__7743\ : InMux
    port map (
            O => \N__37007\,
            I => \N__37004\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__37004\,
            I => \N__37001\
        );

    \I__7741\ : Span4Mux_v
    port map (
            O => \N__37001\,
            I => \N__36998\
        );

    \I__7740\ : Span4Mux_h
    port map (
            O => \N__36998\,
            I => \N__36995\
        );

    \I__7739\ : Span4Mux_h
    port map (
            O => \N__36995\,
            I => \N__36992\
        );

    \I__7738\ : Odrv4
    port map (
            O => \N__36992\,
            I => \pwm_generator_inst.O_8\
        );

    \I__7737\ : InMux
    port map (
            O => \N__36989\,
            I => \N__36986\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__36986\,
            I => \pwm_generator_inst.un15_threshold_1_axb_8\
        );

    \I__7735\ : InMux
    port map (
            O => \N__36983\,
            I => \N__36980\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__36980\,
            I => \N__36977\
        );

    \I__7733\ : Span4Mux_h
    port map (
            O => \N__36977\,
            I => \N__36974\
        );

    \I__7732\ : Span4Mux_h
    port map (
            O => \N__36974\,
            I => \N__36971\
        );

    \I__7731\ : Span4Mux_h
    port map (
            O => \N__36971\,
            I => \N__36968\
        );

    \I__7730\ : Odrv4
    port map (
            O => \N__36968\,
            I => \pwm_generator_inst.O_9\
        );

    \I__7729\ : InMux
    port map (
            O => \N__36965\,
            I => \N__36962\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__36962\,
            I => \pwm_generator_inst.un15_threshold_1_axb_9\
        );

    \I__7727\ : CascadeMux
    port map (
            O => \N__36959\,
            I => \N__36955\
        );

    \I__7726\ : InMux
    port map (
            O => \N__36958\,
            I => \N__36951\
        );

    \I__7725\ : InMux
    port map (
            O => \N__36955\,
            I => \N__36948\
        );

    \I__7724\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36945\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__36951\,
            I => \N__36938\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__36948\,
            I => \N__36938\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__36945\,
            I => \N__36938\
        );

    \I__7720\ : Odrv4
    port map (
            O => \N__36938\,
            I => \il_max_comp1_D2\
        );

    \I__7719\ : InMux
    port map (
            O => \N__36935\,
            I => \N__36932\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__36932\,
            I => \N__36928\
        );

    \I__7717\ : InMux
    port map (
            O => \N__36931\,
            I => \N__36925\
        );

    \I__7716\ : Span4Mux_h
    port map (
            O => \N__36928\,
            I => \N__36922\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__36925\,
            I => \N__36919\
        );

    \I__7714\ : Span4Mux_h
    port map (
            O => \N__36922\,
            I => \N__36916\
        );

    \I__7713\ : Span4Mux_s3_h
    port map (
            O => \N__36919\,
            I => \N__36913\
        );

    \I__7712\ : Span4Mux_v
    port map (
            O => \N__36916\,
            I => \N__36908\
        );

    \I__7711\ : Span4Mux_h
    port map (
            O => \N__36913\,
            I => \N__36908\
        );

    \I__7710\ : Odrv4
    port map (
            O => \N__36908\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__7709\ : InMux
    port map (
            O => \N__36905\,
            I => \N__36902\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__36902\,
            I => \N__36898\
        );

    \I__7707\ : InMux
    port map (
            O => \N__36901\,
            I => \N__36895\
        );

    \I__7706\ : Span4Mux_h
    port map (
            O => \N__36898\,
            I => \N__36892\
        );

    \I__7705\ : LocalMux
    port map (
            O => \N__36895\,
            I => \N__36889\
        );

    \I__7704\ : Span4Mux_v
    port map (
            O => \N__36892\,
            I => \N__36886\
        );

    \I__7703\ : Span4Mux_s3_h
    port map (
            O => \N__36889\,
            I => \N__36883\
        );

    \I__7702\ : Span4Mux_v
    port map (
            O => \N__36886\,
            I => \N__36880\
        );

    \I__7701\ : Span4Mux_h
    port map (
            O => \N__36883\,
            I => \N__36877\
        );

    \I__7700\ : Odrv4
    port map (
            O => \N__36880\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__7699\ : Odrv4
    port map (
            O => \N__36877\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__7698\ : CascadeMux
    port map (
            O => \N__36872\,
            I => \N__36869\
        );

    \I__7697\ : InMux
    port map (
            O => \N__36869\,
            I => \N__36861\
        );

    \I__7696\ : InMux
    port map (
            O => \N__36868\,
            I => \N__36861\
        );

    \I__7695\ : InMux
    port map (
            O => \N__36867\,
            I => \N__36858\
        );

    \I__7694\ : InMux
    port map (
            O => \N__36866\,
            I => \N__36855\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__36861\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__36858\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__36855\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__7690\ : InMux
    port map (
            O => \N__36848\,
            I => \N__36842\
        );

    \I__7689\ : InMux
    port map (
            O => \N__36847\,
            I => \N__36835\
        );

    \I__7688\ : InMux
    port map (
            O => \N__36846\,
            I => \N__36835\
        );

    \I__7687\ : InMux
    port map (
            O => \N__36845\,
            I => \N__36835\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__36842\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__36835\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7684\ : InMux
    port map (
            O => \N__36830\,
            I => \N__36826\
        );

    \I__7683\ : InMux
    port map (
            O => \N__36829\,
            I => \N__36823\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__36826\,
            I => \N__36820\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__36823\,
            I => \N__36817\
        );

    \I__7680\ : Span4Mux_h
    port map (
            O => \N__36820\,
            I => \N__36814\
        );

    \I__7679\ : Span12Mux_v
    port map (
            O => \N__36817\,
            I => \N__36811\
        );

    \I__7678\ : Span4Mux_h
    port map (
            O => \N__36814\,
            I => \N__36808\
        );

    \I__7677\ : Odrv12
    port map (
            O => \N__36811\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__7676\ : Odrv4
    port map (
            O => \N__36808\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__7675\ : InMux
    port map (
            O => \N__36803\,
            I => \N__36800\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__36800\,
            I => \N__36797\
        );

    \I__7673\ : Span4Mux_h
    port map (
            O => \N__36797\,
            I => \N__36794\
        );

    \I__7672\ : Span4Mux_h
    port map (
            O => \N__36794\,
            I => \N__36791\
        );

    \I__7671\ : Span4Mux_h
    port map (
            O => \N__36791\,
            I => \N__36788\
        );

    \I__7670\ : Odrv4
    port map (
            O => \N__36788\,
            I => \pwm_generator_inst.O_0\
        );

    \I__7669\ : InMux
    port map (
            O => \N__36785\,
            I => \N__36782\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__36782\,
            I => \pwm_generator_inst.un15_threshold_1_axb_0\
        );

    \I__7667\ : InMux
    port map (
            O => \N__36779\,
            I => \N__36776\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__36776\,
            I => \N__36773\
        );

    \I__7665\ : Span4Mux_h
    port map (
            O => \N__36773\,
            I => \N__36770\
        );

    \I__7664\ : Span4Mux_h
    port map (
            O => \N__36770\,
            I => \N__36767\
        );

    \I__7663\ : Span4Mux_h
    port map (
            O => \N__36767\,
            I => \N__36764\
        );

    \I__7662\ : Odrv4
    port map (
            O => \N__36764\,
            I => \pwm_generator_inst.O_1\
        );

    \I__7661\ : InMux
    port map (
            O => \N__36761\,
            I => \N__36758\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__36758\,
            I => \pwm_generator_inst.un15_threshold_1_axb_1\
        );

    \I__7659\ : InMux
    port map (
            O => \N__36755\,
            I => \N__36752\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__36752\,
            I => \N__36749\
        );

    \I__7657\ : Span12Mux_h
    port map (
            O => \N__36749\,
            I => \N__36746\
        );

    \I__7656\ : Odrv12
    port map (
            O => \N__36746\,
            I => \pwm_generator_inst.O_2\
        );

    \I__7655\ : InMux
    port map (
            O => \N__36743\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__7654\ : InMux
    port map (
            O => \N__36740\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__7653\ : InMux
    port map (
            O => \N__36737\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__7652\ : InMux
    port map (
            O => \N__36734\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__7651\ : InMux
    port map (
            O => \N__36731\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__7650\ : InMux
    port map (
            O => \N__36728\,
            I => \N__36690\
        );

    \I__7649\ : InMux
    port map (
            O => \N__36727\,
            I => \N__36690\
        );

    \I__7648\ : InMux
    port map (
            O => \N__36726\,
            I => \N__36690\
        );

    \I__7647\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36690\
        );

    \I__7646\ : InMux
    port map (
            O => \N__36724\,
            I => \N__36681\
        );

    \I__7645\ : InMux
    port map (
            O => \N__36723\,
            I => \N__36681\
        );

    \I__7644\ : InMux
    port map (
            O => \N__36722\,
            I => \N__36681\
        );

    \I__7643\ : InMux
    port map (
            O => \N__36721\,
            I => \N__36681\
        );

    \I__7642\ : InMux
    port map (
            O => \N__36720\,
            I => \N__36672\
        );

    \I__7641\ : InMux
    port map (
            O => \N__36719\,
            I => \N__36672\
        );

    \I__7640\ : InMux
    port map (
            O => \N__36718\,
            I => \N__36672\
        );

    \I__7639\ : InMux
    port map (
            O => \N__36717\,
            I => \N__36672\
        );

    \I__7638\ : InMux
    port map (
            O => \N__36716\,
            I => \N__36663\
        );

    \I__7637\ : InMux
    port map (
            O => \N__36715\,
            I => \N__36663\
        );

    \I__7636\ : InMux
    port map (
            O => \N__36714\,
            I => \N__36663\
        );

    \I__7635\ : InMux
    port map (
            O => \N__36713\,
            I => \N__36663\
        );

    \I__7634\ : InMux
    port map (
            O => \N__36712\,
            I => \N__36654\
        );

    \I__7633\ : InMux
    port map (
            O => \N__36711\,
            I => \N__36654\
        );

    \I__7632\ : InMux
    port map (
            O => \N__36710\,
            I => \N__36654\
        );

    \I__7631\ : InMux
    port map (
            O => \N__36709\,
            I => \N__36654\
        );

    \I__7630\ : InMux
    port map (
            O => \N__36708\,
            I => \N__36649\
        );

    \I__7629\ : InMux
    port map (
            O => \N__36707\,
            I => \N__36649\
        );

    \I__7628\ : InMux
    port map (
            O => \N__36706\,
            I => \N__36640\
        );

    \I__7627\ : InMux
    port map (
            O => \N__36705\,
            I => \N__36640\
        );

    \I__7626\ : InMux
    port map (
            O => \N__36704\,
            I => \N__36640\
        );

    \I__7625\ : InMux
    port map (
            O => \N__36703\,
            I => \N__36640\
        );

    \I__7624\ : InMux
    port map (
            O => \N__36702\,
            I => \N__36631\
        );

    \I__7623\ : InMux
    port map (
            O => \N__36701\,
            I => \N__36631\
        );

    \I__7622\ : InMux
    port map (
            O => \N__36700\,
            I => \N__36631\
        );

    \I__7621\ : InMux
    port map (
            O => \N__36699\,
            I => \N__36631\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__36690\,
            I => \N__36626\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__36681\,
            I => \N__36626\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__36672\,
            I => \N__36619\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__36663\,
            I => \N__36619\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__36654\,
            I => \N__36619\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__36649\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__36640\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__36631\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7612\ : Odrv4
    port map (
            O => \N__36626\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7611\ : Odrv12
    port map (
            O => \N__36619\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__7610\ : CEMux
    port map (
            O => \N__36608\,
            I => \N__36602\
        );

    \I__7609\ : CEMux
    port map (
            O => \N__36607\,
            I => \N__36598\
        );

    \I__7608\ : CEMux
    port map (
            O => \N__36606\,
            I => \N__36590\
        );

    \I__7607\ : CEMux
    port map (
            O => \N__36605\,
            I => \N__36587\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__36602\,
            I => \N__36584\
        );

    \I__7605\ : CEMux
    port map (
            O => \N__36601\,
            I => \N__36581\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__36598\,
            I => \N__36555\
        );

    \I__7603\ : CEMux
    port map (
            O => \N__36597\,
            I => \N__36552\
        );

    \I__7602\ : CEMux
    port map (
            O => \N__36596\,
            I => \N__36549\
        );

    \I__7601\ : CEMux
    port map (
            O => \N__36595\,
            I => \N__36539\
        );

    \I__7600\ : CEMux
    port map (
            O => \N__36594\,
            I => \N__36535\
        );

    \I__7599\ : CEMux
    port map (
            O => \N__36593\,
            I => \N__36532\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__36590\,
            I => \N__36522\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__36587\,
            I => \N__36522\
        );

    \I__7596\ : Span4Mux_v
    port map (
            O => \N__36584\,
            I => \N__36522\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__36581\,
            I => \N__36522\
        );

    \I__7594\ : InMux
    port map (
            O => \N__36580\,
            I => \N__36513\
        );

    \I__7593\ : InMux
    port map (
            O => \N__36579\,
            I => \N__36513\
        );

    \I__7592\ : InMux
    port map (
            O => \N__36578\,
            I => \N__36513\
        );

    \I__7591\ : InMux
    port map (
            O => \N__36577\,
            I => \N__36513\
        );

    \I__7590\ : InMux
    port map (
            O => \N__36576\,
            I => \N__36506\
        );

    \I__7589\ : InMux
    port map (
            O => \N__36575\,
            I => \N__36506\
        );

    \I__7588\ : InMux
    port map (
            O => \N__36574\,
            I => \N__36506\
        );

    \I__7587\ : InMux
    port map (
            O => \N__36573\,
            I => \N__36497\
        );

    \I__7586\ : InMux
    port map (
            O => \N__36572\,
            I => \N__36497\
        );

    \I__7585\ : InMux
    port map (
            O => \N__36571\,
            I => \N__36497\
        );

    \I__7584\ : InMux
    port map (
            O => \N__36570\,
            I => \N__36497\
        );

    \I__7583\ : InMux
    port map (
            O => \N__36569\,
            I => \N__36488\
        );

    \I__7582\ : InMux
    port map (
            O => \N__36568\,
            I => \N__36488\
        );

    \I__7581\ : InMux
    port map (
            O => \N__36567\,
            I => \N__36488\
        );

    \I__7580\ : InMux
    port map (
            O => \N__36566\,
            I => \N__36488\
        );

    \I__7579\ : InMux
    port map (
            O => \N__36565\,
            I => \N__36479\
        );

    \I__7578\ : InMux
    port map (
            O => \N__36564\,
            I => \N__36479\
        );

    \I__7577\ : InMux
    port map (
            O => \N__36563\,
            I => \N__36479\
        );

    \I__7576\ : InMux
    port map (
            O => \N__36562\,
            I => \N__36479\
        );

    \I__7575\ : InMux
    port map (
            O => \N__36561\,
            I => \N__36470\
        );

    \I__7574\ : InMux
    port map (
            O => \N__36560\,
            I => \N__36470\
        );

    \I__7573\ : InMux
    port map (
            O => \N__36559\,
            I => \N__36470\
        );

    \I__7572\ : InMux
    port map (
            O => \N__36558\,
            I => \N__36470\
        );

    \I__7571\ : Span4Mux_v
    port map (
            O => \N__36555\,
            I => \N__36464\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__36552\,
            I => \N__36464\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__36549\,
            I => \N__36461\
        );

    \I__7568\ : InMux
    port map (
            O => \N__36548\,
            I => \N__36454\
        );

    \I__7567\ : InMux
    port map (
            O => \N__36547\,
            I => \N__36454\
        );

    \I__7566\ : InMux
    port map (
            O => \N__36546\,
            I => \N__36454\
        );

    \I__7565\ : InMux
    port map (
            O => \N__36545\,
            I => \N__36445\
        );

    \I__7564\ : InMux
    port map (
            O => \N__36544\,
            I => \N__36445\
        );

    \I__7563\ : InMux
    port map (
            O => \N__36543\,
            I => \N__36445\
        );

    \I__7562\ : InMux
    port map (
            O => \N__36542\,
            I => \N__36445\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__36539\,
            I => \N__36441\
        );

    \I__7560\ : CEMux
    port map (
            O => \N__36538\,
            I => \N__36438\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__36535\,
            I => \N__36435\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__36532\,
            I => \N__36432\
        );

    \I__7557\ : CEMux
    port map (
            O => \N__36531\,
            I => \N__36429\
        );

    \I__7556\ : Span4Mux_v
    port map (
            O => \N__36522\,
            I => \N__36426\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__36513\,
            I => \N__36417\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__36506\,
            I => \N__36417\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__36497\,
            I => \N__36417\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__36488\,
            I => \N__36417\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__36479\,
            I => \N__36412\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__36470\,
            I => \N__36412\
        );

    \I__7549\ : InMux
    port map (
            O => \N__36469\,
            I => \N__36409\
        );

    \I__7548\ : Span4Mux_h
    port map (
            O => \N__36464\,
            I => \N__36404\
        );

    \I__7547\ : Span4Mux_v
    port map (
            O => \N__36461\,
            I => \N__36404\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__36454\,
            I => \N__36399\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__36445\,
            I => \N__36399\
        );

    \I__7544\ : CEMux
    port map (
            O => \N__36444\,
            I => \N__36396\
        );

    \I__7543\ : Span4Mux_h
    port map (
            O => \N__36441\,
            I => \N__36393\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__36438\,
            I => \N__36386\
        );

    \I__7541\ : Span4Mux_v
    port map (
            O => \N__36435\,
            I => \N__36386\
        );

    \I__7540\ : Span4Mux_h
    port map (
            O => \N__36432\,
            I => \N__36386\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__36429\,
            I => \N__36383\
        );

    \I__7538\ : Span4Mux_v
    port map (
            O => \N__36426\,
            I => \N__36380\
        );

    \I__7537\ : Span4Mux_v
    port map (
            O => \N__36417\,
            I => \N__36375\
        );

    \I__7536\ : Span4Mux_v
    port map (
            O => \N__36412\,
            I => \N__36375\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__36409\,
            I => \N__36372\
        );

    \I__7534\ : Span4Mux_h
    port map (
            O => \N__36404\,
            I => \N__36367\
        );

    \I__7533\ : Span4Mux_h
    port map (
            O => \N__36399\,
            I => \N__36367\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__36396\,
            I => \N__36364\
        );

    \I__7531\ : Span4Mux_h
    port map (
            O => \N__36393\,
            I => \N__36357\
        );

    \I__7530\ : Span4Mux_v
    port map (
            O => \N__36386\,
            I => \N__36357\
        );

    \I__7529\ : Span4Mux_v
    port map (
            O => \N__36383\,
            I => \N__36357\
        );

    \I__7528\ : Span4Mux_h
    port map (
            O => \N__36380\,
            I => \N__36354\
        );

    \I__7527\ : Span4Mux_v
    port map (
            O => \N__36375\,
            I => \N__36351\
        );

    \I__7526\ : Span4Mux_h
    port map (
            O => \N__36372\,
            I => \N__36346\
        );

    \I__7525\ : Span4Mux_v
    port map (
            O => \N__36367\,
            I => \N__36346\
        );

    \I__7524\ : Span12Mux_h
    port map (
            O => \N__36364\,
            I => \N__36341\
        );

    \I__7523\ : Sp12to4
    port map (
            O => \N__36357\,
            I => \N__36341\
        );

    \I__7522\ : Span4Mux_h
    port map (
            O => \N__36354\,
            I => \N__36338\
        );

    \I__7521\ : Span4Mux_v
    port map (
            O => \N__36351\,
            I => \N__36335\
        );

    \I__7520\ : Span4Mux_v
    port map (
            O => \N__36346\,
            I => \N__36332\
        );

    \I__7519\ : Odrv12
    port map (
            O => \N__36341\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__7518\ : Odrv4
    port map (
            O => \N__36338\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__7517\ : Odrv4
    port map (
            O => \N__36335\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__7516\ : Odrv4
    port map (
            O => \N__36332\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__7515\ : InMux
    port map (
            O => \N__36323\,
            I => \N__36320\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__36320\,
            I => \N__36317\
        );

    \I__7513\ : Span4Mux_v
    port map (
            O => \N__36317\,
            I => \N__36313\
        );

    \I__7512\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36310\
        );

    \I__7511\ : Span4Mux_h
    port map (
            O => \N__36313\,
            I => \N__36307\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__36310\,
            I => \N__36304\
        );

    \I__7509\ : Span4Mux_h
    port map (
            O => \N__36307\,
            I => \N__36301\
        );

    \I__7508\ : Span12Mux_v
    port map (
            O => \N__36304\,
            I => \N__36298\
        );

    \I__7507\ : Odrv4
    port map (
            O => \N__36301\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__7506\ : Odrv12
    port map (
            O => \N__36298\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__7505\ : InMux
    port map (
            O => \N__36293\,
            I => \N__36290\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__36290\,
            I => \N__36287\
        );

    \I__7503\ : Span4Mux_v
    port map (
            O => \N__36287\,
            I => \N__36284\
        );

    \I__7502\ : Span4Mux_v
    port map (
            O => \N__36284\,
            I => \N__36280\
        );

    \I__7501\ : InMux
    port map (
            O => \N__36283\,
            I => \N__36277\
        );

    \I__7500\ : Span4Mux_v
    port map (
            O => \N__36280\,
            I => \N__36274\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__36277\,
            I => state_ns_i_a3_1
        );

    \I__7498\ : Odrv4
    port map (
            O => \N__36274\,
            I => state_ns_i_a3_1
        );

    \I__7497\ : InMux
    port map (
            O => \N__36269\,
            I => \bfn_14_16_0_\
        );

    \I__7496\ : InMux
    port map (
            O => \N__36266\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__7495\ : InMux
    port map (
            O => \N__36263\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__7494\ : InMux
    port map (
            O => \N__36260\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__7493\ : InMux
    port map (
            O => \N__36257\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__7492\ : InMux
    port map (
            O => \N__36254\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__7491\ : InMux
    port map (
            O => \N__36251\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__7490\ : InMux
    port map (
            O => \N__36248\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__7489\ : InMux
    port map (
            O => \N__36245\,
            I => \bfn_14_17_0_\
        );

    \I__7488\ : InMux
    port map (
            O => \N__36242\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__7487\ : InMux
    port map (
            O => \N__36239\,
            I => \bfn_14_15_0_\
        );

    \I__7486\ : InMux
    port map (
            O => \N__36236\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__7485\ : InMux
    port map (
            O => \N__36233\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__7484\ : InMux
    port map (
            O => \N__36230\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__7483\ : InMux
    port map (
            O => \N__36227\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__7482\ : InMux
    port map (
            O => \N__36224\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__7481\ : InMux
    port map (
            O => \N__36221\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__7480\ : InMux
    port map (
            O => \N__36218\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36215\,
            I => \N__36209\
        );

    \I__7478\ : InMux
    port map (
            O => \N__36214\,
            I => \N__36202\
        );

    \I__7477\ : InMux
    port map (
            O => \N__36213\,
            I => \N__36202\
        );

    \I__7476\ : InMux
    port map (
            O => \N__36212\,
            I => \N__36202\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__36209\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__36202\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__7473\ : InMux
    port map (
            O => \N__36197\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__7472\ : InMux
    port map (
            O => \N__36194\,
            I => \N__36160\
        );

    \I__7471\ : InMux
    port map (
            O => \N__36193\,
            I => \N__36160\
        );

    \I__7470\ : InMux
    port map (
            O => \N__36192\,
            I => \N__36160\
        );

    \I__7469\ : InMux
    port map (
            O => \N__36191\,
            I => \N__36160\
        );

    \I__7468\ : InMux
    port map (
            O => \N__36190\,
            I => \N__36151\
        );

    \I__7467\ : InMux
    port map (
            O => \N__36189\,
            I => \N__36151\
        );

    \I__7466\ : InMux
    port map (
            O => \N__36188\,
            I => \N__36151\
        );

    \I__7465\ : InMux
    port map (
            O => \N__36187\,
            I => \N__36151\
        );

    \I__7464\ : InMux
    port map (
            O => \N__36186\,
            I => \N__36142\
        );

    \I__7463\ : InMux
    port map (
            O => \N__36185\,
            I => \N__36142\
        );

    \I__7462\ : InMux
    port map (
            O => \N__36184\,
            I => \N__36142\
        );

    \I__7461\ : InMux
    port map (
            O => \N__36183\,
            I => \N__36142\
        );

    \I__7460\ : InMux
    port map (
            O => \N__36182\,
            I => \N__36135\
        );

    \I__7459\ : InMux
    port map (
            O => \N__36181\,
            I => \N__36135\
        );

    \I__7458\ : InMux
    port map (
            O => \N__36180\,
            I => \N__36135\
        );

    \I__7457\ : InMux
    port map (
            O => \N__36179\,
            I => \N__36126\
        );

    \I__7456\ : InMux
    port map (
            O => \N__36178\,
            I => \N__36126\
        );

    \I__7455\ : InMux
    port map (
            O => \N__36177\,
            I => \N__36126\
        );

    \I__7454\ : InMux
    port map (
            O => \N__36176\,
            I => \N__36126\
        );

    \I__7453\ : InMux
    port map (
            O => \N__36175\,
            I => \N__36113\
        );

    \I__7452\ : InMux
    port map (
            O => \N__36174\,
            I => \N__36113\
        );

    \I__7451\ : InMux
    port map (
            O => \N__36173\,
            I => \N__36113\
        );

    \I__7450\ : InMux
    port map (
            O => \N__36172\,
            I => \N__36104\
        );

    \I__7449\ : InMux
    port map (
            O => \N__36171\,
            I => \N__36104\
        );

    \I__7448\ : InMux
    port map (
            O => \N__36170\,
            I => \N__36104\
        );

    \I__7447\ : InMux
    port map (
            O => \N__36169\,
            I => \N__36104\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__36160\,
            I => \N__36093\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__36151\,
            I => \N__36093\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__36142\,
            I => \N__36093\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__36135\,
            I => \N__36093\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__36126\,
            I => \N__36093\
        );

    \I__7441\ : IoInMux
    port map (
            O => \N__36125\,
            I => \N__36090\
        );

    \I__7440\ : InMux
    port map (
            O => \N__36124\,
            I => \N__36081\
        );

    \I__7439\ : InMux
    port map (
            O => \N__36123\,
            I => \N__36081\
        );

    \I__7438\ : InMux
    port map (
            O => \N__36122\,
            I => \N__36081\
        );

    \I__7437\ : InMux
    port map (
            O => \N__36121\,
            I => \N__36081\
        );

    \I__7436\ : InMux
    port map (
            O => \N__36120\,
            I => \N__36078\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__36113\,
            I => \N__36071\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__36104\,
            I => \N__36071\
        );

    \I__7433\ : Span4Mux_v
    port map (
            O => \N__36093\,
            I => \N__36071\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__36090\,
            I => \N__36068\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__36081\,
            I => \N__36065\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__36078\,
            I => \N__36060\
        );

    \I__7429\ : Span4Mux_v
    port map (
            O => \N__36071\,
            I => \N__36060\
        );

    \I__7428\ : IoSpan4Mux
    port map (
            O => \N__36068\,
            I => \N__36057\
        );

    \I__7427\ : Odrv12
    port map (
            O => \N__36065\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__7426\ : Odrv4
    port map (
            O => \N__36060\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__7425\ : Odrv4
    port map (
            O => \N__36057\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__7424\ : InMux
    port map (
            O => \N__36050\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__7423\ : CascadeMux
    port map (
            O => \N__36047\,
            I => \N__36042\
        );

    \I__7422\ : CascadeMux
    port map (
            O => \N__36046\,
            I => \N__36038\
        );

    \I__7421\ : InMux
    port map (
            O => \N__36045\,
            I => \N__36035\
        );

    \I__7420\ : InMux
    port map (
            O => \N__36042\,
            I => \N__36028\
        );

    \I__7419\ : InMux
    port map (
            O => \N__36041\,
            I => \N__36028\
        );

    \I__7418\ : InMux
    port map (
            O => \N__36038\,
            I => \N__36028\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__36035\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__36028\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__7415\ : InMux
    port map (
            O => \N__36023\,
            I => \bfn_14_14_0_\
        );

    \I__7414\ : InMux
    port map (
            O => \N__36020\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__7413\ : InMux
    port map (
            O => \N__36017\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__7412\ : InMux
    port map (
            O => \N__36014\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__7411\ : InMux
    port map (
            O => \N__36011\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__7410\ : InMux
    port map (
            O => \N__36008\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__7409\ : InMux
    port map (
            O => \N__36005\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__7408\ : InMux
    port map (
            O => \N__36002\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__7407\ : InMux
    port map (
            O => \N__35999\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__7406\ : InMux
    port map (
            O => \N__35996\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__7405\ : InMux
    port map (
            O => \N__35993\,
            I => \bfn_14_13_0_\
        );

    \I__7404\ : InMux
    port map (
            O => \N__35990\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__7403\ : InMux
    port map (
            O => \N__35987\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__7402\ : CascadeMux
    port map (
            O => \N__35984\,
            I => \N__35979\
        );

    \I__7401\ : InMux
    port map (
            O => \N__35983\,
            I => \N__35976\
        );

    \I__7400\ : InMux
    port map (
            O => \N__35982\,
            I => \N__35971\
        );

    \I__7399\ : InMux
    port map (
            O => \N__35979\,
            I => \N__35971\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__35976\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__35971\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__7396\ : InMux
    port map (
            O => \N__35966\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__7395\ : CascadeMux
    port map (
            O => \N__35963\,
            I => \N__35959\
        );

    \I__7394\ : InMux
    port map (
            O => \N__35962\,
            I => \N__35955\
        );

    \I__7393\ : InMux
    port map (
            O => \N__35959\,
            I => \N__35952\
        );

    \I__7392\ : InMux
    port map (
            O => \N__35958\,
            I => \N__35949\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__35955\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__35952\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__7389\ : LocalMux
    port map (
            O => \N__35949\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__7388\ : InMux
    port map (
            O => \N__35942\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__7387\ : InMux
    port map (
            O => \N__35939\,
            I => \N__35935\
        );

    \I__7386\ : InMux
    port map (
            O => \N__35938\,
            I => \N__35932\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__35935\,
            I => \N__35929\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__35932\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7383\ : Odrv4
    port map (
            O => \N__35929\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7382\ : InMux
    port map (
            O => \N__35924\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__7381\ : InMux
    port map (
            O => \N__35921\,
            I => \N__35917\
        );

    \I__7380\ : InMux
    port map (
            O => \N__35920\,
            I => \N__35914\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__35917\,
            I => \N__35911\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__35914\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7377\ : Odrv4
    port map (
            O => \N__35911\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__7376\ : InMux
    port map (
            O => \N__35906\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__7375\ : InMux
    port map (
            O => \N__35903\,
            I => \N__35899\
        );

    \I__7374\ : InMux
    port map (
            O => \N__35902\,
            I => \N__35896\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__35899\,
            I => \N__35893\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__35896\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7371\ : Odrv12
    port map (
            O => \N__35893\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__7370\ : InMux
    port map (
            O => \N__35888\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__7369\ : CascadeMux
    port map (
            O => \N__35885\,
            I => \N__35880\
        );

    \I__7368\ : InMux
    port map (
            O => \N__35884\,
            I => \N__35877\
        );

    \I__7367\ : InMux
    port map (
            O => \N__35883\,
            I => \N__35872\
        );

    \I__7366\ : InMux
    port map (
            O => \N__35880\,
            I => \N__35872\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__35877\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__35872\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__7363\ : InMux
    port map (
            O => \N__35867\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__7362\ : InMux
    port map (
            O => \N__35864\,
            I => \N__35859\
        );

    \I__7361\ : InMux
    port map (
            O => \N__35863\,
            I => \N__35856\
        );

    \I__7360\ : InMux
    port map (
            O => \N__35862\,
            I => \N__35853\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__35859\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__35856\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__35853\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__7356\ : InMux
    port map (
            O => \N__35846\,
            I => \bfn_14_12_0_\
        );

    \I__7355\ : InMux
    port map (
            O => \N__35843\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__7354\ : InMux
    port map (
            O => \N__35840\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__7353\ : InMux
    port map (
            O => \N__35837\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__7352\ : InMux
    port map (
            O => \N__35834\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__7351\ : InMux
    port map (
            O => \N__35831\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__7350\ : InMux
    port map (
            O => \N__35828\,
            I => \N__35825\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__35825\,
            I => \N__35821\
        );

    \I__7348\ : InMux
    port map (
            O => \N__35824\,
            I => \N__35818\
        );

    \I__7347\ : Span4Mux_v
    port map (
            O => \N__35821\,
            I => \N__35815\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__35818\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7345\ : Odrv4
    port map (
            O => \N__35815\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__7344\ : InMux
    port map (
            O => \N__35810\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__7343\ : InMux
    port map (
            O => \N__35807\,
            I => \N__35803\
        );

    \I__7342\ : InMux
    port map (
            O => \N__35806\,
            I => \N__35800\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__35803\,
            I => \N__35797\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__35800\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7339\ : Odrv4
    port map (
            O => \N__35797\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7338\ : InMux
    port map (
            O => \N__35792\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__7337\ : InMux
    port map (
            O => \N__35789\,
            I => \N__35785\
        );

    \I__7336\ : InMux
    port map (
            O => \N__35788\,
            I => \N__35782\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__35785\,
            I => \N__35779\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__35782\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7333\ : Odrv12
    port map (
            O => \N__35779\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7332\ : InMux
    port map (
            O => \N__35774\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__7331\ : InMux
    port map (
            O => \N__35771\,
            I => \N__35767\
        );

    \I__7330\ : InMux
    port map (
            O => \N__35770\,
            I => \N__35764\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__35767\,
            I => \N__35761\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__35764\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7327\ : Odrv12
    port map (
            O => \N__35761\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7326\ : InMux
    port map (
            O => \N__35756\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__7325\ : InMux
    port map (
            O => \N__35753\,
            I => \N__35749\
        );

    \I__7324\ : InMux
    port map (
            O => \N__35752\,
            I => \N__35746\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__35749\,
            I => \N__35743\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__35746\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7321\ : Odrv4
    port map (
            O => \N__35743\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7320\ : InMux
    port map (
            O => \N__35738\,
            I => \bfn_14_11_0_\
        );

    \I__7319\ : InMux
    port map (
            O => \N__35735\,
            I => \N__35731\
        );

    \I__7318\ : InMux
    port map (
            O => \N__35734\,
            I => \N__35728\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__35731\,
            I => \N__35725\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__35728\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7315\ : Odrv4
    port map (
            O => \N__35725\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7314\ : InMux
    port map (
            O => \N__35720\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__7313\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35713\
        );

    \I__7312\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35710\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__35713\,
            I => \N__35707\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__35710\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7309\ : Odrv4
    port map (
            O => \N__35707\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7308\ : InMux
    port map (
            O => \N__35702\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__7307\ : InMux
    port map (
            O => \N__35699\,
            I => \N__35695\
        );

    \I__7306\ : InMux
    port map (
            O => \N__35698\,
            I => \N__35692\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__35695\,
            I => \N__35689\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__35692\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7303\ : Odrv4
    port map (
            O => \N__35689\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__7302\ : InMux
    port map (
            O => \N__35684\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__7301\ : InMux
    port map (
            O => \N__35681\,
            I => \N__35678\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__35678\,
            I => \N__35675\
        );

    \I__7299\ : Span4Mux_h
    port map (
            O => \N__35675\,
            I => \N__35672\
        );

    \I__7298\ : Odrv4
    port map (
            O => \N__35672\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt28\
        );

    \I__7297\ : CascadeMux
    port map (
            O => \N__35669\,
            I => \N__35666\
        );

    \I__7296\ : InMux
    port map (
            O => \N__35666\,
            I => \N__35663\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__35663\,
            I => \N__35660\
        );

    \I__7294\ : Span4Mux_h
    port map (
            O => \N__35660\,
            I => \N__35657\
        );

    \I__7293\ : Odrv4
    port map (
            O => \N__35657\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\
        );

    \I__7292\ : InMux
    port map (
            O => \N__35654\,
            I => \N__35651\
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__35651\,
            I => \N__35648\
        );

    \I__7290\ : Span4Mux_v
    port map (
            O => \N__35648\,
            I => \N__35645\
        );

    \I__7289\ : Odrv4
    port map (
            O => \N__35645\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\
        );

    \I__7288\ : CascadeMux
    port map (
            O => \N__35642\,
            I => \N__35639\
        );

    \I__7287\ : InMux
    port map (
            O => \N__35639\,
            I => \N__35635\
        );

    \I__7286\ : CascadeMux
    port map (
            O => \N__35638\,
            I => \N__35632\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__35635\,
            I => \N__35629\
        );

    \I__7284\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35626\
        );

    \I__7283\ : Span4Mux_v
    port map (
            O => \N__35629\,
            I => \N__35623\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__35626\,
            I => \N__35620\
        );

    \I__7281\ : Odrv4
    port map (
            O => \N__35623\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt30\
        );

    \I__7280\ : Odrv12
    port map (
            O => \N__35620\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt30\
        );

    \I__7279\ : InMux
    port map (
            O => \N__35615\,
            I => \N__35612\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__35612\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\
        );

    \I__7277\ : InMux
    port map (
            O => \N__35609\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_28\
        );

    \I__7276\ : InMux
    port map (
            O => \N__35606\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30\
        );

    \I__7275\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35600\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__35600\,
            I => \N__35596\
        );

    \I__7273\ : InMux
    port map (
            O => \N__35599\,
            I => \N__35593\
        );

    \I__7272\ : Span4Mux_v
    port map (
            O => \N__35596\,
            I => \N__35590\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__35593\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__7270\ : Odrv4
    port map (
            O => \N__35590\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__7269\ : InMux
    port map (
            O => \N__35585\,
            I => \N__35582\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__35582\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\
        );

    \I__7267\ : CascadeMux
    port map (
            O => \N__35579\,
            I => \N__35575\
        );

    \I__7266\ : CascadeMux
    port map (
            O => \N__35578\,
            I => \N__35572\
        );

    \I__7265\ : InMux
    port map (
            O => \N__35575\,
            I => \N__35569\
        );

    \I__7264\ : InMux
    port map (
            O => \N__35572\,
            I => \N__35565\
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__35569\,
            I => \N__35562\
        );

    \I__7262\ : InMux
    port map (
            O => \N__35568\,
            I => \N__35559\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__35565\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7260\ : Odrv12
    port map (
            O => \N__35562\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__35559\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__7258\ : InMux
    port map (
            O => \N__35552\,
            I => \N__35548\
        );

    \I__7257\ : InMux
    port map (
            O => \N__35551\,
            I => \N__35545\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__35548\,
            I => \N__35542\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__35545\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7254\ : Odrv4
    port map (
            O => \N__35542\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__7253\ : InMux
    port map (
            O => \N__35537\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__7252\ : CascadeMux
    port map (
            O => \N__35534\,
            I => \N__35531\
        );

    \I__7251\ : InMux
    port map (
            O => \N__35531\,
            I => \N__35528\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__35528\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28\
        );

    \I__7249\ : InMux
    port map (
            O => \N__35525\,
            I => \N__35521\
        );

    \I__7248\ : InMux
    port map (
            O => \N__35524\,
            I => \N__35518\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__35521\,
            I => \N__35515\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__35518\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7245\ : Odrv4
    port map (
            O => \N__35515\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__7244\ : InMux
    port map (
            O => \N__35510\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__7243\ : InMux
    port map (
            O => \N__35507\,
            I => \N__35503\
        );

    \I__7242\ : InMux
    port map (
            O => \N__35506\,
            I => \N__35500\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__35503\,
            I => \N__35497\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__35500\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7239\ : Odrv4
    port map (
            O => \N__35497\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__7238\ : CascadeMux
    port map (
            O => \N__35492\,
            I => \N__35489\
        );

    \I__7237\ : InMux
    port map (
            O => \N__35489\,
            I => \N__35486\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__35486\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__7235\ : InMux
    port map (
            O => \N__35483\,
            I => \N__35480\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__35480\,
            I => \N__35477\
        );

    \I__7233\ : Span4Mux_h
    port map (
            O => \N__35477\,
            I => \N__35474\
        );

    \I__7232\ : Span4Mux_v
    port map (
            O => \N__35474\,
            I => \N__35471\
        );

    \I__7231\ : Odrv4
    port map (
            O => \N__35471\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__7230\ : CascadeMux
    port map (
            O => \N__35468\,
            I => \N__35465\
        );

    \I__7229\ : InMux
    port map (
            O => \N__35465\,
            I => \N__35462\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__35462\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__7227\ : InMux
    port map (
            O => \N__35459\,
            I => \N__35456\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__35456\,
            I => \N__35453\
        );

    \I__7225\ : Span4Mux_v
    port map (
            O => \N__35453\,
            I => \N__35450\
        );

    \I__7224\ : Odrv4
    port map (
            O => \N__35450\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__7223\ : CascadeMux
    port map (
            O => \N__35447\,
            I => \N__35444\
        );

    \I__7222\ : InMux
    port map (
            O => \N__35444\,
            I => \N__35441\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__35441\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__7220\ : InMux
    port map (
            O => \N__35438\,
            I => \N__35435\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__35435\,
            I => \N__35432\
        );

    \I__7218\ : Span4Mux_h
    port map (
            O => \N__35432\,
            I => \N__35429\
        );

    \I__7217\ : Odrv4
    port map (
            O => \N__35429\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__7216\ : CascadeMux
    port map (
            O => \N__35426\,
            I => \N__35423\
        );

    \I__7215\ : InMux
    port map (
            O => \N__35423\,
            I => \N__35420\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__35420\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__7213\ : InMux
    port map (
            O => \N__35417\,
            I => \N__35414\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__35414\,
            I => \N__35411\
        );

    \I__7211\ : Odrv4
    port map (
            O => \N__35411\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt16\
        );

    \I__7210\ : CascadeMux
    port map (
            O => \N__35408\,
            I => \N__35405\
        );

    \I__7209\ : InMux
    port map (
            O => \N__35405\,
            I => \N__35402\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__35402\,
            I => \N__35399\
        );

    \I__7207\ : Span4Mux_h
    port map (
            O => \N__35399\,
            I => \N__35396\
        );

    \I__7206\ : Odrv4
    port map (
            O => \N__35396\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\
        );

    \I__7205\ : CascadeMux
    port map (
            O => \N__35393\,
            I => \N__35390\
        );

    \I__7204\ : InMux
    port map (
            O => \N__35390\,
            I => \N__35387\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__35387\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__7202\ : CascadeMux
    port map (
            O => \N__35384\,
            I => \N__35381\
        );

    \I__7201\ : InMux
    port map (
            O => \N__35381\,
            I => \N__35378\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__35378\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__7199\ : InMux
    port map (
            O => \N__35375\,
            I => \N__35372\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__35372\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__7197\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35366\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__35366\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__7195\ : CascadeMux
    port map (
            O => \N__35363\,
            I => \N__35360\
        );

    \I__7194\ : InMux
    port map (
            O => \N__35360\,
            I => \N__35357\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__35357\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__7192\ : CascadeMux
    port map (
            O => \N__35354\,
            I => \N__35351\
        );

    \I__7191\ : InMux
    port map (
            O => \N__35351\,
            I => \N__35348\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__35348\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__7189\ : CascadeMux
    port map (
            O => \N__35345\,
            I => \N__35342\
        );

    \I__7188\ : InMux
    port map (
            O => \N__35342\,
            I => \N__35339\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__35339\,
            I => \N__35336\
        );

    \I__7186\ : Odrv4
    port map (
            O => \N__35336\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__7185\ : CascadeMux
    port map (
            O => \N__35333\,
            I => \N__35330\
        );

    \I__7184\ : InMux
    port map (
            O => \N__35330\,
            I => \N__35327\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__35327\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__7182\ : CascadeMux
    port map (
            O => \N__35324\,
            I => \N__35316\
        );

    \I__7181\ : CascadeMux
    port map (
            O => \N__35323\,
            I => \N__35312\
        );

    \I__7180\ : CascadeMux
    port map (
            O => \N__35322\,
            I => \N__35308\
        );

    \I__7179\ : InMux
    port map (
            O => \N__35321\,
            I => \N__35303\
        );

    \I__7178\ : InMux
    port map (
            O => \N__35320\,
            I => \N__35303\
        );

    \I__7177\ : InMux
    port map (
            O => \N__35319\,
            I => \N__35290\
        );

    \I__7176\ : InMux
    port map (
            O => \N__35316\,
            I => \N__35290\
        );

    \I__7175\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35290\
        );

    \I__7174\ : InMux
    port map (
            O => \N__35312\,
            I => \N__35290\
        );

    \I__7173\ : InMux
    port map (
            O => \N__35311\,
            I => \N__35290\
        );

    \I__7172\ : InMux
    port map (
            O => \N__35308\,
            I => \N__35290\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__35303\,
            I => \N__35287\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__35290\,
            I => \N__35284\
        );

    \I__7169\ : Span12Mux_h
    port map (
            O => \N__35287\,
            I => \N__35279\
        );

    \I__7168\ : Span12Mux_s7_v
    port map (
            O => \N__35284\,
            I => \N__35279\
        );

    \I__7167\ : Span12Mux_h
    port map (
            O => \N__35279\,
            I => \N__35276\
        );

    \I__7166\ : Odrv12
    port map (
            O => \N__35276\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__7165\ : CascadeMux
    port map (
            O => \N__35273\,
            I => \N__35270\
        );

    \I__7164\ : InMux
    port map (
            O => \N__35270\,
            I => \N__35267\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__35267\,
            I => \N__35264\
        );

    \I__7162\ : Span4Mux_s2_v
    port map (
            O => \N__35264\,
            I => \N__35261\
        );

    \I__7161\ : Span4Mux_v
    port map (
            O => \N__35261\,
            I => \N__35258\
        );

    \I__7160\ : Odrv4
    port map (
            O => \N__35258\,
            I => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\
        );

    \I__7159\ : InMux
    port map (
            O => \N__35255\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_14\
        );

    \I__7158\ : InMux
    port map (
            O => \N__35252\,
            I => \N__35249\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__35249\,
            I => \N__35246\
        );

    \I__7156\ : Span4Mux_v
    port map (
            O => \N__35246\,
            I => \N__35243\
        );

    \I__7155\ : Odrv4
    port map (
            O => \N__35243\,
            I => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35240\,
            I => \bfn_13_30_0_\
        );

    \I__7153\ : CascadeMux
    port map (
            O => \N__35237\,
            I => \N__35233\
        );

    \I__7152\ : InMux
    port map (
            O => \N__35236\,
            I => \N__35230\
        );

    \I__7151\ : InMux
    port map (
            O => \N__35233\,
            I => \N__35227\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__35230\,
            I => \N__35224\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__35227\,
            I => \N__35219\
        );

    \I__7148\ : Span4Mux_h
    port map (
            O => \N__35224\,
            I => \N__35219\
        );

    \I__7147\ : Span4Mux_v
    port map (
            O => \N__35219\,
            I => \N__35213\
        );

    \I__7146\ : InMux
    port map (
            O => \N__35218\,
            I => \N__35206\
        );

    \I__7145\ : InMux
    port map (
            O => \N__35217\,
            I => \N__35206\
        );

    \I__7144\ : InMux
    port map (
            O => \N__35216\,
            I => \N__35206\
        );

    \I__7143\ : Odrv4
    port map (
            O => \N__35213\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__35206\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__7141\ : InMux
    port map (
            O => \N__35201\,
            I => \N__35198\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__35198\,
            I => \N__35195\
        );

    \I__7139\ : Span4Mux_h
    port map (
            O => \N__35195\,
            I => \N__35192\
        );

    \I__7138\ : Span4Mux_v
    port map (
            O => \N__35192\,
            I => \N__35186\
        );

    \I__7137\ : InMux
    port map (
            O => \N__35191\,
            I => \N__35179\
        );

    \I__7136\ : InMux
    port map (
            O => \N__35190\,
            I => \N__35179\
        );

    \I__7135\ : InMux
    port map (
            O => \N__35189\,
            I => \N__35179\
        );

    \I__7134\ : Odrv4
    port map (
            O => \N__35186\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__35179\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__7132\ : InMux
    port map (
            O => \N__35174\,
            I => \N__35169\
        );

    \I__7131\ : InMux
    port map (
            O => \N__35173\,
            I => \N__35166\
        );

    \I__7130\ : CascadeMux
    port map (
            O => \N__35172\,
            I => \N__35163\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__35169\,
            I => \N__35158\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__35166\,
            I => \N__35158\
        );

    \I__7127\ : InMux
    port map (
            O => \N__35163\,
            I => \N__35153\
        );

    \I__7126\ : Span4Mux_h
    port map (
            O => \N__35158\,
            I => \N__35150\
        );

    \I__7125\ : InMux
    port map (
            O => \N__35157\,
            I => \N__35145\
        );

    \I__7124\ : InMux
    port map (
            O => \N__35156\,
            I => \N__35145\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__35153\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__7122\ : Odrv4
    port map (
            O => \N__35150\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__35145\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__7120\ : InMux
    port map (
            O => \N__35138\,
            I => \N__35135\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__35135\,
            I => \N__35132\
        );

    \I__7118\ : Span4Mux_h
    port map (
            O => \N__35132\,
            I => \N__35128\
        );

    \I__7117\ : InMux
    port map (
            O => \N__35131\,
            I => \N__35125\
        );

    \I__7116\ : Odrv4
    port map (
            O => \N__35128\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__35125\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__7114\ : InMux
    port map (
            O => \N__35120\,
            I => \N__35117\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__35117\,
            I => \N__35113\
        );

    \I__7112\ : InMux
    port map (
            O => \N__35116\,
            I => \N__35110\
        );

    \I__7111\ : Span4Mux_v
    port map (
            O => \N__35113\,
            I => \N__35107\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__35110\,
            I => \N__35104\
        );

    \I__7109\ : Span4Mux_v
    port map (
            O => \N__35107\,
            I => \N__35101\
        );

    \I__7108\ : Span4Mux_h
    port map (
            O => \N__35104\,
            I => \N__35098\
        );

    \I__7107\ : Odrv4
    port map (
            O => \N__35101\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__35098\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__7105\ : CascadeMux
    port map (
            O => \N__35093\,
            I => \N__35089\
        );

    \I__7104\ : InMux
    port map (
            O => \N__35092\,
            I => \N__35086\
        );

    \I__7103\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35083\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__35086\,
            I => \N__35080\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__35083\,
            I => \N__35077\
        );

    \I__7100\ : Span12Mux_h
    port map (
            O => \N__35080\,
            I => \N__35071\
        );

    \I__7099\ : Span4Mux_v
    port map (
            O => \N__35077\,
            I => \N__35068\
        );

    \I__7098\ : InMux
    port map (
            O => \N__35076\,
            I => \N__35063\
        );

    \I__7097\ : InMux
    port map (
            O => \N__35075\,
            I => \N__35063\
        );

    \I__7096\ : InMux
    port map (
            O => \N__35074\,
            I => \N__35060\
        );

    \I__7095\ : Span12Mux_v
    port map (
            O => \N__35071\,
            I => \N__35057\
        );

    \I__7094\ : Span4Mux_v
    port map (
            O => \N__35068\,
            I => \N__35052\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__35063\,
            I => \N__35052\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__35060\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7091\ : Odrv12
    port map (
            O => \N__35057\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7090\ : Odrv4
    port map (
            O => \N__35052\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7089\ : CascadeMux
    port map (
            O => \N__35045\,
            I => \N__35042\
        );

    \I__7088\ : InMux
    port map (
            O => \N__35042\,
            I => \N__35038\
        );

    \I__7087\ : InMux
    port map (
            O => \N__35041\,
            I => \N__35035\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__35038\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__35035\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__7084\ : CascadeMux
    port map (
            O => \N__35030\,
            I => \N__35027\
        );

    \I__7083\ : InMux
    port map (
            O => \N__35027\,
            I => \N__35024\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__35024\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__7081\ : InMux
    port map (
            O => \N__35021\,
            I => \N__35018\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__35018\,
            I => \N__35015\
        );

    \I__7079\ : Span4Mux_v
    port map (
            O => \N__35015\,
            I => \N__35012\
        );

    \I__7078\ : Odrv4
    port map (
            O => \N__35012\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__7077\ : CascadeMux
    port map (
            O => \N__35009\,
            I => \N__35006\
        );

    \I__7076\ : InMux
    port map (
            O => \N__35006\,
            I => \N__35003\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__35003\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__7074\ : InMux
    port map (
            O => \N__35000\,
            I => \N__34997\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__34997\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__7072\ : InMux
    port map (
            O => \N__34994\,
            I => \N__34991\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__34991\,
            I => \N__34988\
        );

    \I__7070\ : Span4Mux_v
    port map (
            O => \N__34988\,
            I => \N__34985\
        );

    \I__7069\ : Sp12to4
    port map (
            O => \N__34985\,
            I => \N__34982\
        );

    \I__7068\ : Span12Mux_h
    port map (
            O => \N__34982\,
            I => \N__34979\
        );

    \I__7067\ : Odrv12
    port map (
            O => \N__34979\,
            I => \pwm_generator_inst.un2_threshold_2_7\
        );

    \I__7066\ : CascadeMux
    port map (
            O => \N__34976\,
            I => \N__34973\
        );

    \I__7065\ : InMux
    port map (
            O => \N__34973\,
            I => \N__34970\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__34970\,
            I => \N__34967\
        );

    \I__7063\ : Span4Mux_v
    port map (
            O => \N__34967\,
            I => \N__34964\
        );

    \I__7062\ : Sp12to4
    port map (
            O => \N__34964\,
            I => \N__34961\
        );

    \I__7061\ : Odrv12
    port map (
            O => \N__34961\,
            I => \pwm_generator_inst.un2_threshold_1_22\
        );

    \I__7060\ : InMux
    port map (
            O => \N__34958\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6\
        );

    \I__7059\ : InMux
    port map (
            O => \N__34955\,
            I => \N__34952\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__34952\,
            I => \N__34949\
        );

    \I__7057\ : Span4Mux_v
    port map (
            O => \N__34949\,
            I => \N__34946\
        );

    \I__7056\ : Span4Mux_h
    port map (
            O => \N__34946\,
            I => \N__34943\
        );

    \I__7055\ : Span4Mux_h
    port map (
            O => \N__34943\,
            I => \N__34940\
        );

    \I__7054\ : Span4Mux_h
    port map (
            O => \N__34940\,
            I => \N__34937\
        );

    \I__7053\ : Odrv4
    port map (
            O => \N__34937\,
            I => \pwm_generator_inst.un2_threshold_2_8\
        );

    \I__7052\ : CascadeMux
    port map (
            O => \N__34934\,
            I => \N__34931\
        );

    \I__7051\ : InMux
    port map (
            O => \N__34931\,
            I => \N__34928\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__34928\,
            I => \N__34925\
        );

    \I__7049\ : Span12Mux_s10_v
    port map (
            O => \N__34925\,
            I => \N__34922\
        );

    \I__7048\ : Span12Mux_h
    port map (
            O => \N__34922\,
            I => \N__34919\
        );

    \I__7047\ : Odrv12
    port map (
            O => \N__34919\,
            I => \pwm_generator_inst.un2_threshold_1_23\
        );

    \I__7046\ : InMux
    port map (
            O => \N__34916\,
            I => \bfn_13_29_0_\
        );

    \I__7045\ : InMux
    port map (
            O => \N__34913\,
            I => \N__34910\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__34910\,
            I => \N__34907\
        );

    \I__7043\ : Span4Mux_v
    port map (
            O => \N__34907\,
            I => \N__34904\
        );

    \I__7042\ : Span4Mux_h
    port map (
            O => \N__34904\,
            I => \N__34901\
        );

    \I__7041\ : Span4Mux_h
    port map (
            O => \N__34901\,
            I => \N__34898\
        );

    \I__7040\ : Span4Mux_h
    port map (
            O => \N__34898\,
            I => \N__34895\
        );

    \I__7039\ : Odrv4
    port map (
            O => \N__34895\,
            I => \pwm_generator_inst.un2_threshold_2_9\
        );

    \I__7038\ : CascadeMux
    port map (
            O => \N__34892\,
            I => \N__34889\
        );

    \I__7037\ : InMux
    port map (
            O => \N__34889\,
            I => \N__34886\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__34886\,
            I => \N__34883\
        );

    \I__7035\ : Span12Mux_s8_v
    port map (
            O => \N__34883\,
            I => \N__34880\
        );

    \I__7034\ : Span12Mux_h
    port map (
            O => \N__34880\,
            I => \N__34877\
        );

    \I__7033\ : Odrv12
    port map (
            O => \N__34877\,
            I => \pwm_generator_inst.un2_threshold_1_24\
        );

    \I__7032\ : InMux
    port map (
            O => \N__34874\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8\
        );

    \I__7031\ : InMux
    port map (
            O => \N__34871\,
            I => \N__34868\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__34868\,
            I => \N__34865\
        );

    \I__7029\ : Span4Mux_v
    port map (
            O => \N__34865\,
            I => \N__34862\
        );

    \I__7028\ : Sp12to4
    port map (
            O => \N__34862\,
            I => \N__34859\
        );

    \I__7027\ : Span12Mux_h
    port map (
            O => \N__34859\,
            I => \N__34856\
        );

    \I__7026\ : Odrv12
    port map (
            O => \N__34856\,
            I => \pwm_generator_inst.un2_threshold_2_10\
        );

    \I__7025\ : InMux
    port map (
            O => \N__34853\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9\
        );

    \I__7024\ : CascadeMux
    port map (
            O => \N__34850\,
            I => \N__34847\
        );

    \I__7023\ : InMux
    port map (
            O => \N__34847\,
            I => \N__34844\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__34844\,
            I => \N__34841\
        );

    \I__7021\ : Span4Mux_s3_v
    port map (
            O => \N__34841\,
            I => \N__34838\
        );

    \I__7020\ : Sp12to4
    port map (
            O => \N__34838\,
            I => \N__34835\
        );

    \I__7019\ : Span12Mux_h
    port map (
            O => \N__34835\,
            I => \N__34832\
        );

    \I__7018\ : Odrv12
    port map (
            O => \N__34832\,
            I => \pwm_generator_inst.un2_threshold_2_11\
        );

    \I__7017\ : InMux
    port map (
            O => \N__34829\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10\
        );

    \I__7016\ : InMux
    port map (
            O => \N__34826\,
            I => \N__34823\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__34823\,
            I => \N__34820\
        );

    \I__7014\ : Span4Mux_s2_v
    port map (
            O => \N__34820\,
            I => \N__34817\
        );

    \I__7013\ : Span4Mux_v
    port map (
            O => \N__34817\,
            I => \N__34814\
        );

    \I__7012\ : Sp12to4
    port map (
            O => \N__34814\,
            I => \N__34811\
        );

    \I__7011\ : Odrv12
    port map (
            O => \N__34811\,
            I => \pwm_generator_inst.un2_threshold_2_12\
        );

    \I__7010\ : InMux
    port map (
            O => \N__34808\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11\
        );

    \I__7009\ : CascadeMux
    port map (
            O => \N__34805\,
            I => \N__34802\
        );

    \I__7008\ : InMux
    port map (
            O => \N__34802\,
            I => \N__34799\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__34799\,
            I => \N__34796\
        );

    \I__7006\ : Sp12to4
    port map (
            O => \N__34796\,
            I => \N__34793\
        );

    \I__7005\ : Span12Mux_h
    port map (
            O => \N__34793\,
            I => \N__34790\
        );

    \I__7004\ : Odrv12
    port map (
            O => \N__34790\,
            I => \pwm_generator_inst.un2_threshold_2_13\
        );

    \I__7003\ : InMux
    port map (
            O => \N__34787\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_12\
        );

    \I__7002\ : InMux
    port map (
            O => \N__34784\,
            I => \N__34781\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__34781\,
            I => \N__34778\
        );

    \I__7000\ : Span4Mux_v
    port map (
            O => \N__34778\,
            I => \N__34775\
        );

    \I__6999\ : Sp12to4
    port map (
            O => \N__34775\,
            I => \N__34772\
        );

    \I__6998\ : Span12Mux_h
    port map (
            O => \N__34772\,
            I => \N__34769\
        );

    \I__6997\ : Odrv12
    port map (
            O => \N__34769\,
            I => \pwm_generator_inst.un2_threshold_2_14\
        );

    \I__6996\ : InMux
    port map (
            O => \N__34766\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_13\
        );

    \I__6995\ : InMux
    port map (
            O => \N__34763\,
            I => \N__34760\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__34760\,
            I => \N__34757\
        );

    \I__6993\ : Odrv12
    port map (
            O => \N__34757\,
            I => \pwm_generator_inst.un19_threshold_axb_7\
        );

    \I__6992\ : InMux
    port map (
            O => \N__34754\,
            I => \N__34751\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__34751\,
            I => \N__34748\
        );

    \I__6990\ : Span4Mux_v
    port map (
            O => \N__34748\,
            I => \N__34745\
        );

    \I__6989\ : Span4Mux_h
    port map (
            O => \N__34745\,
            I => \N__34742\
        );

    \I__6988\ : Span4Mux_h
    port map (
            O => \N__34742\,
            I => \N__34739\
        );

    \I__6987\ : Span4Mux_h
    port map (
            O => \N__34739\,
            I => \N__34736\
        );

    \I__6986\ : Odrv4
    port map (
            O => \N__34736\,
            I => \pwm_generator_inst.un2_threshold_2_0\
        );

    \I__6985\ : CascadeMux
    port map (
            O => \N__34733\,
            I => \N__34730\
        );

    \I__6984\ : InMux
    port map (
            O => \N__34730\,
            I => \N__34727\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__34727\,
            I => \N__34724\
        );

    \I__6982\ : Span12Mux_s11_v
    port map (
            O => \N__34724\,
            I => \N__34721\
        );

    \I__6981\ : Span12Mux_h
    port map (
            O => \N__34721\,
            I => \N__34718\
        );

    \I__6980\ : Odrv12
    port map (
            O => \N__34718\,
            I => \pwm_generator_inst.un2_threshold_1_15\
        );

    \I__6979\ : InMux
    port map (
            O => \N__34715\,
            I => \N__34712\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__34712\,
            I => \N__34709\
        );

    \I__6977\ : Span4Mux_v
    port map (
            O => \N__34709\,
            I => \N__34706\
        );

    \I__6976\ : Sp12to4
    port map (
            O => \N__34706\,
            I => \N__34703\
        );

    \I__6975\ : Span12Mux_h
    port map (
            O => \N__34703\,
            I => \N__34700\
        );

    \I__6974\ : Odrv12
    port map (
            O => \N__34700\,
            I => \pwm_generator_inst.un2_threshold_2_1\
        );

    \I__6973\ : CascadeMux
    port map (
            O => \N__34697\,
            I => \N__34694\
        );

    \I__6972\ : InMux
    port map (
            O => \N__34694\,
            I => \N__34691\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__34691\,
            I => \N__34688\
        );

    \I__6970\ : Span12Mux_s9_v
    port map (
            O => \N__34688\,
            I => \N__34685\
        );

    \I__6969\ : Span12Mux_h
    port map (
            O => \N__34685\,
            I => \N__34682\
        );

    \I__6968\ : Odrv12
    port map (
            O => \N__34682\,
            I => \pwm_generator_inst.un2_threshold_1_16\
        );

    \I__6967\ : InMux
    port map (
            O => \N__34679\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0\
        );

    \I__6966\ : InMux
    port map (
            O => \N__34676\,
            I => \N__34673\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__34673\,
            I => \N__34670\
        );

    \I__6964\ : Span4Mux_v
    port map (
            O => \N__34670\,
            I => \N__34667\
        );

    \I__6963\ : Span4Mux_h
    port map (
            O => \N__34667\,
            I => \N__34664\
        );

    \I__6962\ : Span4Mux_h
    port map (
            O => \N__34664\,
            I => \N__34661\
        );

    \I__6961\ : Span4Mux_h
    port map (
            O => \N__34661\,
            I => \N__34658\
        );

    \I__6960\ : Odrv4
    port map (
            O => \N__34658\,
            I => \pwm_generator_inst.un2_threshold_2_2\
        );

    \I__6959\ : CascadeMux
    port map (
            O => \N__34655\,
            I => \N__34652\
        );

    \I__6958\ : InMux
    port map (
            O => \N__34652\,
            I => \N__34649\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__34649\,
            I => \N__34646\
        );

    \I__6956\ : Span12Mux_s4_v
    port map (
            O => \N__34646\,
            I => \N__34643\
        );

    \I__6955\ : Span12Mux_h
    port map (
            O => \N__34643\,
            I => \N__34640\
        );

    \I__6954\ : Odrv12
    port map (
            O => \N__34640\,
            I => \pwm_generator_inst.un2_threshold_1_17\
        );

    \I__6953\ : InMux
    port map (
            O => \N__34637\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1\
        );

    \I__6952\ : InMux
    port map (
            O => \N__34634\,
            I => \N__34631\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__34631\,
            I => \N__34628\
        );

    \I__6950\ : Span4Mux_v
    port map (
            O => \N__34628\,
            I => \N__34625\
        );

    \I__6949\ : Sp12to4
    port map (
            O => \N__34625\,
            I => \N__34622\
        );

    \I__6948\ : Span12Mux_h
    port map (
            O => \N__34622\,
            I => \N__34619\
        );

    \I__6947\ : Odrv12
    port map (
            O => \N__34619\,
            I => \pwm_generator_inst.un2_threshold_2_3\
        );

    \I__6946\ : CascadeMux
    port map (
            O => \N__34616\,
            I => \N__34613\
        );

    \I__6945\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34610\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__34610\,
            I => \N__34607\
        );

    \I__6943\ : Span4Mux_h
    port map (
            O => \N__34607\,
            I => \N__34604\
        );

    \I__6942\ : Span4Mux_h
    port map (
            O => \N__34604\,
            I => \N__34601\
        );

    \I__6941\ : Span4Mux_h
    port map (
            O => \N__34601\,
            I => \N__34598\
        );

    \I__6940\ : Odrv4
    port map (
            O => \N__34598\,
            I => \pwm_generator_inst.un2_threshold_1_18\
        );

    \I__6939\ : InMux
    port map (
            O => \N__34595\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2\
        );

    \I__6938\ : InMux
    port map (
            O => \N__34592\,
            I => \N__34589\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__34589\,
            I => \N__34586\
        );

    \I__6936\ : Span4Mux_s3_v
    port map (
            O => \N__34586\,
            I => \N__34583\
        );

    \I__6935\ : Span4Mux_v
    port map (
            O => \N__34583\,
            I => \N__34580\
        );

    \I__6934\ : Sp12to4
    port map (
            O => \N__34580\,
            I => \N__34577\
        );

    \I__6933\ : Odrv12
    port map (
            O => \N__34577\,
            I => \pwm_generator_inst.un2_threshold_2_4\
        );

    \I__6932\ : CascadeMux
    port map (
            O => \N__34574\,
            I => \N__34571\
        );

    \I__6931\ : InMux
    port map (
            O => \N__34571\,
            I => \N__34568\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__34568\,
            I => \N__34565\
        );

    \I__6929\ : Span12Mux_h
    port map (
            O => \N__34565\,
            I => \N__34562\
        );

    \I__6928\ : Odrv12
    port map (
            O => \N__34562\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__6927\ : InMux
    port map (
            O => \N__34559\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3\
        );

    \I__6926\ : InMux
    port map (
            O => \N__34556\,
            I => \N__34553\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__34553\,
            I => \N__34550\
        );

    \I__6924\ : Span12Mux_h
    port map (
            O => \N__34550\,
            I => \N__34547\
        );

    \I__6923\ : Span12Mux_h
    port map (
            O => \N__34547\,
            I => \N__34544\
        );

    \I__6922\ : Odrv12
    port map (
            O => \N__34544\,
            I => \pwm_generator_inst.un2_threshold_2_5\
        );

    \I__6921\ : CascadeMux
    port map (
            O => \N__34541\,
            I => \N__34538\
        );

    \I__6920\ : InMux
    port map (
            O => \N__34538\,
            I => \N__34535\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__34535\,
            I => \N__34532\
        );

    \I__6918\ : Span4Mux_h
    port map (
            O => \N__34532\,
            I => \N__34529\
        );

    \I__6917\ : Span4Mux_h
    port map (
            O => \N__34529\,
            I => \N__34526\
        );

    \I__6916\ : Span4Mux_h
    port map (
            O => \N__34526\,
            I => \N__34523\
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__34523\,
            I => \pwm_generator_inst.un2_threshold_1_20\
        );

    \I__6914\ : InMux
    port map (
            O => \N__34520\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4\
        );

    \I__6913\ : InMux
    port map (
            O => \N__34517\,
            I => \N__34514\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__34514\,
            I => \N__34511\
        );

    \I__6911\ : Span4Mux_v
    port map (
            O => \N__34511\,
            I => \N__34508\
        );

    \I__6910\ : Sp12to4
    port map (
            O => \N__34508\,
            I => \N__34505\
        );

    \I__6909\ : Span12Mux_h
    port map (
            O => \N__34505\,
            I => \N__34502\
        );

    \I__6908\ : Odrv12
    port map (
            O => \N__34502\,
            I => \pwm_generator_inst.un2_threshold_2_6\
        );

    \I__6907\ : CascadeMux
    port map (
            O => \N__34499\,
            I => \N__34496\
        );

    \I__6906\ : InMux
    port map (
            O => \N__34496\,
            I => \N__34493\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__34493\,
            I => \N__34490\
        );

    \I__6904\ : Span4Mux_h
    port map (
            O => \N__34490\,
            I => \N__34487\
        );

    \I__6903\ : Span4Mux_h
    port map (
            O => \N__34487\,
            I => \N__34484\
        );

    \I__6902\ : Span4Mux_h
    port map (
            O => \N__34484\,
            I => \N__34481\
        );

    \I__6901\ : Odrv4
    port map (
            O => \N__34481\,
            I => \pwm_generator_inst.un2_threshold_1_21\
        );

    \I__6900\ : InMux
    port map (
            O => \N__34478\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5\
        );

    \I__6899\ : InMux
    port map (
            O => \N__34475\,
            I => \pwm_generator_inst.un19_threshold_cry_8\
        );

    \I__6898\ : InMux
    port map (
            O => \N__34472\,
            I => \N__34469\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__34469\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\
        );

    \I__6896\ : InMux
    port map (
            O => \N__34466\,
            I => \N__34463\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__34463\,
            I => \pwm_generator_inst.un19_threshold_axb_5\
        );

    \I__6894\ : InMux
    port map (
            O => \N__34460\,
            I => \N__34457\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__34457\,
            I => \pwm_generator_inst.un19_threshold_axb_3\
        );

    \I__6892\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34451\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__34451\,
            I => \pwm_generator_inst.un19_threshold_axb_6\
        );

    \I__6890\ : InMux
    port map (
            O => \N__34448\,
            I => \N__34445\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__34445\,
            I => \pwm_generator_inst.un19_threshold_axb_4\
        );

    \I__6888\ : InMux
    port map (
            O => \N__34442\,
            I => \N__34439\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__34439\,
            I => \pwm_generator_inst.un19_threshold_axb_0\
        );

    \I__6886\ : InMux
    port map (
            O => \N__34436\,
            I => \N__34433\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__34433\,
            I => \pwm_generator_inst.un19_threshold_axb_8\
        );

    \I__6884\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34427\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__34427\,
            I => \N__34424\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__34424\,
            I => \pwm_generator_inst.un19_threshold_axb_2\
        );

    \I__6881\ : CascadeMux
    port map (
            O => \N__34421\,
            I => \N__34418\
        );

    \I__6880\ : InMux
    port map (
            O => \N__34418\,
            I => \N__34415\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__34415\,
            I => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\
        );

    \I__6878\ : InMux
    port map (
            O => \N__34412\,
            I => \pwm_generator_inst.un19_threshold_cry_0\
        );

    \I__6877\ : CascadeMux
    port map (
            O => \N__34409\,
            I => \N__34406\
        );

    \I__6876\ : InMux
    port map (
            O => \N__34406\,
            I => \N__34403\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__34403\,
            I => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\
        );

    \I__6874\ : InMux
    port map (
            O => \N__34400\,
            I => \pwm_generator_inst.un19_threshold_cry_1\
        );

    \I__6873\ : InMux
    port map (
            O => \N__34397\,
            I => \N__34394\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__34394\,
            I => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\
        );

    \I__6871\ : InMux
    port map (
            O => \N__34391\,
            I => \pwm_generator_inst.un19_threshold_cry_2\
        );

    \I__6870\ : InMux
    port map (
            O => \N__34388\,
            I => \N__34385\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__34385\,
            I => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\
        );

    \I__6868\ : InMux
    port map (
            O => \N__34382\,
            I => \pwm_generator_inst.un19_threshold_cry_3\
        );

    \I__6867\ : CascadeMux
    port map (
            O => \N__34379\,
            I => \N__34376\
        );

    \I__6866\ : InMux
    port map (
            O => \N__34376\,
            I => \N__34373\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__34373\,
            I => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\
        );

    \I__6864\ : InMux
    port map (
            O => \N__34370\,
            I => \pwm_generator_inst.un19_threshold_cry_4\
        );

    \I__6863\ : InMux
    port map (
            O => \N__34367\,
            I => \N__34364\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__34364\,
            I => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\
        );

    \I__6861\ : InMux
    port map (
            O => \N__34361\,
            I => \pwm_generator_inst.un19_threshold_cry_5\
        );

    \I__6860\ : InMux
    port map (
            O => \N__34358\,
            I => \N__34355\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__34355\,
            I => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\
        );

    \I__6858\ : InMux
    port map (
            O => \N__34352\,
            I => \pwm_generator_inst.un19_threshold_cry_6\
        );

    \I__6857\ : CascadeMux
    port map (
            O => \N__34349\,
            I => \N__34346\
        );

    \I__6856\ : InMux
    port map (
            O => \N__34346\,
            I => \N__34343\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__34343\,
            I => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\
        );

    \I__6854\ : InMux
    port map (
            O => \N__34340\,
            I => \bfn_13_25_0_\
        );

    \I__6853\ : InMux
    port map (
            O => \N__34337\,
            I => \N__34334\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__34334\,
            I => \N__34329\
        );

    \I__6851\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34326\
        );

    \I__6850\ : InMux
    port map (
            O => \N__34332\,
            I => \N__34323\
        );

    \I__6849\ : Span4Mux_v
    port map (
            O => \N__34329\,
            I => \N__34320\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__34326\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__34323\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__6846\ : Odrv4
    port map (
            O => \N__34320\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__6845\ : InMux
    port map (
            O => \N__34313\,
            I => \N__34309\
        );

    \I__6844\ : InMux
    port map (
            O => \N__34312\,
            I => \N__34305\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__34309\,
            I => \N__34302\
        );

    \I__6842\ : InMux
    port map (
            O => \N__34308\,
            I => \N__34299\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__34305\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__6840\ : Odrv4
    port map (
            O => \N__34302\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__34299\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__6838\ : InMux
    port map (
            O => \N__34292\,
            I => \N__34287\
        );

    \I__6837\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34284\
        );

    \I__6836\ : InMux
    port map (
            O => \N__34290\,
            I => \N__34281\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__34287\,
            I => \N__34278\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__34284\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__34281\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__6832\ : Odrv4
    port map (
            O => \N__34278\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__6831\ : InMux
    port map (
            O => \N__34271\,
            I => \N__34266\
        );

    \I__6830\ : InMux
    port map (
            O => \N__34270\,
            I => \N__34263\
        );

    \I__6829\ : InMux
    port map (
            O => \N__34269\,
            I => \N__34260\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__34266\,
            I => \N__34257\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__34263\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__34260\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__6825\ : Odrv4
    port map (
            O => \N__34257\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__6824\ : CascadeMux
    port map (
            O => \N__34250\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__6823\ : InMux
    port map (
            O => \N__34247\,
            I => \N__34242\
        );

    \I__6822\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34239\
        );

    \I__6821\ : InMux
    port map (
            O => \N__34245\,
            I => \N__34236\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__34242\,
            I => \N__34233\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__34239\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__34236\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__6817\ : Odrv4
    port map (
            O => \N__34233\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__6816\ : InMux
    port map (
            O => \N__34226\,
            I => \N__34210\
        );

    \I__6815\ : InMux
    port map (
            O => \N__34225\,
            I => \N__34210\
        );

    \I__6814\ : InMux
    port map (
            O => \N__34224\,
            I => \N__34210\
        );

    \I__6813\ : InMux
    port map (
            O => \N__34223\,
            I => \N__34210\
        );

    \I__6812\ : InMux
    port map (
            O => \N__34222\,
            I => \N__34195\
        );

    \I__6811\ : InMux
    port map (
            O => \N__34221\,
            I => \N__34195\
        );

    \I__6810\ : InMux
    port map (
            O => \N__34220\,
            I => \N__34195\
        );

    \I__6809\ : InMux
    port map (
            O => \N__34219\,
            I => \N__34195\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__34210\,
            I => \N__34188\
        );

    \I__6807\ : InMux
    port map (
            O => \N__34209\,
            I => \N__34183\
        );

    \I__6806\ : InMux
    port map (
            O => \N__34208\,
            I => \N__34183\
        );

    \I__6805\ : InMux
    port map (
            O => \N__34207\,
            I => \N__34174\
        );

    \I__6804\ : InMux
    port map (
            O => \N__34206\,
            I => \N__34174\
        );

    \I__6803\ : InMux
    port map (
            O => \N__34205\,
            I => \N__34174\
        );

    \I__6802\ : InMux
    port map (
            O => \N__34204\,
            I => \N__34174\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__34195\,
            I => \N__34171\
        );

    \I__6800\ : InMux
    port map (
            O => \N__34194\,
            I => \N__34162\
        );

    \I__6799\ : InMux
    port map (
            O => \N__34193\,
            I => \N__34162\
        );

    \I__6798\ : InMux
    port map (
            O => \N__34192\,
            I => \N__34162\
        );

    \I__6797\ : InMux
    port map (
            O => \N__34191\,
            I => \N__34162\
        );

    \I__6796\ : Span4Mux_v
    port map (
            O => \N__34188\,
            I => \N__34143\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__34183\,
            I => \N__34143\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__34174\,
            I => \N__34143\
        );

    \I__6793\ : Span4Mux_v
    port map (
            O => \N__34171\,
            I => \N__34143\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__34162\,
            I => \N__34143\
        );

    \I__6791\ : InMux
    port map (
            O => \N__34161\,
            I => \N__34134\
        );

    \I__6790\ : InMux
    port map (
            O => \N__34160\,
            I => \N__34134\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34159\,
            I => \N__34134\
        );

    \I__6788\ : InMux
    port map (
            O => \N__34158\,
            I => \N__34134\
        );

    \I__6787\ : InMux
    port map (
            O => \N__34157\,
            I => \N__34125\
        );

    \I__6786\ : InMux
    port map (
            O => \N__34156\,
            I => \N__34125\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34155\,
            I => \N__34125\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34154\,
            I => \N__34125\
        );

    \I__6783\ : Span4Mux_v
    port map (
            O => \N__34143\,
            I => \N__34116\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__34134\,
            I => \N__34116\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__34125\,
            I => \N__34113\
        );

    \I__6780\ : InMux
    port map (
            O => \N__34124\,
            I => \N__34104\
        );

    \I__6779\ : InMux
    port map (
            O => \N__34123\,
            I => \N__34104\
        );

    \I__6778\ : InMux
    port map (
            O => \N__34122\,
            I => \N__34104\
        );

    \I__6777\ : InMux
    port map (
            O => \N__34121\,
            I => \N__34104\
        );

    \I__6776\ : Span4Mux_h
    port map (
            O => \N__34116\,
            I => \N__34099\
        );

    \I__6775\ : Span4Mux_h
    port map (
            O => \N__34113\,
            I => \N__34099\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__34104\,
            I => \N__34096\
        );

    \I__6773\ : Span4Mux_h
    port map (
            O => \N__34099\,
            I => \N__34093\
        );

    \I__6772\ : Odrv12
    port map (
            O => \N__34096\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__6771\ : Odrv4
    port map (
            O => \N__34093\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__6770\ : InMux
    port map (
            O => \N__34088\,
            I => \N__34083\
        );

    \I__6769\ : InMux
    port map (
            O => \N__34087\,
            I => \N__34080\
        );

    \I__6768\ : InMux
    port map (
            O => \N__34086\,
            I => \N__34077\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__34083\,
            I => \N__34074\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__34080\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__34077\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__6764\ : Odrv4
    port map (
            O => \N__34074\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__6763\ : InMux
    port map (
            O => \N__34067\,
            I => \N__34063\
        );

    \I__6762\ : InMux
    port map (
            O => \N__34066\,
            I => \N__34059\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__34063\,
            I => \N__34056\
        );

    \I__6760\ : InMux
    port map (
            O => \N__34062\,
            I => \N__34053\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__34059\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__6758\ : Odrv4
    port map (
            O => \N__34056\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__34053\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__6756\ : InMux
    port map (
            O => \N__34046\,
            I => \N__34041\
        );

    \I__6755\ : InMux
    port map (
            O => \N__34045\,
            I => \N__34038\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34044\,
            I => \N__34035\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__34041\,
            I => \N__34032\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__34038\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__34035\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__6750\ : Odrv4
    port map (
            O => \N__34032\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__6749\ : InMux
    port map (
            O => \N__34025\,
            I => \N__34020\
        );

    \I__6748\ : InMux
    port map (
            O => \N__34024\,
            I => \N__34017\
        );

    \I__6747\ : InMux
    port map (
            O => \N__34023\,
            I => \N__34014\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__34020\,
            I => \N__34011\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__34017\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__34014\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__6743\ : Odrv4
    port map (
            O => \N__34011\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__6742\ : InMux
    port map (
            O => \N__34004\,
            I => \N__33999\
        );

    \I__6741\ : InMux
    port map (
            O => \N__34003\,
            I => \N__33996\
        );

    \I__6740\ : InMux
    port map (
            O => \N__34002\,
            I => \N__33993\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__33999\,
            I => \N__33990\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__33996\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__33993\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__6736\ : Odrv4
    port map (
            O => \N__33990\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__6735\ : CascadeMux
    port map (
            O => \N__33983\,
            I => \pwm_generator_inst.un1_counterlto9_2_cascade_\
        );

    \I__6734\ : InMux
    port map (
            O => \N__33980\,
            I => \N__33977\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__33977\,
            I => \pwm_generator_inst.un1_counterlt9\
        );

    \I__6732\ : InMux
    port map (
            O => \N__33974\,
            I => \N__33956\
        );

    \I__6731\ : InMux
    port map (
            O => \N__33973\,
            I => \N__33956\
        );

    \I__6730\ : InMux
    port map (
            O => \N__33972\,
            I => \N__33956\
        );

    \I__6729\ : InMux
    port map (
            O => \N__33971\,
            I => \N__33956\
        );

    \I__6728\ : InMux
    port map (
            O => \N__33970\,
            I => \N__33951\
        );

    \I__6727\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33951\
        );

    \I__6726\ : InMux
    port map (
            O => \N__33968\,
            I => \N__33942\
        );

    \I__6725\ : InMux
    port map (
            O => \N__33967\,
            I => \N__33942\
        );

    \I__6724\ : InMux
    port map (
            O => \N__33966\,
            I => \N__33942\
        );

    \I__6723\ : InMux
    port map (
            O => \N__33965\,
            I => \N__33942\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__33956\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__33951\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__33942\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__6719\ : InMux
    port map (
            O => \N__33935\,
            I => \N__33932\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__33932\,
            I => \N__33928\
        );

    \I__6717\ : InMux
    port map (
            O => \N__33931\,
            I => \N__33925\
        );

    \I__6716\ : Span4Mux_h
    port map (
            O => \N__33928\,
            I => \N__33922\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__33925\,
            I => \N__33919\
        );

    \I__6714\ : Sp12to4
    port map (
            O => \N__33922\,
            I => \N__33916\
        );

    \I__6713\ : Span4Mux_s3_h
    port map (
            O => \N__33919\,
            I => \N__33913\
        );

    \I__6712\ : Span12Mux_v
    port map (
            O => \N__33916\,
            I => \N__33910\
        );

    \I__6711\ : Span4Mux_h
    port map (
            O => \N__33913\,
            I => \N__33907\
        );

    \I__6710\ : Odrv12
    port map (
            O => \N__33910\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__6709\ : Odrv4
    port map (
            O => \N__33907\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__6708\ : InMux
    port map (
            O => \N__33902\,
            I => \N__33899\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__33899\,
            I => \N__33895\
        );

    \I__6706\ : InMux
    port map (
            O => \N__33898\,
            I => \N__33892\
        );

    \I__6705\ : Span4Mux_v
    port map (
            O => \N__33895\,
            I => \N__33889\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__33892\,
            I => \N__33886\
        );

    \I__6703\ : Sp12to4
    port map (
            O => \N__33889\,
            I => \N__33883\
        );

    \I__6702\ : Span4Mux_s3_h
    port map (
            O => \N__33886\,
            I => \N__33880\
        );

    \I__6701\ : Span12Mux_h
    port map (
            O => \N__33883\,
            I => \N__33877\
        );

    \I__6700\ : Span4Mux_h
    port map (
            O => \N__33880\,
            I => \N__33874\
        );

    \I__6699\ : Odrv12
    port map (
            O => \N__33877\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__6698\ : Odrv4
    port map (
            O => \N__33874\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__6697\ : InMux
    port map (
            O => \N__33869\,
            I => \N__33866\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__33866\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\
        );

    \I__6695\ : CascadeMux
    port map (
            O => \N__33863\,
            I => \N__33860\
        );

    \I__6694\ : InMux
    port map (
            O => \N__33860\,
            I => \N__33856\
        );

    \I__6693\ : CascadeMux
    port map (
            O => \N__33859\,
            I => \N__33853\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__33856\,
            I => \N__33850\
        );

    \I__6691\ : InMux
    port map (
            O => \N__33853\,
            I => \N__33845\
        );

    \I__6690\ : Span4Mux_v
    port map (
            O => \N__33850\,
            I => \N__33842\
        );

    \I__6689\ : InMux
    port map (
            O => \N__33849\,
            I => \N__33839\
        );

    \I__6688\ : InMux
    port map (
            O => \N__33848\,
            I => \N__33836\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__33845\,
            I => \N__33833\
        );

    \I__6686\ : Span4Mux_h
    port map (
            O => \N__33842\,
            I => \N__33826\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__33839\,
            I => \N__33826\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__33836\,
            I => \N__33826\
        );

    \I__6683\ : Span4Mux_v
    port map (
            O => \N__33833\,
            I => \N__33823\
        );

    \I__6682\ : Span4Mux_v
    port map (
            O => \N__33826\,
            I => \N__33820\
        );

    \I__6681\ : Odrv4
    port map (
            O => \N__33823\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__6680\ : Odrv4
    port map (
            O => \N__33820\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__6679\ : InMux
    port map (
            O => \N__33815\,
            I => \N__33812\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__33812\,
            I => \N__33807\
        );

    \I__6677\ : CascadeMux
    port map (
            O => \N__33811\,
            I => \N__33804\
        );

    \I__6676\ : InMux
    port map (
            O => \N__33810\,
            I => \N__33801\
        );

    \I__6675\ : Span4Mux_h
    port map (
            O => \N__33807\,
            I => \N__33798\
        );

    \I__6674\ : InMux
    port map (
            O => \N__33804\,
            I => \N__33795\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__33801\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__6672\ : Odrv4
    port map (
            O => \N__33798\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__33795\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__6670\ : InMux
    port map (
            O => \N__33788\,
            I => \N__33785\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__33785\,
            I => \N__33782\
        );

    \I__6668\ : Odrv4
    port map (
            O => \N__33782\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__6667\ : InMux
    port map (
            O => \N__33779\,
            I => \N__33776\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__33776\,
            I => \N__33773\
        );

    \I__6665\ : Span4Mux_h
    port map (
            O => \N__33773\,
            I => \N__33768\
        );

    \I__6664\ : InMux
    port map (
            O => \N__33772\,
            I => \N__33765\
        );

    \I__6663\ : InMux
    port map (
            O => \N__33771\,
            I => \N__33762\
        );

    \I__6662\ : Span4Mux_v
    port map (
            O => \N__33768\,
            I => \N__33759\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__33765\,
            I => \N__33754\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__33762\,
            I => \N__33754\
        );

    \I__6659\ : Span4Mux_h
    port map (
            O => \N__33759\,
            I => \N__33751\
        );

    \I__6658\ : Span4Mux_v
    port map (
            O => \N__33754\,
            I => \N__33748\
        );

    \I__6657\ : Odrv4
    port map (
            O => \N__33751\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__6656\ : Odrv4
    port map (
            O => \N__33748\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__6655\ : CEMux
    port map (
            O => \N__33743\,
            I => \N__33719\
        );

    \I__6654\ : CEMux
    port map (
            O => \N__33742\,
            I => \N__33719\
        );

    \I__6653\ : CEMux
    port map (
            O => \N__33741\,
            I => \N__33719\
        );

    \I__6652\ : CEMux
    port map (
            O => \N__33740\,
            I => \N__33719\
        );

    \I__6651\ : CEMux
    port map (
            O => \N__33739\,
            I => \N__33719\
        );

    \I__6650\ : CEMux
    port map (
            O => \N__33738\,
            I => \N__33719\
        );

    \I__6649\ : CEMux
    port map (
            O => \N__33737\,
            I => \N__33719\
        );

    \I__6648\ : CEMux
    port map (
            O => \N__33736\,
            I => \N__33719\
        );

    \I__6647\ : GlobalMux
    port map (
            O => \N__33719\,
            I => \N__33716\
        );

    \I__6646\ : gio2CtrlBuf
    port map (
            O => \N__33716\,
            I => \current_shift_inst.timer_s1.N_162_i_g\
        );

    \I__6645\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33709\
        );

    \I__6644\ : CascadeMux
    port map (
            O => \N__33712\,
            I => \N__33705\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__33709\,
            I => \N__33702\
        );

    \I__6642\ : InMux
    port map (
            O => \N__33708\,
            I => \N__33699\
        );

    \I__6641\ : InMux
    port map (
            O => \N__33705\,
            I => \N__33696\
        );

    \I__6640\ : Span4Mux_h
    port map (
            O => \N__33702\,
            I => \N__33688\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__33699\,
            I => \N__33688\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__33696\,
            I => \N__33688\
        );

    \I__6637\ : InMux
    port map (
            O => \N__33695\,
            I => \N__33685\
        );

    \I__6636\ : Span4Mux_h
    port map (
            O => \N__33688\,
            I => \N__33682\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__33685\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__6634\ : Odrv4
    port map (
            O => \N__33682\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__6633\ : InMux
    port map (
            O => \N__33677\,
            I => \N__33674\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__33674\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__6631\ : CascadeMux
    port map (
            O => \N__33671\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__6630\ : InMux
    port map (
            O => \N__33668\,
            I => \N__33664\
        );

    \I__6629\ : InMux
    port map (
            O => \N__33667\,
            I => \N__33661\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__33664\,
            I => \N__33658\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__33661\,
            I => \N__33655\
        );

    \I__6626\ : Span4Mux_v
    port map (
            O => \N__33658\,
            I => \N__33650\
        );

    \I__6625\ : Span4Mux_v
    port map (
            O => \N__33655\,
            I => \N__33650\
        );

    \I__6624\ : Span4Mux_h
    port map (
            O => \N__33650\,
            I => \N__33645\
        );

    \I__6623\ : InMux
    port map (
            O => \N__33649\,
            I => \N__33642\
        );

    \I__6622\ : InMux
    port map (
            O => \N__33648\,
            I => \N__33639\
        );

    \I__6621\ : Odrv4
    port map (
            O => \N__33645\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__33642\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__33639\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6618\ : CascadeMux
    port map (
            O => \N__33632\,
            I => \N__33629\
        );

    \I__6617\ : InMux
    port map (
            O => \N__33629\,
            I => \N__33626\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__33626\,
            I => \N__33623\
        );

    \I__6615\ : Span4Mux_v
    port map (
            O => \N__33623\,
            I => \N__33620\
        );

    \I__6614\ : Odrv4
    port map (
            O => \N__33620\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__6613\ : CascadeMux
    port map (
            O => \N__33617\,
            I => \N__33612\
        );

    \I__6612\ : CascadeMux
    port map (
            O => \N__33616\,
            I => \N__33597\
        );

    \I__6611\ : InMux
    port map (
            O => \N__33615\,
            I => \N__33582\
        );

    \I__6610\ : InMux
    port map (
            O => \N__33612\,
            I => \N__33582\
        );

    \I__6609\ : InMux
    port map (
            O => \N__33611\,
            I => \N__33582\
        );

    \I__6608\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33573\
        );

    \I__6607\ : InMux
    port map (
            O => \N__33609\,
            I => \N__33573\
        );

    \I__6606\ : InMux
    port map (
            O => \N__33608\,
            I => \N__33573\
        );

    \I__6605\ : InMux
    port map (
            O => \N__33607\,
            I => \N__33573\
        );

    \I__6604\ : InMux
    port map (
            O => \N__33606\,
            I => \N__33562\
        );

    \I__6603\ : InMux
    port map (
            O => \N__33605\,
            I => \N__33562\
        );

    \I__6602\ : InMux
    port map (
            O => \N__33604\,
            I => \N__33542\
        );

    \I__6601\ : InMux
    port map (
            O => \N__33603\,
            I => \N__33542\
        );

    \I__6600\ : InMux
    port map (
            O => \N__33602\,
            I => \N__33529\
        );

    \I__6599\ : InMux
    port map (
            O => \N__33601\,
            I => \N__33529\
        );

    \I__6598\ : InMux
    port map (
            O => \N__33600\,
            I => \N__33529\
        );

    \I__6597\ : InMux
    port map (
            O => \N__33597\,
            I => \N__33529\
        );

    \I__6596\ : InMux
    port map (
            O => \N__33596\,
            I => \N__33529\
        );

    \I__6595\ : InMux
    port map (
            O => \N__33595\,
            I => \N__33529\
        );

    \I__6594\ : InMux
    port map (
            O => \N__33594\,
            I => \N__33518\
        );

    \I__6593\ : InMux
    port map (
            O => \N__33593\,
            I => \N__33518\
        );

    \I__6592\ : InMux
    port map (
            O => \N__33592\,
            I => \N__33518\
        );

    \I__6591\ : InMux
    port map (
            O => \N__33591\,
            I => \N__33518\
        );

    \I__6590\ : InMux
    port map (
            O => \N__33590\,
            I => \N__33518\
        );

    \I__6589\ : InMux
    port map (
            O => \N__33589\,
            I => \N__33512\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__33582\,
            I => \N__33509\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__33573\,
            I => \N__33506\
        );

    \I__6586\ : InMux
    port map (
            O => \N__33572\,
            I => \N__33493\
        );

    \I__6585\ : InMux
    port map (
            O => \N__33571\,
            I => \N__33493\
        );

    \I__6584\ : InMux
    port map (
            O => \N__33570\,
            I => \N__33493\
        );

    \I__6583\ : InMux
    port map (
            O => \N__33569\,
            I => \N__33493\
        );

    \I__6582\ : InMux
    port map (
            O => \N__33568\,
            I => \N__33493\
        );

    \I__6581\ : InMux
    port map (
            O => \N__33567\,
            I => \N__33493\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__33562\,
            I => \N__33489\
        );

    \I__6579\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33486\
        );

    \I__6578\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33471\
        );

    \I__6577\ : InMux
    port map (
            O => \N__33559\,
            I => \N__33471\
        );

    \I__6576\ : InMux
    port map (
            O => \N__33558\,
            I => \N__33471\
        );

    \I__6575\ : InMux
    port map (
            O => \N__33557\,
            I => \N__33471\
        );

    \I__6574\ : InMux
    port map (
            O => \N__33556\,
            I => \N__33471\
        );

    \I__6573\ : InMux
    port map (
            O => \N__33555\,
            I => \N__33471\
        );

    \I__6572\ : InMux
    port map (
            O => \N__33554\,
            I => \N__33471\
        );

    \I__6571\ : InMux
    port map (
            O => \N__33553\,
            I => \N__33455\
        );

    \I__6570\ : InMux
    port map (
            O => \N__33552\,
            I => \N__33455\
        );

    \I__6569\ : InMux
    port map (
            O => \N__33551\,
            I => \N__33455\
        );

    \I__6568\ : InMux
    port map (
            O => \N__33550\,
            I => \N__33455\
        );

    \I__6567\ : InMux
    port map (
            O => \N__33549\,
            I => \N__33455\
        );

    \I__6566\ : InMux
    port map (
            O => \N__33548\,
            I => \N__33447\
        );

    \I__6565\ : InMux
    port map (
            O => \N__33547\,
            I => \N__33444\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__33542\,
            I => \N__33441\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__33529\,
            I => \N__33436\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__33518\,
            I => \N__33436\
        );

    \I__6561\ : InMux
    port map (
            O => \N__33517\,
            I => \N__33426\
        );

    \I__6560\ : InMux
    port map (
            O => \N__33516\,
            I => \N__33426\
        );

    \I__6559\ : InMux
    port map (
            O => \N__33515\,
            I => \N__33426\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__33512\,
            I => \N__33417\
        );

    \I__6557\ : Span4Mux_v
    port map (
            O => \N__33509\,
            I => \N__33417\
        );

    \I__6556\ : Span4Mux_v
    port map (
            O => \N__33506\,
            I => \N__33417\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__33493\,
            I => \N__33417\
        );

    \I__6554\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33414\
        );

    \I__6553\ : Span4Mux_v
    port map (
            O => \N__33489\,
            I => \N__33407\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__33486\,
            I => \N__33407\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__33471\,
            I => \N__33407\
        );

    \I__6550\ : InMux
    port map (
            O => \N__33470\,
            I => \N__33389\
        );

    \I__6549\ : InMux
    port map (
            O => \N__33469\,
            I => \N__33389\
        );

    \I__6548\ : InMux
    port map (
            O => \N__33468\,
            I => \N__33389\
        );

    \I__6547\ : InMux
    port map (
            O => \N__33467\,
            I => \N__33389\
        );

    \I__6546\ : InMux
    port map (
            O => \N__33466\,
            I => \N__33389\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__33455\,
            I => \N__33386\
        );

    \I__6544\ : InMux
    port map (
            O => \N__33454\,
            I => \N__33372\
        );

    \I__6543\ : InMux
    port map (
            O => \N__33453\,
            I => \N__33372\
        );

    \I__6542\ : InMux
    port map (
            O => \N__33452\,
            I => \N__33372\
        );

    \I__6541\ : InMux
    port map (
            O => \N__33451\,
            I => \N__33372\
        );

    \I__6540\ : InMux
    port map (
            O => \N__33450\,
            I => \N__33372\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__33447\,
            I => \N__33367\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__33444\,
            I => \N__33367\
        );

    \I__6537\ : Span4Mux_h
    port map (
            O => \N__33441\,
            I => \N__33364\
        );

    \I__6536\ : Span4Mux_v
    port map (
            O => \N__33436\,
            I => \N__33361\
        );

    \I__6535\ : InMux
    port map (
            O => \N__33435\,
            I => \N__33354\
        );

    \I__6534\ : InMux
    port map (
            O => \N__33434\,
            I => \N__33354\
        );

    \I__6533\ : InMux
    port map (
            O => \N__33433\,
            I => \N__33354\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__33426\,
            I => \N__33349\
        );

    \I__6531\ : Span4Mux_h
    port map (
            O => \N__33417\,
            I => \N__33349\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__33414\,
            I => \N__33344\
        );

    \I__6529\ : Span4Mux_v
    port map (
            O => \N__33407\,
            I => \N__33344\
        );

    \I__6528\ : InMux
    port map (
            O => \N__33406\,
            I => \N__33329\
        );

    \I__6527\ : InMux
    port map (
            O => \N__33405\,
            I => \N__33329\
        );

    \I__6526\ : InMux
    port map (
            O => \N__33404\,
            I => \N__33329\
        );

    \I__6525\ : InMux
    port map (
            O => \N__33403\,
            I => \N__33329\
        );

    \I__6524\ : InMux
    port map (
            O => \N__33402\,
            I => \N__33329\
        );

    \I__6523\ : InMux
    port map (
            O => \N__33401\,
            I => \N__33329\
        );

    \I__6522\ : InMux
    port map (
            O => \N__33400\,
            I => \N__33329\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__33389\,
            I => \N__33324\
        );

    \I__6520\ : Span4Mux_h
    port map (
            O => \N__33386\,
            I => \N__33324\
        );

    \I__6519\ : InMux
    port map (
            O => \N__33385\,
            I => \N__33317\
        );

    \I__6518\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33317\
        );

    \I__6517\ : InMux
    port map (
            O => \N__33383\,
            I => \N__33317\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__33372\,
            I => \N__33310\
        );

    \I__6515\ : Span4Mux_h
    port map (
            O => \N__33367\,
            I => \N__33310\
        );

    \I__6514\ : Span4Mux_v
    port map (
            O => \N__33364\,
            I => \N__33310\
        );

    \I__6513\ : Odrv4
    port map (
            O => \N__33361\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__33354\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6511\ : Odrv4
    port map (
            O => \N__33349\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6510\ : Odrv4
    port map (
            O => \N__33344\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__33329\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6508\ : Odrv4
    port map (
            O => \N__33324\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__33317\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6506\ : Odrv4
    port map (
            O => \N__33310\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__6505\ : CascadeMux
    port map (
            O => \N__33293\,
            I => \N__33282\
        );

    \I__6504\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33255\
        );

    \I__6503\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33242\
        );

    \I__6502\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33242\
        );

    \I__6501\ : InMux
    port map (
            O => \N__33289\,
            I => \N__33242\
        );

    \I__6500\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33242\
        );

    \I__6499\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33242\
        );

    \I__6498\ : InMux
    port map (
            O => \N__33286\,
            I => \N__33242\
        );

    \I__6497\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33235\
        );

    \I__6496\ : InMux
    port map (
            O => \N__33282\,
            I => \N__33235\
        );

    \I__6495\ : InMux
    port map (
            O => \N__33281\,
            I => \N__33235\
        );

    \I__6494\ : CascadeMux
    port map (
            O => \N__33280\,
            I => \N__33231\
        );

    \I__6493\ : CascadeMux
    port map (
            O => \N__33279\,
            I => \N__33225\
        );

    \I__6492\ : CascadeMux
    port map (
            O => \N__33278\,
            I => \N__33215\
        );

    \I__6491\ : CascadeMux
    port map (
            O => \N__33277\,
            I => \N__33212\
        );

    \I__6490\ : CascadeMux
    port map (
            O => \N__33276\,
            I => \N__33205\
        );

    \I__6489\ : CascadeMux
    port map (
            O => \N__33275\,
            I => \N__33202\
        );

    \I__6488\ : CascadeMux
    port map (
            O => \N__33274\,
            I => \N__33199\
        );

    \I__6487\ : InMux
    port map (
            O => \N__33273\,
            I => \N__33194\
        );

    \I__6486\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33194\
        );

    \I__6485\ : CascadeMux
    port map (
            O => \N__33271\,
            I => \N__33188\
        );

    \I__6484\ : CascadeMux
    port map (
            O => \N__33270\,
            I => \N__33181\
        );

    \I__6483\ : CascadeMux
    port map (
            O => \N__33269\,
            I => \N__33176\
        );

    \I__6482\ : CascadeMux
    port map (
            O => \N__33268\,
            I => \N__33173\
        );

    \I__6481\ : CascadeMux
    port map (
            O => \N__33267\,
            I => \N__33170\
        );

    \I__6480\ : CascadeMux
    port map (
            O => \N__33266\,
            I => \N__33162\
        );

    \I__6479\ : CascadeMux
    port map (
            O => \N__33265\,
            I => \N__33157\
        );

    \I__6478\ : CascadeMux
    port map (
            O => \N__33264\,
            I => \N__33153\
        );

    \I__6477\ : CascadeMux
    port map (
            O => \N__33263\,
            I => \N__33149\
        );

    \I__6476\ : CascadeMux
    port map (
            O => \N__33262\,
            I => \N__33144\
        );

    \I__6475\ : CascadeMux
    port map (
            O => \N__33261\,
            I => \N__33140\
        );

    \I__6474\ : CascadeMux
    port map (
            O => \N__33260\,
            I => \N__33136\
        );

    \I__6473\ : CascadeMux
    port map (
            O => \N__33259\,
            I => \N__33132\
        );

    \I__6472\ : CascadeMux
    port map (
            O => \N__33258\,
            I => \N__33115\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__33255\,
            I => \N__33111\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__33242\,
            I => \N__33106\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__33235\,
            I => \N__33106\
        );

    \I__6468\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33103\
        );

    \I__6467\ : InMux
    port map (
            O => \N__33231\,
            I => \N__33092\
        );

    \I__6466\ : InMux
    port map (
            O => \N__33230\,
            I => \N__33092\
        );

    \I__6465\ : InMux
    port map (
            O => \N__33229\,
            I => \N__33092\
        );

    \I__6464\ : InMux
    port map (
            O => \N__33228\,
            I => \N__33092\
        );

    \I__6463\ : InMux
    port map (
            O => \N__33225\,
            I => \N__33092\
        );

    \I__6462\ : InMux
    port map (
            O => \N__33224\,
            I => \N__33087\
        );

    \I__6461\ : InMux
    port map (
            O => \N__33223\,
            I => \N__33087\
        );

    \I__6460\ : CascadeMux
    port map (
            O => \N__33222\,
            I => \N__33083\
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__33221\,
            I => \N__33080\
        );

    \I__6458\ : CascadeMux
    port map (
            O => \N__33220\,
            I => \N__33076\
        );

    \I__6457\ : CascadeMux
    port map (
            O => \N__33219\,
            I => \N__33072\
        );

    \I__6456\ : CascadeMux
    port map (
            O => \N__33218\,
            I => \N__33069\
        );

    \I__6455\ : InMux
    port map (
            O => \N__33215\,
            I => \N__33060\
        );

    \I__6454\ : InMux
    port map (
            O => \N__33212\,
            I => \N__33060\
        );

    \I__6453\ : InMux
    port map (
            O => \N__33211\,
            I => \N__33045\
        );

    \I__6452\ : InMux
    port map (
            O => \N__33210\,
            I => \N__33045\
        );

    \I__6451\ : InMux
    port map (
            O => \N__33209\,
            I => \N__33045\
        );

    \I__6450\ : InMux
    port map (
            O => \N__33208\,
            I => \N__33045\
        );

    \I__6449\ : InMux
    port map (
            O => \N__33205\,
            I => \N__33045\
        );

    \I__6448\ : InMux
    port map (
            O => \N__33202\,
            I => \N__33045\
        );

    \I__6447\ : InMux
    port map (
            O => \N__33199\,
            I => \N__33045\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__33194\,
            I => \N__33042\
        );

    \I__6445\ : CascadeMux
    port map (
            O => \N__33193\,
            I => \N__33038\
        );

    \I__6444\ : CascadeMux
    port map (
            O => \N__33192\,
            I => \N__33034\
        );

    \I__6443\ : CascadeMux
    port map (
            O => \N__33191\,
            I => \N__33030\
        );

    \I__6442\ : InMux
    port map (
            O => \N__33188\,
            I => \N__33024\
        );

    \I__6441\ : InMux
    port map (
            O => \N__33187\,
            I => \N__33024\
        );

    \I__6440\ : InMux
    port map (
            O => \N__33186\,
            I => \N__33011\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33185\,
            I => \N__33011\
        );

    \I__6438\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33011\
        );

    \I__6437\ : InMux
    port map (
            O => \N__33181\,
            I => \N__33011\
        );

    \I__6436\ : InMux
    port map (
            O => \N__33180\,
            I => \N__33011\
        );

    \I__6435\ : InMux
    port map (
            O => \N__33179\,
            I => \N__33011\
        );

    \I__6434\ : InMux
    port map (
            O => \N__33176\,
            I => \N__33004\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33173\,
            I => \N__33004\
        );

    \I__6432\ : InMux
    port map (
            O => \N__33170\,
            I => \N__33004\
        );

    \I__6431\ : InMux
    port map (
            O => \N__33169\,
            I => \N__32991\
        );

    \I__6430\ : InMux
    port map (
            O => \N__33168\,
            I => \N__32991\
        );

    \I__6429\ : InMux
    port map (
            O => \N__33167\,
            I => \N__32991\
        );

    \I__6428\ : InMux
    port map (
            O => \N__33166\,
            I => \N__32991\
        );

    \I__6427\ : InMux
    port map (
            O => \N__33165\,
            I => \N__32991\
        );

    \I__6426\ : InMux
    port map (
            O => \N__33162\,
            I => \N__32991\
        );

    \I__6425\ : InMux
    port map (
            O => \N__33161\,
            I => \N__32974\
        );

    \I__6424\ : InMux
    port map (
            O => \N__33160\,
            I => \N__32974\
        );

    \I__6423\ : InMux
    port map (
            O => \N__33157\,
            I => \N__32974\
        );

    \I__6422\ : InMux
    port map (
            O => \N__33156\,
            I => \N__32974\
        );

    \I__6421\ : InMux
    port map (
            O => \N__33153\,
            I => \N__32974\
        );

    \I__6420\ : InMux
    port map (
            O => \N__33152\,
            I => \N__32974\
        );

    \I__6419\ : InMux
    port map (
            O => \N__33149\,
            I => \N__32974\
        );

    \I__6418\ : InMux
    port map (
            O => \N__33148\,
            I => \N__32974\
        );

    \I__6417\ : InMux
    port map (
            O => \N__33147\,
            I => \N__32957\
        );

    \I__6416\ : InMux
    port map (
            O => \N__33144\,
            I => \N__32957\
        );

    \I__6415\ : InMux
    port map (
            O => \N__33143\,
            I => \N__32957\
        );

    \I__6414\ : InMux
    port map (
            O => \N__33140\,
            I => \N__32957\
        );

    \I__6413\ : InMux
    port map (
            O => \N__33139\,
            I => \N__32957\
        );

    \I__6412\ : InMux
    port map (
            O => \N__33136\,
            I => \N__32957\
        );

    \I__6411\ : InMux
    port map (
            O => \N__33135\,
            I => \N__32957\
        );

    \I__6410\ : InMux
    port map (
            O => \N__33132\,
            I => \N__32957\
        );

    \I__6409\ : CascadeMux
    port map (
            O => \N__33131\,
            I => \N__32954\
        );

    \I__6408\ : CascadeMux
    port map (
            O => \N__33130\,
            I => \N__32950\
        );

    \I__6407\ : CascadeMux
    port map (
            O => \N__33129\,
            I => \N__32946\
        );

    \I__6406\ : CascadeMux
    port map (
            O => \N__33128\,
            I => \N__32942\
        );

    \I__6405\ : CascadeMux
    port map (
            O => \N__33127\,
            I => \N__32937\
        );

    \I__6404\ : CascadeMux
    port map (
            O => \N__33126\,
            I => \N__32933\
        );

    \I__6403\ : CascadeMux
    port map (
            O => \N__33125\,
            I => \N__32929\
        );

    \I__6402\ : CascadeMux
    port map (
            O => \N__33124\,
            I => \N__32925\
        );

    \I__6401\ : CascadeMux
    port map (
            O => \N__33123\,
            I => \N__32921\
        );

    \I__6400\ : CascadeMux
    port map (
            O => \N__33122\,
            I => \N__32917\
        );

    \I__6399\ : CascadeMux
    port map (
            O => \N__33121\,
            I => \N__32913\
        );

    \I__6398\ : InMux
    port map (
            O => \N__33120\,
            I => \N__32899\
        );

    \I__6397\ : InMux
    port map (
            O => \N__33119\,
            I => \N__32899\
        );

    \I__6396\ : InMux
    port map (
            O => \N__33118\,
            I => \N__32899\
        );

    \I__6395\ : InMux
    port map (
            O => \N__33115\,
            I => \N__32899\
        );

    \I__6394\ : InMux
    port map (
            O => \N__33114\,
            I => \N__32899\
        );

    \I__6393\ : Span4Mux_v
    port map (
            O => \N__33111\,
            I => \N__32892\
        );

    \I__6392\ : Span4Mux_v
    port map (
            O => \N__33106\,
            I => \N__32892\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__33103\,
            I => \N__32892\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__33092\,
            I => \N__32889\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__33087\,
            I => \N__32886\
        );

    \I__6388\ : InMux
    port map (
            O => \N__33086\,
            I => \N__32883\
        );

    \I__6387\ : InMux
    port map (
            O => \N__33083\,
            I => \N__32878\
        );

    \I__6386\ : InMux
    port map (
            O => \N__33080\,
            I => \N__32878\
        );

    \I__6385\ : InMux
    port map (
            O => \N__33079\,
            I => \N__32867\
        );

    \I__6384\ : InMux
    port map (
            O => \N__33076\,
            I => \N__32867\
        );

    \I__6383\ : InMux
    port map (
            O => \N__33075\,
            I => \N__32867\
        );

    \I__6382\ : InMux
    port map (
            O => \N__33072\,
            I => \N__32867\
        );

    \I__6381\ : InMux
    port map (
            O => \N__33069\,
            I => \N__32867\
        );

    \I__6380\ : CascadeMux
    port map (
            O => \N__33068\,
            I => \N__32864\
        );

    \I__6379\ : CascadeMux
    port map (
            O => \N__33067\,
            I => \N__32860\
        );

    \I__6378\ : CascadeMux
    port map (
            O => \N__33066\,
            I => \N__32856\
        );

    \I__6377\ : CascadeMux
    port map (
            O => \N__33065\,
            I => \N__32852\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__33060\,
            I => \N__32848\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__33045\,
            I => \N__32843\
        );

    \I__6374\ : Span4Mux_v
    port map (
            O => \N__33042\,
            I => \N__32843\
        );

    \I__6373\ : InMux
    port map (
            O => \N__33041\,
            I => \N__32828\
        );

    \I__6372\ : InMux
    port map (
            O => \N__33038\,
            I => \N__32828\
        );

    \I__6371\ : InMux
    port map (
            O => \N__33037\,
            I => \N__32828\
        );

    \I__6370\ : InMux
    port map (
            O => \N__33034\,
            I => \N__32828\
        );

    \I__6369\ : InMux
    port map (
            O => \N__33033\,
            I => \N__32828\
        );

    \I__6368\ : InMux
    port map (
            O => \N__33030\,
            I => \N__32828\
        );

    \I__6367\ : InMux
    port map (
            O => \N__33029\,
            I => \N__32828\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__33024\,
            I => \N__32815\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__33011\,
            I => \N__32815\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__33004\,
            I => \N__32815\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__32991\,
            I => \N__32815\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__32974\,
            I => \N__32815\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__32957\,
            I => \N__32815\
        );

    \I__6360\ : InMux
    port map (
            O => \N__32954\,
            I => \N__32798\
        );

    \I__6359\ : InMux
    port map (
            O => \N__32953\,
            I => \N__32798\
        );

    \I__6358\ : InMux
    port map (
            O => \N__32950\,
            I => \N__32798\
        );

    \I__6357\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32798\
        );

    \I__6356\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32798\
        );

    \I__6355\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32798\
        );

    \I__6354\ : InMux
    port map (
            O => \N__32942\,
            I => \N__32798\
        );

    \I__6353\ : InMux
    port map (
            O => \N__32941\,
            I => \N__32798\
        );

    \I__6352\ : InMux
    port map (
            O => \N__32940\,
            I => \N__32781\
        );

    \I__6351\ : InMux
    port map (
            O => \N__32937\,
            I => \N__32781\
        );

    \I__6350\ : InMux
    port map (
            O => \N__32936\,
            I => \N__32781\
        );

    \I__6349\ : InMux
    port map (
            O => \N__32933\,
            I => \N__32781\
        );

    \I__6348\ : InMux
    port map (
            O => \N__32932\,
            I => \N__32781\
        );

    \I__6347\ : InMux
    port map (
            O => \N__32929\,
            I => \N__32781\
        );

    \I__6346\ : InMux
    port map (
            O => \N__32928\,
            I => \N__32781\
        );

    \I__6345\ : InMux
    port map (
            O => \N__32925\,
            I => \N__32781\
        );

    \I__6344\ : InMux
    port map (
            O => \N__32924\,
            I => \N__32768\
        );

    \I__6343\ : InMux
    port map (
            O => \N__32921\,
            I => \N__32768\
        );

    \I__6342\ : InMux
    port map (
            O => \N__32920\,
            I => \N__32768\
        );

    \I__6341\ : InMux
    port map (
            O => \N__32917\,
            I => \N__32768\
        );

    \I__6340\ : InMux
    port map (
            O => \N__32916\,
            I => \N__32768\
        );

    \I__6339\ : InMux
    port map (
            O => \N__32913\,
            I => \N__32768\
        );

    \I__6338\ : CascadeMux
    port map (
            O => \N__32912\,
            I => \N__32765\
        );

    \I__6337\ : CascadeMux
    port map (
            O => \N__32911\,
            I => \N__32761\
        );

    \I__6336\ : CascadeMux
    port map (
            O => \N__32910\,
            I => \N__32757\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__32899\,
            I => \N__32753\
        );

    \I__6334\ : Span4Mux_v
    port map (
            O => \N__32892\,
            I => \N__32750\
        );

    \I__6333\ : Span4Mux_h
    port map (
            O => \N__32889\,
            I => \N__32747\
        );

    \I__6332\ : Span4Mux_v
    port map (
            O => \N__32886\,
            I => \N__32738\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__32883\,
            I => \N__32738\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__32878\,
            I => \N__32738\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__32867\,
            I => \N__32738\
        );

    \I__6328\ : InMux
    port map (
            O => \N__32864\,
            I => \N__32721\
        );

    \I__6327\ : InMux
    port map (
            O => \N__32863\,
            I => \N__32721\
        );

    \I__6326\ : InMux
    port map (
            O => \N__32860\,
            I => \N__32721\
        );

    \I__6325\ : InMux
    port map (
            O => \N__32859\,
            I => \N__32721\
        );

    \I__6324\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32721\
        );

    \I__6323\ : InMux
    port map (
            O => \N__32855\,
            I => \N__32721\
        );

    \I__6322\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32721\
        );

    \I__6321\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32721\
        );

    \I__6320\ : Span4Mux_h
    port map (
            O => \N__32848\,
            I => \N__32706\
        );

    \I__6319\ : Span4Mux_h
    port map (
            O => \N__32843\,
            I => \N__32706\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__32828\,
            I => \N__32706\
        );

    \I__6317\ : Span4Mux_v
    port map (
            O => \N__32815\,
            I => \N__32706\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__32798\,
            I => \N__32706\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__32781\,
            I => \N__32706\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__32768\,
            I => \N__32706\
        );

    \I__6313\ : InMux
    port map (
            O => \N__32765\,
            I => \N__32693\
        );

    \I__6312\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32693\
        );

    \I__6311\ : InMux
    port map (
            O => \N__32761\,
            I => \N__32693\
        );

    \I__6310\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32693\
        );

    \I__6309\ : InMux
    port map (
            O => \N__32757\,
            I => \N__32693\
        );

    \I__6308\ : InMux
    port map (
            O => \N__32756\,
            I => \N__32693\
        );

    \I__6307\ : Odrv12
    port map (
            O => \N__32753\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__32750\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6305\ : Odrv4
    port map (
            O => \N__32747\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6304\ : Odrv4
    port map (
            O => \N__32738\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__32721\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6302\ : Odrv4
    port map (
            O => \N__32706\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__32693\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__6300\ : CascadeMux
    port map (
            O => \N__32678\,
            I => \N__32675\
        );

    \I__6299\ : InMux
    port map (
            O => \N__32675\,
            I => \N__32671\
        );

    \I__6298\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32668\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__32671\,
            I => \N__32662\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__32668\,
            I => \N__32662\
        );

    \I__6295\ : InMux
    port map (
            O => \N__32667\,
            I => \N__32659\
        );

    \I__6294\ : Span4Mux_h
    port map (
            O => \N__32662\,
            I => \N__32656\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__32659\,
            I => \N__32653\
        );

    \I__6292\ : Span4Mux_h
    port map (
            O => \N__32656\,
            I => \N__32649\
        );

    \I__6291\ : Span4Mux_h
    port map (
            O => \N__32653\,
            I => \N__32646\
        );

    \I__6290\ : InMux
    port map (
            O => \N__32652\,
            I => \N__32643\
        );

    \I__6289\ : Odrv4
    port map (
            O => \N__32649\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__6288\ : Odrv4
    port map (
            O => \N__32646\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__32643\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__6286\ : InMux
    port map (
            O => \N__32636\,
            I => \N__32633\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__32633\,
            I => \N__32629\
        );

    \I__6284\ : InMux
    port map (
            O => \N__32632\,
            I => \N__32626\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__32629\,
            I => \N__32620\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__32626\,
            I => \N__32620\
        );

    \I__6281\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32617\
        );

    \I__6280\ : Odrv4
    port map (
            O => \N__32620\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__32617\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__6278\ : InMux
    port map (
            O => \N__32612\,
            I => \N__32609\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__32609\,
            I => \N__32606\
        );

    \I__6276\ : Span4Mux_h
    port map (
            O => \N__32606\,
            I => \N__32603\
        );

    \I__6275\ : Odrv4
    port map (
            O => \N__32603\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__6274\ : IoInMux
    port map (
            O => \N__32600\,
            I => \N__32597\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__32597\,
            I => \N__32594\
        );

    \I__6272\ : Span12Mux_s0_v
    port map (
            O => \N__32594\,
            I => \N__32591\
        );

    \I__6271\ : Odrv12
    port map (
            O => \N__32591\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__6270\ : CEMux
    port map (
            O => \N__32588\,
            I => \N__32585\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__32585\,
            I => \N__32579\
        );

    \I__6268\ : CEMux
    port map (
            O => \N__32584\,
            I => \N__32576\
        );

    \I__6267\ : CEMux
    port map (
            O => \N__32583\,
            I => \N__32573\
        );

    \I__6266\ : CEMux
    port map (
            O => \N__32582\,
            I => \N__32570\
        );

    \I__6265\ : Span4Mux_v
    port map (
            O => \N__32579\,
            I => \N__32565\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__32576\,
            I => \N__32565\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__32573\,
            I => \N__32562\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__32570\,
            I => \N__32559\
        );

    \I__6261\ : Span4Mux_v
    port map (
            O => \N__32565\,
            I => \N__32556\
        );

    \I__6260\ : Span4Mux_h
    port map (
            O => \N__32562\,
            I => \N__32551\
        );

    \I__6259\ : Span4Mux_v
    port map (
            O => \N__32559\,
            I => \N__32551\
        );

    \I__6258\ : Sp12to4
    port map (
            O => \N__32556\,
            I => \N__32548\
        );

    \I__6257\ : Span4Mux_h
    port map (
            O => \N__32551\,
            I => \N__32545\
        );

    \I__6256\ : Odrv12
    port map (
            O => \N__32548\,
            I => \current_shift_inst.timer_s1.N_163_i\
        );

    \I__6255\ : Odrv4
    port map (
            O => \N__32545\,
            I => \current_shift_inst.timer_s1.N_163_i\
        );

    \I__6254\ : CascadeMux
    port map (
            O => \N__32540\,
            I => \N__32537\
        );

    \I__6253\ : InMux
    port map (
            O => \N__32537\,
            I => \N__32534\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__32534\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__6251\ : CascadeMux
    port map (
            O => \N__32531\,
            I => \N__32528\
        );

    \I__6250\ : InMux
    port map (
            O => \N__32528\,
            I => \N__32525\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__32525\,
            I => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\
        );

    \I__6248\ : InMux
    port map (
            O => \N__32522\,
            I => \N__32519\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__32519\,
            I => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\
        );

    \I__6246\ : InMux
    port map (
            O => \N__32516\,
            I => \N__32512\
        );

    \I__6245\ : InMux
    port map (
            O => \N__32515\,
            I => \N__32509\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__32512\,
            I => \N__32506\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__32509\,
            I => \N__32503\
        );

    \I__6242\ : Span4Mux_v
    port map (
            O => \N__32506\,
            I => \N__32500\
        );

    \I__6241\ : Span4Mux_h
    port map (
            O => \N__32503\,
            I => \N__32496\
        );

    \I__6240\ : Span4Mux_h
    port map (
            O => \N__32500\,
            I => \N__32493\
        );

    \I__6239\ : InMux
    port map (
            O => \N__32499\,
            I => \N__32490\
        );

    \I__6238\ : Odrv4
    port map (
            O => \N__32496\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__6237\ : Odrv4
    port map (
            O => \N__32493\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__32490\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__6235\ : CascadeMux
    port map (
            O => \N__32483\,
            I => \N__32479\
        );

    \I__6234\ : CascadeMux
    port map (
            O => \N__32482\,
            I => \N__32476\
        );

    \I__6233\ : InMux
    port map (
            O => \N__32479\,
            I => \N__32473\
        );

    \I__6232\ : InMux
    port map (
            O => \N__32476\,
            I => \N__32470\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__32473\,
            I => \N__32467\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__32470\,
            I => \N__32464\
        );

    \I__6229\ : Span4Mux_v
    port map (
            O => \N__32467\,
            I => \N__32461\
        );

    \I__6228\ : Span4Mux_h
    port map (
            O => \N__32464\,
            I => \N__32456\
        );

    \I__6227\ : Span4Mux_v
    port map (
            O => \N__32461\,
            I => \N__32453\
        );

    \I__6226\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32450\
        );

    \I__6225\ : InMux
    port map (
            O => \N__32459\,
            I => \N__32447\
        );

    \I__6224\ : Span4Mux_h
    port map (
            O => \N__32456\,
            I => \N__32444\
        );

    \I__6223\ : Sp12to4
    port map (
            O => \N__32453\,
            I => \N__32437\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__32450\,
            I => \N__32437\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__32447\,
            I => \N__32437\
        );

    \I__6220\ : Odrv4
    port map (
            O => \N__32444\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__6219\ : Odrv12
    port map (
            O => \N__32437\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__6218\ : InMux
    port map (
            O => \N__32432\,
            I => \N__32429\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__32429\,
            I => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\
        );

    \I__6216\ : InMux
    port map (
            O => \N__32426\,
            I => \N__32423\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__32423\,
            I => \N__32419\
        );

    \I__6214\ : InMux
    port map (
            O => \N__32422\,
            I => \N__32415\
        );

    \I__6213\ : Span4Mux_v
    port map (
            O => \N__32419\,
            I => \N__32412\
        );

    \I__6212\ : InMux
    port map (
            O => \N__32418\,
            I => \N__32409\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__32415\,
            I => \N__32406\
        );

    \I__6210\ : Span4Mux_h
    port map (
            O => \N__32412\,
            I => \N__32401\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__32409\,
            I => \N__32401\
        );

    \I__6208\ : Span12Mux_v
    port map (
            O => \N__32406\,
            I => \N__32397\
        );

    \I__6207\ : Span4Mux_v
    port map (
            O => \N__32401\,
            I => \N__32394\
        );

    \I__6206\ : InMux
    port map (
            O => \N__32400\,
            I => \N__32391\
        );

    \I__6205\ : Odrv12
    port map (
            O => \N__32397\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__6204\ : Odrv4
    port map (
            O => \N__32394\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__32391\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__6202\ : CascadeMux
    port map (
            O => \N__32384\,
            I => \N__32381\
        );

    \I__6201\ : InMux
    port map (
            O => \N__32381\,
            I => \N__32378\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__32378\,
            I => \N__32375\
        );

    \I__6199\ : Span4Mux_v
    port map (
            O => \N__32375\,
            I => \N__32371\
        );

    \I__6198\ : InMux
    port map (
            O => \N__32374\,
            I => \N__32368\
        );

    \I__6197\ : Span4Mux_h
    port map (
            O => \N__32371\,
            I => \N__32363\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__32368\,
            I => \N__32363\
        );

    \I__6195\ : Span4Mux_h
    port map (
            O => \N__32363\,
            I => \N__32359\
        );

    \I__6194\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32356\
        );

    \I__6193\ : Odrv4
    port map (
            O => \N__32359\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__32356\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__6191\ : CascadeMux
    port map (
            O => \N__32351\,
            I => \N__32348\
        );

    \I__6190\ : InMux
    port map (
            O => \N__32348\,
            I => \N__32345\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__32345\,
            I => \N__32342\
        );

    \I__6188\ : Odrv4
    port map (
            O => \N__32342\,
            I => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\
        );

    \I__6187\ : InMux
    port map (
            O => \N__32339\,
            I => \N__32335\
        );

    \I__6186\ : InMux
    port map (
            O => \N__32338\,
            I => \N__32332\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__32335\,
            I => \N__32329\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__32332\,
            I => \N__32325\
        );

    \I__6183\ : Span4Mux_h
    port map (
            O => \N__32329\,
            I => \N__32322\
        );

    \I__6182\ : InMux
    port map (
            O => \N__32328\,
            I => \N__32319\
        );

    \I__6181\ : Span4Mux_h
    port map (
            O => \N__32325\,
            I => \N__32315\
        );

    \I__6180\ : Span4Mux_v
    port map (
            O => \N__32322\,
            I => \N__32310\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__32319\,
            I => \N__32310\
        );

    \I__6178\ : InMux
    port map (
            O => \N__32318\,
            I => \N__32307\
        );

    \I__6177\ : Span4Mux_v
    port map (
            O => \N__32315\,
            I => \N__32302\
        );

    \I__6176\ : Span4Mux_h
    port map (
            O => \N__32310\,
            I => \N__32302\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__32307\,
            I => \N__32299\
        );

    \I__6174\ : Odrv4
    port map (
            O => \N__32302\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__6173\ : Odrv4
    port map (
            O => \N__32299\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__6172\ : InMux
    port map (
            O => \N__32294\,
            I => \N__32291\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__32291\,
            I => \N__32287\
        );

    \I__6170\ : InMux
    port map (
            O => \N__32290\,
            I => \N__32284\
        );

    \I__6169\ : Span4Mux_h
    port map (
            O => \N__32287\,
            I => \N__32280\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__32284\,
            I => \N__32277\
        );

    \I__6167\ : InMux
    port map (
            O => \N__32283\,
            I => \N__32274\
        );

    \I__6166\ : Odrv4
    port map (
            O => \N__32280\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__6165\ : Odrv4
    port map (
            O => \N__32277\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__32274\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__6163\ : CascadeMux
    port map (
            O => \N__32267\,
            I => \N__32264\
        );

    \I__6162\ : InMux
    port map (
            O => \N__32264\,
            I => \N__32261\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__32261\,
            I => \N__32258\
        );

    \I__6160\ : Span4Mux_h
    port map (
            O => \N__32258\,
            I => \N__32255\
        );

    \I__6159\ : Odrv4
    port map (
            O => \N__32255\,
            I => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\
        );

    \I__6158\ : CascadeMux
    port map (
            O => \N__32252\,
            I => \N__32249\
        );

    \I__6157\ : InMux
    port map (
            O => \N__32249\,
            I => \N__32245\
        );

    \I__6156\ : InMux
    port map (
            O => \N__32248\,
            I => \N__32242\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__32245\,
            I => \N__32239\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__32242\,
            I => \N__32235\
        );

    \I__6153\ : Span4Mux_h
    port map (
            O => \N__32239\,
            I => \N__32231\
        );

    \I__6152\ : InMux
    port map (
            O => \N__32238\,
            I => \N__32228\
        );

    \I__6151\ : Span4Mux_h
    port map (
            O => \N__32235\,
            I => \N__32225\
        );

    \I__6150\ : InMux
    port map (
            O => \N__32234\,
            I => \N__32222\
        );

    \I__6149\ : Span4Mux_v
    port map (
            O => \N__32231\,
            I => \N__32219\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__32228\,
            I => \N__32216\
        );

    \I__6147\ : Span4Mux_v
    port map (
            O => \N__32225\,
            I => \N__32211\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__32222\,
            I => \N__32211\
        );

    \I__6145\ : Span4Mux_h
    port map (
            O => \N__32219\,
            I => \N__32208\
        );

    \I__6144\ : Span4Mux_h
    port map (
            O => \N__32216\,
            I => \N__32205\
        );

    \I__6143\ : Span4Mux_h
    port map (
            O => \N__32211\,
            I => \N__32202\
        );

    \I__6142\ : Odrv4
    port map (
            O => \N__32208\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__6141\ : Odrv4
    port map (
            O => \N__32205\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__6140\ : Odrv4
    port map (
            O => \N__32202\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__6139\ : InMux
    port map (
            O => \N__32195\,
            I => \N__32191\
        );

    \I__6138\ : InMux
    port map (
            O => \N__32194\,
            I => \N__32188\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__32191\,
            I => \N__32184\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__32188\,
            I => \N__32181\
        );

    \I__6135\ : InMux
    port map (
            O => \N__32187\,
            I => \N__32178\
        );

    \I__6134\ : Span4Mux_v
    port map (
            O => \N__32184\,
            I => \N__32175\
        );

    \I__6133\ : Span4Mux_h
    port map (
            O => \N__32181\,
            I => \N__32170\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__32178\,
            I => \N__32170\
        );

    \I__6131\ : Odrv4
    port map (
            O => \N__32175\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__6130\ : Odrv4
    port map (
            O => \N__32170\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__6129\ : InMux
    port map (
            O => \N__32165\,
            I => \N__32162\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__32162\,
            I => \N__32159\
        );

    \I__6127\ : Odrv4
    port map (
            O => \N__32159\,
            I => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\
        );

    \I__6126\ : InMux
    port map (
            O => \N__32156\,
            I => \N__32152\
        );

    \I__6125\ : InMux
    port map (
            O => \N__32155\,
            I => \N__32149\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__32152\,
            I => \N__32144\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__32149\,
            I => \N__32144\
        );

    \I__6122\ : Span4Mux_v
    port map (
            O => \N__32144\,
            I => \N__32140\
        );

    \I__6121\ : InMux
    port map (
            O => \N__32143\,
            I => \N__32136\
        );

    \I__6120\ : Span4Mux_v
    port map (
            O => \N__32140\,
            I => \N__32133\
        );

    \I__6119\ : InMux
    port map (
            O => \N__32139\,
            I => \N__32130\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__32136\,
            I => \N__32127\
        );

    \I__6117\ : Span4Mux_h
    port map (
            O => \N__32133\,
            I => \N__32122\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__32130\,
            I => \N__32122\
        );

    \I__6115\ : Odrv12
    port map (
            O => \N__32127\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__6114\ : Odrv4
    port map (
            O => \N__32122\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__6113\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32114\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__32114\,
            I => \N__32109\
        );

    \I__6111\ : InMux
    port map (
            O => \N__32113\,
            I => \N__32106\
        );

    \I__6110\ : InMux
    port map (
            O => \N__32112\,
            I => \N__32103\
        );

    \I__6109\ : Span4Mux_h
    port map (
            O => \N__32109\,
            I => \N__32098\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__32106\,
            I => \N__32098\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__32103\,
            I => \N__32095\
        );

    \I__6106\ : Span4Mux_v
    port map (
            O => \N__32098\,
            I => \N__32092\
        );

    \I__6105\ : Span4Mux_h
    port map (
            O => \N__32095\,
            I => \N__32089\
        );

    \I__6104\ : Odrv4
    port map (
            O => \N__32092\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__6103\ : Odrv4
    port map (
            O => \N__32089\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__6102\ : CascadeMux
    port map (
            O => \N__32084\,
            I => \N__32081\
        );

    \I__6101\ : InMux
    port map (
            O => \N__32081\,
            I => \N__32078\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__32078\,
            I => \N__32075\
        );

    \I__6099\ : Odrv4
    port map (
            O => \N__32075\,
            I => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\
        );

    \I__6098\ : InMux
    port map (
            O => \N__32072\,
            I => \N__32069\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__32069\,
            I => \N__32066\
        );

    \I__6096\ : Span4Mux_h
    port map (
            O => \N__32066\,
            I => \N__32063\
        );

    \I__6095\ : Sp12to4
    port map (
            O => \N__32063\,
            I => \N__32060\
        );

    \I__6094\ : Span12Mux_v
    port map (
            O => \N__32060\,
            I => \N__32057\
        );

    \I__6093\ : Odrv12
    port map (
            O => \N__32057\,
            I => \il_max_comp1_D1\
        );

    \I__6092\ : InMux
    port map (
            O => \N__32054\,
            I => \N__32050\
        );

    \I__6091\ : InMux
    port map (
            O => \N__32053\,
            I => \N__32047\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__32050\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__32047\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\
        );

    \I__6088\ : InMux
    port map (
            O => \N__32042\,
            I => \N__32036\
        );

    \I__6087\ : InMux
    port map (
            O => \N__32041\,
            I => \N__32036\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__32036\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\
        );

    \I__6085\ : InMux
    port map (
            O => \N__32033\,
            I => \N__32030\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__32030\,
            I => \N__32027\
        );

    \I__6083\ : Odrv12
    port map (
            O => \N__32027\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df30\
        );

    \I__6082\ : InMux
    port map (
            O => \N__32024\,
            I => \N__32015\
        );

    \I__6081\ : InMux
    port map (
            O => \N__32023\,
            I => \N__32015\
        );

    \I__6080\ : InMux
    port map (
            O => \N__32022\,
            I => \N__32015\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__32015\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\
        );

    \I__6078\ : CascadeMux
    port map (
            O => \N__32012\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\
        );

    \I__6077\ : InMux
    port map (
            O => \N__32009\,
            I => \N__32006\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__32006\,
            I => \N__32003\
        );

    \I__6075\ : Span4Mux_h
    port map (
            O => \N__32003\,
            I => \N__32000\
        );

    \I__6074\ : Span4Mux_v
    port map (
            O => \N__32000\,
            I => \N__31996\
        );

    \I__6073\ : InMux
    port map (
            O => \N__31999\,
            I => \N__31993\
        );

    \I__6072\ : Odrv4
    port map (
            O => \N__31996\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__31993\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__6070\ : CascadeMux
    port map (
            O => \N__31988\,
            I => \N__31985\
        );

    \I__6069\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31979\
        );

    \I__6068\ : InMux
    port map (
            O => \N__31984\,
            I => \N__31974\
        );

    \I__6067\ : InMux
    port map (
            O => \N__31983\,
            I => \N__31974\
        );

    \I__6066\ : InMux
    port map (
            O => \N__31982\,
            I => \N__31971\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__31979\,
            I => \N__31968\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__31974\,
            I => \N__31965\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__31971\,
            I => \N__31962\
        );

    \I__6062\ : Span4Mux_v
    port map (
            O => \N__31968\,
            I => \N__31959\
        );

    \I__6061\ : Span4Mux_h
    port map (
            O => \N__31965\,
            I => \N__31955\
        );

    \I__6060\ : Span12Mux_v
    port map (
            O => \N__31962\,
            I => \N__31952\
        );

    \I__6059\ : Span4Mux_h
    port map (
            O => \N__31959\,
            I => \N__31949\
        );

    \I__6058\ : InMux
    port map (
            O => \N__31958\,
            I => \N__31946\
        );

    \I__6057\ : Span4Mux_h
    port map (
            O => \N__31955\,
            I => \N__31943\
        );

    \I__6056\ : Odrv12
    port map (
            O => \N__31952\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__6055\ : Odrv4
    port map (
            O => \N__31949\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__31946\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__6053\ : Odrv4
    port map (
            O => \N__31943\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__6052\ : InMux
    port map (
            O => \N__31934\,
            I => \N__31928\
        );

    \I__6051\ : InMux
    port map (
            O => \N__31933\,
            I => \N__31928\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__31928\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__6049\ : CascadeMux
    port map (
            O => \N__31925\,
            I => \N__31922\
        );

    \I__6048\ : InMux
    port map (
            O => \N__31922\,
            I => \N__31918\
        );

    \I__6047\ : InMux
    port map (
            O => \N__31921\,
            I => \N__31915\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__31918\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__31915\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__6044\ : InMux
    port map (
            O => \N__31910\,
            I => \N__31907\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__31907\,
            I => \N__31903\
        );

    \I__6042\ : InMux
    port map (
            O => \N__31906\,
            I => \N__31900\
        );

    \I__6041\ : Odrv4
    port map (
            O => \N__31903\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__31900\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__31895\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\
        );

    \I__6038\ : InMux
    port map (
            O => \N__31892\,
            I => \N__31885\
        );

    \I__6037\ : InMux
    port map (
            O => \N__31891\,
            I => \N__31885\
        );

    \I__6036\ : InMux
    port map (
            O => \N__31890\,
            I => \N__31882\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__31885\,
            I => \N__31879\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__31882\,
            I => \N__31873\
        );

    \I__6033\ : Span4Mux_v
    port map (
            O => \N__31879\,
            I => \N__31873\
        );

    \I__6032\ : InMux
    port map (
            O => \N__31878\,
            I => \N__31870\
        );

    \I__6031\ : Span4Mux_h
    port map (
            O => \N__31873\,
            I => \N__31865\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__31870\,
            I => \N__31865\
        );

    \I__6029\ : Span4Mux_v
    port map (
            O => \N__31865\,
            I => \N__31862\
        );

    \I__6028\ : Odrv4
    port map (
            O => \N__31862\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__6027\ : InMux
    port map (
            O => \N__31859\,
            I => \N__31856\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__31856\,
            I => \N__31853\
        );

    \I__6025\ : Span4Mux_h
    port map (
            O => \N__31853\,
            I => \N__31849\
        );

    \I__6024\ : InMux
    port map (
            O => \N__31852\,
            I => \N__31846\
        );

    \I__6023\ : Odrv4
    port map (
            O => \N__31849\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__31846\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\
        );

    \I__6021\ : InMux
    port map (
            O => \N__31841\,
            I => \N__31838\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__31838\,
            I => \N__31834\
        );

    \I__6019\ : InMux
    port map (
            O => \N__31837\,
            I => \N__31831\
        );

    \I__6018\ : Span4Mux_v
    port map (
            O => \N__31834\,
            I => \N__31825\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__31831\,
            I => \N__31825\
        );

    \I__6016\ : InMux
    port map (
            O => \N__31830\,
            I => \N__31822\
        );

    \I__6015\ : Span4Mux_v
    port map (
            O => \N__31825\,
            I => \N__31819\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__31822\,
            I => \N__31816\
        );

    \I__6013\ : Sp12to4
    port map (
            O => \N__31819\,
            I => \N__31813\
        );

    \I__6012\ : Span12Mux_v
    port map (
            O => \N__31816\,
            I => \N__31808\
        );

    \I__6011\ : Span12Mux_h
    port map (
            O => \N__31813\,
            I => \N__31808\
        );

    \I__6010\ : Odrv12
    port map (
            O => \N__31808\,
            I => il_min_comp2_c
        );

    \I__6009\ : InMux
    port map (
            O => \N__31805\,
            I => \N__31802\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__31802\,
            I => \N__31796\
        );

    \I__6007\ : InMux
    port map (
            O => \N__31801\,
            I => \N__31793\
        );

    \I__6006\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31790\
        );

    \I__6005\ : InMux
    port map (
            O => \N__31799\,
            I => \N__31787\
        );

    \I__6004\ : Span4Mux_v
    port map (
            O => \N__31796\,
            I => \N__31784\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__31793\,
            I => \N__31781\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__31790\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__31787\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__6000\ : Odrv4
    port map (
            O => \N__31784\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__5999\ : Odrv12
    port map (
            O => \N__31781\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__5998\ : CascadeMux
    port map (
            O => \N__31772\,
            I => \N__31769\
        );

    \I__5997\ : InMux
    port map (
            O => \N__31769\,
            I => \N__31765\
        );

    \I__5996\ : InMux
    port map (
            O => \N__31768\,
            I => \N__31762\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__31765\,
            I => \N__31758\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__31762\,
            I => \N__31755\
        );

    \I__5993\ : CascadeMux
    port map (
            O => \N__31761\,
            I => \N__31752\
        );

    \I__5992\ : Span4Mux_h
    port map (
            O => \N__31758\,
            I => \N__31749\
        );

    \I__5991\ : Span4Mux_v
    port map (
            O => \N__31755\,
            I => \N__31746\
        );

    \I__5990\ : InMux
    port map (
            O => \N__31752\,
            I => \N__31743\
        );

    \I__5989\ : Span4Mux_v
    port map (
            O => \N__31749\,
            I => \N__31738\
        );

    \I__5988\ : Span4Mux_h
    port map (
            O => \N__31746\,
            I => \N__31738\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__31743\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__5986\ : Odrv4
    port map (
            O => \N__31738\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__5985\ : InMux
    port map (
            O => \N__31733\,
            I => \N__31728\
        );

    \I__5984\ : InMux
    port map (
            O => \N__31732\,
            I => \N__31725\
        );

    \I__5983\ : InMux
    port map (
            O => \N__31731\,
            I => \N__31722\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__31728\,
            I => \N__31719\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__31725\,
            I => \N__31716\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__31722\,
            I => \N__31712\
        );

    \I__5979\ : Span4Mux_h
    port map (
            O => \N__31719\,
            I => \N__31709\
        );

    \I__5978\ : Span12Mux_s4_v
    port map (
            O => \N__31716\,
            I => \N__31706\
        );

    \I__5977\ : InMux
    port map (
            O => \N__31715\,
            I => \N__31703\
        );

    \I__5976\ : Span4Mux_h
    port map (
            O => \N__31712\,
            I => \N__31698\
        );

    \I__5975\ : Span4Mux_v
    port map (
            O => \N__31709\,
            I => \N__31698\
        );

    \I__5974\ : Span12Mux_v
    port map (
            O => \N__31706\,
            I => \N__31695\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__31703\,
            I => \N__31690\
        );

    \I__5972\ : Span4Mux_v
    port map (
            O => \N__31698\,
            I => \N__31690\
        );

    \I__5971\ : Odrv12
    port map (
            O => \N__31695\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__5970\ : Odrv4
    port map (
            O => \N__31690\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__5969\ : InMux
    port map (
            O => \N__31685\,
            I => \N__31682\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__31682\,
            I => \N__31679\
        );

    \I__5967\ : Odrv12
    port map (
            O => \N__31679\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__5966\ : CascadeMux
    port map (
            O => \N__31676\,
            I => \phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_\
        );

    \I__5965\ : InMux
    port map (
            O => \N__31673\,
            I => \N__31667\
        );

    \I__5964\ : InMux
    port map (
            O => \N__31672\,
            I => \N__31667\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__31667\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__5962\ : CascadeMux
    port map (
            O => \N__31664\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__5961\ : CascadeMux
    port map (
            O => \N__31661\,
            I => \N__31656\
        );

    \I__5960\ : InMux
    port map (
            O => \N__31660\,
            I => \N__31653\
        );

    \I__5959\ : InMux
    port map (
            O => \N__31659\,
            I => \N__31648\
        );

    \I__5958\ : InMux
    port map (
            O => \N__31656\,
            I => \N__31648\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__31653\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__31648\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__5955\ : CascadeMux
    port map (
            O => \N__31643\,
            I => \N__31638\
        );

    \I__5954\ : InMux
    port map (
            O => \N__31642\,
            I => \N__31635\
        );

    \I__5953\ : InMux
    port map (
            O => \N__31641\,
            I => \N__31630\
        );

    \I__5952\ : InMux
    port map (
            O => \N__31638\,
            I => \N__31630\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__31635\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__31630\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__5949\ : InMux
    port map (
            O => \N__31625\,
            I => \N__31622\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__31622\,
            I => \N__31619\
        );

    \I__5947\ : Span4Mux_h
    port map (
            O => \N__31619\,
            I => \N__31616\
        );

    \I__5946\ : Odrv4
    port map (
            O => \N__31616\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\
        );

    \I__5945\ : InMux
    port map (
            O => \N__31613\,
            I => \N__31609\
        );

    \I__5944\ : InMux
    port map (
            O => \N__31612\,
            I => \N__31605\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__31609\,
            I => \N__31602\
        );

    \I__5942\ : InMux
    port map (
            O => \N__31608\,
            I => \N__31599\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__31605\,
            I => \N__31592\
        );

    \I__5940\ : Span12Mux_h
    port map (
            O => \N__31602\,
            I => \N__31592\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__31599\,
            I => \N__31592\
        );

    \I__5938\ : Odrv12
    port map (
            O => \N__31592\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__5937\ : InMux
    port map (
            O => \N__31589\,
            I => \N__31586\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__31586\,
            I => \N__31581\
        );

    \I__5935\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31578\
        );

    \I__5934\ : InMux
    port map (
            O => \N__31584\,
            I => \N__31575\
        );

    \I__5933\ : Span4Mux_v
    port map (
            O => \N__31581\,
            I => \N__31571\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__31578\,
            I => \N__31568\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__31575\,
            I => \N__31565\
        );

    \I__5930\ : InMux
    port map (
            O => \N__31574\,
            I => \N__31562\
        );

    \I__5929\ : Span4Mux_h
    port map (
            O => \N__31571\,
            I => \N__31555\
        );

    \I__5928\ : Span4Mux_h
    port map (
            O => \N__31568\,
            I => \N__31555\
        );

    \I__5927\ : Span4Mux_v
    port map (
            O => \N__31565\,
            I => \N__31555\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__31562\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__31555\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__5924\ : InMux
    port map (
            O => \N__31550\,
            I => \N__31544\
        );

    \I__5923\ : InMux
    port map (
            O => \N__31549\,
            I => \N__31544\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__31544\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\
        );

    \I__5921\ : InMux
    port map (
            O => \N__31541\,
            I => \N__31538\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__31538\,
            I => \N__31535\
        );

    \I__5919\ : Span4Mux_h
    port map (
            O => \N__31535\,
            I => \N__31530\
        );

    \I__5918\ : InMux
    port map (
            O => \N__31534\,
            I => \N__31527\
        );

    \I__5917\ : InMux
    port map (
            O => \N__31533\,
            I => \N__31524\
        );

    \I__5916\ : Span4Mux_h
    port map (
            O => \N__31530\,
            I => \N__31521\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__31527\,
            I => \N__31518\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__31524\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__5913\ : Odrv4
    port map (
            O => \N__31521\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__5912\ : Odrv4
    port map (
            O => \N__31518\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__5911\ : InMux
    port map (
            O => \N__31511\,
            I => \N__31507\
        );

    \I__5910\ : InMux
    port map (
            O => \N__31510\,
            I => \N__31504\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__31507\,
            I => \N__31499\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__31504\,
            I => \N__31496\
        );

    \I__5907\ : InMux
    port map (
            O => \N__31503\,
            I => \N__31493\
        );

    \I__5906\ : InMux
    port map (
            O => \N__31502\,
            I => \N__31490\
        );

    \I__5905\ : Span4Mux_v
    port map (
            O => \N__31499\,
            I => \N__31487\
        );

    \I__5904\ : Span4Mux_v
    port map (
            O => \N__31496\,
            I => \N__31482\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__31493\,
            I => \N__31482\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__31490\,
            I => \N__31479\
        );

    \I__5901\ : Span4Mux_h
    port map (
            O => \N__31487\,
            I => \N__31476\
        );

    \I__5900\ : Span4Mux_h
    port map (
            O => \N__31482\,
            I => \N__31471\
        );

    \I__5899\ : Span4Mux_v
    port map (
            O => \N__31479\,
            I => \N__31471\
        );

    \I__5898\ : Odrv4
    port map (
            O => \N__31476\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__5897\ : Odrv4
    port map (
            O => \N__31471\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__5896\ : InMux
    port map (
            O => \N__31466\,
            I => \N__31460\
        );

    \I__5895\ : InMux
    port map (
            O => \N__31465\,
            I => \N__31460\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__31460\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\
        );

    \I__5893\ : InMux
    port map (
            O => \N__31457\,
            I => \N__31454\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__31454\,
            I => \N__31451\
        );

    \I__5891\ : Span4Mux_h
    port map (
            O => \N__31451\,
            I => \N__31448\
        );

    \I__5890\ : Odrv4
    port map (
            O => \N__31448\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt20\
        );

    \I__5889\ : InMux
    port map (
            O => \N__31445\,
            I => \N__31440\
        );

    \I__5888\ : InMux
    port map (
            O => \N__31444\,
            I => \N__31435\
        );

    \I__5887\ : InMux
    port map (
            O => \N__31443\,
            I => \N__31435\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__31440\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__31435\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__5884\ : CascadeMux
    port map (
            O => \N__31430\,
            I => \N__31427\
        );

    \I__5883\ : InMux
    port map (
            O => \N__31427\,
            I => \N__31420\
        );

    \I__5882\ : InMux
    port map (
            O => \N__31426\,
            I => \N__31420\
        );

    \I__5881\ : InMux
    port map (
            O => \N__31425\,
            I => \N__31417\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__31420\,
            I => \N__31414\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__31417\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__5878\ : Odrv4
    port map (
            O => \N__31414\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__5877\ : CascadeMux
    port map (
            O => \N__31409\,
            I => \N__31406\
        );

    \I__5876\ : InMux
    port map (
            O => \N__31406\,
            I => \N__31403\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__31403\,
            I => \N__31400\
        );

    \I__5874\ : Span4Mux_h
    port map (
            O => \N__31400\,
            I => \N__31397\
        );

    \I__5873\ : Odrv4
    port map (
            O => \N__31397\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\
        );

    \I__5872\ : CascadeMux
    port map (
            O => \N__31394\,
            I => \N__31391\
        );

    \I__5871\ : InMux
    port map (
            O => \N__31391\,
            I => \N__31385\
        );

    \I__5870\ : InMux
    port map (
            O => \N__31390\,
            I => \N__31385\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__31385\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\
        );

    \I__5868\ : InMux
    port map (
            O => \N__31382\,
            I => \N__31379\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__31379\,
            I => \N__31375\
        );

    \I__5866\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31371\
        );

    \I__5865\ : Span12Mux_h
    port map (
            O => \N__31375\,
            I => \N__31368\
        );

    \I__5864\ : InMux
    port map (
            O => \N__31374\,
            I => \N__31365\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__31371\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__5862\ : Odrv12
    port map (
            O => \N__31368\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__31365\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__5860\ : InMux
    port map (
            O => \N__31358\,
            I => \N__31353\
        );

    \I__5859\ : InMux
    port map (
            O => \N__31357\,
            I => \N__31350\
        );

    \I__5858\ : InMux
    port map (
            O => \N__31356\,
            I => \N__31347\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__31353\,
            I => \N__31343\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__31350\,
            I => \N__31338\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__31347\,
            I => \N__31338\
        );

    \I__5854\ : CascadeMux
    port map (
            O => \N__31346\,
            I => \N__31335\
        );

    \I__5853\ : Span4Mux_v
    port map (
            O => \N__31343\,
            I => \N__31332\
        );

    \I__5852\ : Span4Mux_v
    port map (
            O => \N__31338\,
            I => \N__31329\
        );

    \I__5851\ : InMux
    port map (
            O => \N__31335\,
            I => \N__31326\
        );

    \I__5850\ : Span4Mux_h
    port map (
            O => \N__31332\,
            I => \N__31319\
        );

    \I__5849\ : Span4Mux_v
    port map (
            O => \N__31329\,
            I => \N__31319\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__31326\,
            I => \N__31319\
        );

    \I__5847\ : Span4Mux_v
    port map (
            O => \N__31319\,
            I => \N__31316\
        );

    \I__5846\ : Odrv4
    port map (
            O => \N__31316\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__5845\ : InMux
    port map (
            O => \N__31313\,
            I => \N__31307\
        );

    \I__5844\ : InMux
    port map (
            O => \N__31312\,
            I => \N__31307\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__31307\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\
        );

    \I__5842\ : InMux
    port map (
            O => \N__31304\,
            I => \N__31299\
        );

    \I__5841\ : InMux
    port map (
            O => \N__31303\,
            I => \N__31296\
        );

    \I__5840\ : InMux
    port map (
            O => \N__31302\,
            I => \N__31293\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__31299\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__31296\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__31293\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__5836\ : CascadeMux
    port map (
            O => \N__31286\,
            I => \N__31282\
        );

    \I__5835\ : CascadeMux
    port map (
            O => \N__31285\,
            I => \N__31279\
        );

    \I__5834\ : InMux
    port map (
            O => \N__31282\,
            I => \N__31276\
        );

    \I__5833\ : InMux
    port map (
            O => \N__31279\,
            I => \N__31273\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__31276\,
            I => \N__31270\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__31273\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\
        );

    \I__5830\ : Odrv12
    port map (
            O => \N__31270\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\
        );

    \I__5829\ : InMux
    port map (
            O => \N__31265\,
            I => \N__31260\
        );

    \I__5828\ : InMux
    port map (
            O => \N__31264\,
            I => \N__31257\
        );

    \I__5827\ : InMux
    port map (
            O => \N__31263\,
            I => \N__31254\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__31260\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__31257\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__31254\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__5823\ : CascadeMux
    port map (
            O => \N__31247\,
            I => \N__31244\
        );

    \I__5822\ : InMux
    port map (
            O => \N__31244\,
            I => \N__31241\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__31241\,
            I => \N__31238\
        );

    \I__5820\ : Odrv12
    port map (
            O => \N__31238\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\
        );

    \I__5819\ : InMux
    port map (
            O => \N__31235\,
            I => \N__31231\
        );

    \I__5818\ : InMux
    port map (
            O => \N__31234\,
            I => \N__31228\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__31231\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__31228\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__5815\ : InMux
    port map (
            O => \N__31223\,
            I => \N__31219\
        );

    \I__5814\ : InMux
    port map (
            O => \N__31222\,
            I => \N__31215\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__31219\,
            I => \N__31212\
        );

    \I__5812\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31209\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__31215\,
            I => \N__31206\
        );

    \I__5810\ : Span4Mux_h
    port map (
            O => \N__31212\,
            I => \N__31203\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__31209\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__5808\ : Odrv4
    port map (
            O => \N__31206\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__5807\ : Odrv4
    port map (
            O => \N__31203\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__5806\ : CascadeMux
    port map (
            O => \N__31196\,
            I => \N__31192\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__31195\,
            I => \N__31189\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31192\,
            I => \N__31186\
        );

    \I__5803\ : InMux
    port map (
            O => \N__31189\,
            I => \N__31183\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__31186\,
            I => \N__31180\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__31183\,
            I => \N__31177\
        );

    \I__5800\ : Span4Mux_h
    port map (
            O => \N__31180\,
            I => \N__31174\
        );

    \I__5799\ : Odrv4
    port map (
            O => \N__31177\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__5798\ : Odrv4
    port map (
            O => \N__31174\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__5797\ : InMux
    port map (
            O => \N__31169\,
            I => \N__31165\
        );

    \I__5796\ : InMux
    port map (
            O => \N__31168\,
            I => \N__31161\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__31165\,
            I => \N__31158\
        );

    \I__5794\ : InMux
    port map (
            O => \N__31164\,
            I => \N__31155\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__31161\,
            I => \N__31152\
        );

    \I__5792\ : Span4Mux_h
    port map (
            O => \N__31158\,
            I => \N__31149\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__31155\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__5790\ : Odrv4
    port map (
            O => \N__31152\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__5789\ : Odrv4
    port map (
            O => \N__31149\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__5788\ : CascadeMux
    port map (
            O => \N__31142\,
            I => \N__31139\
        );

    \I__5787\ : InMux
    port map (
            O => \N__31139\,
            I => \N__31136\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__31136\,
            I => \N__31133\
        );

    \I__5785\ : Span4Mux_v
    port map (
            O => \N__31133\,
            I => \N__31130\
        );

    \I__5784\ : Odrv4
    port map (
            O => \N__31130\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt16\
        );

    \I__5783\ : InMux
    port map (
            O => \N__31127\,
            I => \N__31118\
        );

    \I__5782\ : InMux
    port map (
            O => \N__31126\,
            I => \N__31118\
        );

    \I__5781\ : InMux
    port map (
            O => \N__31125\,
            I => \N__31118\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__31118\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__5779\ : CascadeMux
    port map (
            O => \N__31115\,
            I => \N__31112\
        );

    \I__5778\ : InMux
    port map (
            O => \N__31112\,
            I => \N__31108\
        );

    \I__5777\ : InMux
    port map (
            O => \N__31111\,
            I => \N__31105\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__31108\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__31105\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__5774\ : CascadeMux
    port map (
            O => \N__31100\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_\
        );

    \I__5773\ : InMux
    port map (
            O => \N__31097\,
            I => \N__31094\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__31094\,
            I => \N__31091\
        );

    \I__5771\ : Span4Mux_v
    port map (
            O => \N__31091\,
            I => \N__31088\
        );

    \I__5770\ : Odrv4
    port map (
            O => \N__31088\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa\
        );

    \I__5769\ : InMux
    port map (
            O => \N__31085\,
            I => \N__31082\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__31082\,
            I => \N__31079\
        );

    \I__5767\ : Span4Mux_v
    port map (
            O => \N__31079\,
            I => \N__31076\
        );

    \I__5766\ : Sp12to4
    port map (
            O => \N__31076\,
            I => \N__31073\
        );

    \I__5765\ : Span12Mux_h
    port map (
            O => \N__31073\,
            I => \N__31070\
        );

    \I__5764\ : Span12Mux_v
    port map (
            O => \N__31070\,
            I => \N__31064\
        );

    \I__5763\ : InMux
    port map (
            O => \N__31069\,
            I => \N__31057\
        );

    \I__5762\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31057\
        );

    \I__5761\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31057\
        );

    \I__5760\ : Odrv12
    port map (
            O => \N__31064\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__31057\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__5758\ : InMux
    port map (
            O => \N__31052\,
            I => \N__31043\
        );

    \I__5757\ : InMux
    port map (
            O => \N__31051\,
            I => \N__31043\
        );

    \I__5756\ : InMux
    port map (
            O => \N__31050\,
            I => \N__31043\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__31043\,
            I => \N__31040\
        );

    \I__5754\ : Span4Mux_v
    port map (
            O => \N__31040\,
            I => \N__31037\
        );

    \I__5753\ : Span4Mux_h
    port map (
            O => \N__31037\,
            I => \N__31034\
        );

    \I__5752\ : Span4Mux_h
    port map (
            O => \N__31034\,
            I => \N__31031\
        );

    \I__5751\ : Odrv4
    port map (
            O => \N__31031\,
            I => il_max_comp2_c
        );

    \I__5750\ : CascadeMux
    port map (
            O => \N__31028\,
            I => \N__31025\
        );

    \I__5749\ : InMux
    port map (
            O => \N__31025\,
            I => \N__31022\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__31022\,
            I => \N__31019\
        );

    \I__5747\ : Span4Mux_h
    port map (
            O => \N__31019\,
            I => \N__31016\
        );

    \I__5746\ : Odrv4
    port map (
            O => \N__31016\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt22\
        );

    \I__5745\ : CascadeMux
    port map (
            O => \N__31013\,
            I => \N__31010\
        );

    \I__5744\ : InMux
    port map (
            O => \N__31010\,
            I => \N__31007\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__31007\,
            I => \pwm_generator_inst.un14_counter_1\
        );

    \I__5742\ : CascadeMux
    port map (
            O => \N__31004\,
            I => \N__31001\
        );

    \I__5741\ : InMux
    port map (
            O => \N__31001\,
            I => \N__30998\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__30998\,
            I => \N__30995\
        );

    \I__5739\ : Odrv4
    port map (
            O => \N__30995\,
            I => \pwm_generator_inst.threshold_0\
        );

    \I__5738\ : CascadeMux
    port map (
            O => \N__30992\,
            I => \N__30989\
        );

    \I__5737\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30986\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__30986\,
            I => \pwm_generator_inst.threshold_2\
        );

    \I__5735\ : CascadeMux
    port map (
            O => \N__30983\,
            I => \N__30980\
        );

    \I__5734\ : InMux
    port map (
            O => \N__30980\,
            I => \N__30977\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__30977\,
            I => \N__30974\
        );

    \I__5732\ : Odrv4
    port map (
            O => \N__30974\,
            I => \pwm_generator_inst.un14_counter_8\
        );

    \I__5731\ : InMux
    port map (
            O => \N__30971\,
            I => \N__30947\
        );

    \I__5730\ : InMux
    port map (
            O => \N__30970\,
            I => \N__30947\
        );

    \I__5729\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30940\
        );

    \I__5728\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30940\
        );

    \I__5727\ : InMux
    port map (
            O => \N__30967\,
            I => \N__30940\
        );

    \I__5726\ : InMux
    port map (
            O => \N__30966\,
            I => \N__30922\
        );

    \I__5725\ : InMux
    port map (
            O => \N__30965\,
            I => \N__30922\
        );

    \I__5724\ : InMux
    port map (
            O => \N__30964\,
            I => \N__30922\
        );

    \I__5723\ : InMux
    port map (
            O => \N__30963\,
            I => \N__30922\
        );

    \I__5722\ : InMux
    port map (
            O => \N__30962\,
            I => \N__30922\
        );

    \I__5721\ : InMux
    port map (
            O => \N__30961\,
            I => \N__30922\
        );

    \I__5720\ : InMux
    port map (
            O => \N__30960\,
            I => \N__30922\
        );

    \I__5719\ : InMux
    port map (
            O => \N__30959\,
            I => \N__30922\
        );

    \I__5718\ : InMux
    port map (
            O => \N__30958\,
            I => \N__30907\
        );

    \I__5717\ : InMux
    port map (
            O => \N__30957\,
            I => \N__30907\
        );

    \I__5716\ : InMux
    port map (
            O => \N__30956\,
            I => \N__30907\
        );

    \I__5715\ : InMux
    port map (
            O => \N__30955\,
            I => \N__30907\
        );

    \I__5714\ : InMux
    port map (
            O => \N__30954\,
            I => \N__30907\
        );

    \I__5713\ : InMux
    port map (
            O => \N__30953\,
            I => \N__30907\
        );

    \I__5712\ : InMux
    port map (
            O => \N__30952\,
            I => \N__30907\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__30947\,
            I => \N__30904\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__30940\,
            I => \N__30901\
        );

    \I__5709\ : CascadeMux
    port map (
            O => \N__30939\,
            I => \N__30892\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__30922\,
            I => \N__30886\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__30907\,
            I => \N__30886\
        );

    \I__5706\ : Span4Mux_v
    port map (
            O => \N__30904\,
            I => \N__30881\
        );

    \I__5705\ : Span4Mux_v
    port map (
            O => \N__30901\,
            I => \N__30881\
        );

    \I__5704\ : CascadeMux
    port map (
            O => \N__30900\,
            I => \N__30878\
        );

    \I__5703\ : CascadeMux
    port map (
            O => \N__30899\,
            I => \N__30874\
        );

    \I__5702\ : CascadeMux
    port map (
            O => \N__30898\,
            I => \N__30871\
        );

    \I__5701\ : CascadeMux
    port map (
            O => \N__30897\,
            I => \N__30866\
        );

    \I__5700\ : CascadeMux
    port map (
            O => \N__30896\,
            I => \N__30863\
        );

    \I__5699\ : CascadeMux
    port map (
            O => \N__30895\,
            I => \N__30860\
        );

    \I__5698\ : InMux
    port map (
            O => \N__30892\,
            I => \N__30854\
        );

    \I__5697\ : InMux
    port map (
            O => \N__30891\,
            I => \N__30854\
        );

    \I__5696\ : Span12Mux_s10_v
    port map (
            O => \N__30886\,
            I => \N__30851\
        );

    \I__5695\ : Span4Mux_h
    port map (
            O => \N__30881\,
            I => \N__30848\
        );

    \I__5694\ : InMux
    port map (
            O => \N__30878\,
            I => \N__30845\
        );

    \I__5693\ : InMux
    port map (
            O => \N__30877\,
            I => \N__30832\
        );

    \I__5692\ : InMux
    port map (
            O => \N__30874\,
            I => \N__30832\
        );

    \I__5691\ : InMux
    port map (
            O => \N__30871\,
            I => \N__30832\
        );

    \I__5690\ : InMux
    port map (
            O => \N__30870\,
            I => \N__30832\
        );

    \I__5689\ : InMux
    port map (
            O => \N__30869\,
            I => \N__30832\
        );

    \I__5688\ : InMux
    port map (
            O => \N__30866\,
            I => \N__30832\
        );

    \I__5687\ : InMux
    port map (
            O => \N__30863\,
            I => \N__30825\
        );

    \I__5686\ : InMux
    port map (
            O => \N__30860\,
            I => \N__30825\
        );

    \I__5685\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30825\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__30854\,
            I => \N__30820\
        );

    \I__5683\ : Span12Mux_h
    port map (
            O => \N__30851\,
            I => \N__30820\
        );

    \I__5682\ : Sp12to4
    port map (
            O => \N__30848\,
            I => \N__30817\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__30845\,
            I => \N_19_1\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__30832\,
            I => \N_19_1\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__30825\,
            I => \N_19_1\
        );

    \I__5678\ : Odrv12
    port map (
            O => \N__30820\,
            I => \N_19_1\
        );

    \I__5677\ : Odrv12
    port map (
            O => \N__30817\,
            I => \N_19_1\
        );

    \I__5676\ : CascadeMux
    port map (
            O => \N__30806\,
            I => \N__30803\
        );

    \I__5675\ : InMux
    port map (
            O => \N__30803\,
            I => \N__30800\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__30800\,
            I => \pwm_generator_inst.threshold_9\
        );

    \I__5673\ : IoInMux
    port map (
            O => \N__30797\,
            I => \N__30794\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__30794\,
            I => \N__30791\
        );

    \I__5671\ : IoSpan4Mux
    port map (
            O => \N__30791\,
            I => \N__30788\
        );

    \I__5670\ : Span4Mux_s0_v
    port map (
            O => \N__30788\,
            I => \N__30785\
        );

    \I__5669\ : Odrv4
    port map (
            O => \N__30785\,
            I => \pll_inst.red_c_i\
        );

    \I__5668\ : InMux
    port map (
            O => \N__30782\,
            I => \N__30779\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__30779\,
            I => \N__30776\
        );

    \I__5666\ : Span4Mux_v
    port map (
            O => \N__30776\,
            I => \N__30773\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__30773\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\
        );

    \I__5664\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30764\
        );

    \I__5663\ : CascadeMux
    port map (
            O => \N__30769\,
            I => \N__30761\
        );

    \I__5662\ : InMux
    port map (
            O => \N__30768\,
            I => \N__30758\
        );

    \I__5661\ : InMux
    port map (
            O => \N__30767\,
            I => \N__30755\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__30764\,
            I => \N__30752\
        );

    \I__5659\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30749\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__30758\,
            I => \N__30746\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__30755\,
            I => \N__30741\
        );

    \I__5656\ : Span4Mux_h
    port map (
            O => \N__30752\,
            I => \N__30741\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__30749\,
            I => \N__30738\
        );

    \I__5654\ : Span12Mux_s11_v
    port map (
            O => \N__30746\,
            I => \N__30735\
        );

    \I__5653\ : Span4Mux_v
    port map (
            O => \N__30741\,
            I => \N__30730\
        );

    \I__5652\ : Span4Mux_h
    port map (
            O => \N__30738\,
            I => \N__30730\
        );

    \I__5651\ : Odrv12
    port map (
            O => \N__30735\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__5650\ : Odrv4
    port map (
            O => \N__30730\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__5649\ : InMux
    port map (
            O => \N__30725\,
            I => \N__30722\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__30722\,
            I => \N__30719\
        );

    \I__5647\ : Span4Mux_h
    port map (
            O => \N__30719\,
            I => \N__30715\
        );

    \I__5646\ : InMux
    port map (
            O => \N__30718\,
            I => \N__30711\
        );

    \I__5645\ : Span4Mux_h
    port map (
            O => \N__30715\,
            I => \N__30708\
        );

    \I__5644\ : InMux
    port map (
            O => \N__30714\,
            I => \N__30705\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__30711\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__30708\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__30705\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__5640\ : InMux
    port map (
            O => \N__30698\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__5639\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30692\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__30692\,
            I => \N__30689\
        );

    \I__5637\ : Span12Mux_s9_v
    port map (
            O => \N__30689\,
            I => \N__30686\
        );

    \I__5636\ : Span12Mux_h
    port map (
            O => \N__30686\,
            I => \N__30683\
        );

    \I__5635\ : Odrv12
    port map (
            O => \N__30683\,
            I => \pwm_generator_inst.un2_threshold_2_1_16\
        );

    \I__5634\ : InMux
    port map (
            O => \N__30680\,
            I => \N__30676\
        );

    \I__5633\ : InMux
    port map (
            O => \N__30679\,
            I => \N__30673\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__30676\,
            I => \N__30668\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__30673\,
            I => \N__30668\
        );

    \I__5630\ : Span4Mux_h
    port map (
            O => \N__30668\,
            I => \N__30665\
        );

    \I__5629\ : Span4Mux_h
    port map (
            O => \N__30665\,
            I => \N__30662\
        );

    \I__5628\ : Span4Mux_h
    port map (
            O => \N__30662\,
            I => \N__30659\
        );

    \I__5627\ : Odrv4
    port map (
            O => \N__30659\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__5626\ : CascadeMux
    port map (
            O => \N__30656\,
            I => \N__30653\
        );

    \I__5625\ : InMux
    port map (
            O => \N__30653\,
            I => \N__30650\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__30650\,
            I => \pwm_generator_inst.threshold_3\
        );

    \I__5623\ : CascadeMux
    port map (
            O => \N__30647\,
            I => \N__30644\
        );

    \I__5622\ : InMux
    port map (
            O => \N__30644\,
            I => \N__30641\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__30641\,
            I => \pwm_generator_inst.threshold_4\
        );

    \I__5620\ : CascadeMux
    port map (
            O => \N__30638\,
            I => \N__30635\
        );

    \I__5619\ : InMux
    port map (
            O => \N__30635\,
            I => \N__30632\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__30632\,
            I => \pwm_generator_inst.threshold_5\
        );

    \I__5617\ : CascadeMux
    port map (
            O => \N__30629\,
            I => \N__30626\
        );

    \I__5616\ : InMux
    port map (
            O => \N__30626\,
            I => \N__30623\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__30623\,
            I => \N__30620\
        );

    \I__5614\ : Odrv4
    port map (
            O => \N__30620\,
            I => \pwm_generator_inst.un14_counter_6\
        );

    \I__5613\ : CascadeMux
    port map (
            O => \N__30617\,
            I => \N__30614\
        );

    \I__5612\ : InMux
    port map (
            O => \N__30614\,
            I => \N__30611\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__30611\,
            I => \pwm_generator_inst.un14_counter_7\
        );

    \I__5610\ : InMux
    port map (
            O => \N__30608\,
            I => \bfn_12_21_0_\
        );

    \I__5609\ : InMux
    port map (
            O => \N__30605\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__5608\ : InMux
    port map (
            O => \N__30602\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__5607\ : InMux
    port map (
            O => \N__30599\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__5606\ : InMux
    port map (
            O => \N__30596\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__5605\ : InMux
    port map (
            O => \N__30593\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__5604\ : InMux
    port map (
            O => \N__30590\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__5603\ : InMux
    port map (
            O => \N__30587\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__5602\ : InMux
    port map (
            O => \N__30584\,
            I => \bfn_12_22_0_\
        );

    \I__5601\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30577\
        );

    \I__5600\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30574\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__30577\,
            I => \N__30570\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__30574\,
            I => \N__30567\
        );

    \I__5597\ : InMux
    port map (
            O => \N__30573\,
            I => \N__30564\
        );

    \I__5596\ : Span4Mux_h
    port map (
            O => \N__30570\,
            I => \N__30561\
        );

    \I__5595\ : Span4Mux_v
    port map (
            O => \N__30567\,
            I => \N__30556\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__30564\,
            I => \N__30556\
        );

    \I__5593\ : Span4Mux_h
    port map (
            O => \N__30561\,
            I => \N__30552\
        );

    \I__5592\ : Span4Mux_h
    port map (
            O => \N__30556\,
            I => \N__30549\
        );

    \I__5591\ : InMux
    port map (
            O => \N__30555\,
            I => \N__30546\
        );

    \I__5590\ : Odrv4
    port map (
            O => \N__30552\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__5589\ : Odrv4
    port map (
            O => \N__30549\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__30546\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__5587\ : CascadeMux
    port map (
            O => \N__30539\,
            I => \N__30535\
        );

    \I__5586\ : InMux
    port map (
            O => \N__30538\,
            I => \N__30532\
        );

    \I__5585\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30529\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__30532\,
            I => \N__30526\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__30529\,
            I => \N__30522\
        );

    \I__5582\ : Span4Mux_h
    port map (
            O => \N__30526\,
            I => \N__30519\
        );

    \I__5581\ : InMux
    port map (
            O => \N__30525\,
            I => \N__30516\
        );

    \I__5580\ : Odrv4
    port map (
            O => \N__30522\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__5579\ : Odrv4
    port map (
            O => \N__30519\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__30516\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__5577\ : InMux
    port map (
            O => \N__30509\,
            I => \N__30506\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__30506\,
            I => \N__30503\
        );

    \I__5575\ : Odrv4
    port map (
            O => \N__30503\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__5574\ : InMux
    port map (
            O => \N__30500\,
            I => \N__30496\
        );

    \I__5573\ : InMux
    port map (
            O => \N__30499\,
            I => \N__30492\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__30496\,
            I => \N__30488\
        );

    \I__5571\ : InMux
    port map (
            O => \N__30495\,
            I => \N__30485\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__30492\,
            I => \N__30482\
        );

    \I__5569\ : InMux
    port map (
            O => \N__30491\,
            I => \N__30479\
        );

    \I__5568\ : Span4Mux_v
    port map (
            O => \N__30488\,
            I => \N__30476\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__30485\,
            I => \N__30473\
        );

    \I__5566\ : Span4Mux_h
    port map (
            O => \N__30482\,
            I => \N__30468\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__30479\,
            I => \N__30468\
        );

    \I__5564\ : Span4Mux_h
    port map (
            O => \N__30476\,
            I => \N__30465\
        );

    \I__5563\ : Span4Mux_h
    port map (
            O => \N__30473\,
            I => \N__30462\
        );

    \I__5562\ : Span4Mux_h
    port map (
            O => \N__30468\,
            I => \N__30459\
        );

    \I__5561\ : Odrv4
    port map (
            O => \N__30465\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__5560\ : Odrv4
    port map (
            O => \N__30462\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__5559\ : Odrv4
    port map (
            O => \N__30459\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__5558\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30447\
        );

    \I__5557\ : InMux
    port map (
            O => \N__30451\,
            I => \N__30444\
        );

    \I__5556\ : InMux
    port map (
            O => \N__30450\,
            I => \N__30441\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__30447\,
            I => \N__30438\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__30444\,
            I => \N__30435\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__30441\,
            I => \N__30432\
        );

    \I__5552\ : Odrv4
    port map (
            O => \N__30438\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__5551\ : Odrv4
    port map (
            O => \N__30435\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__5550\ : Odrv4
    port map (
            O => \N__30432\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__5549\ : InMux
    port map (
            O => \N__30425\,
            I => \N__30422\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__30422\,
            I => \N__30419\
        );

    \I__5547\ : Odrv12
    port map (
            O => \N__30419\,
            I => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\
        );

    \I__5546\ : CascadeMux
    port map (
            O => \N__30416\,
            I => \N__30413\
        );

    \I__5545\ : InMux
    port map (
            O => \N__30413\,
            I => \N__30409\
        );

    \I__5544\ : InMux
    port map (
            O => \N__30412\,
            I => \N__30406\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__30409\,
            I => \N__30400\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__30406\,
            I => \N__30400\
        );

    \I__5541\ : InMux
    port map (
            O => \N__30405\,
            I => \N__30397\
        );

    \I__5540\ : Span4Mux_h
    port map (
            O => \N__30400\,
            I => \N__30393\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__30397\,
            I => \N__30390\
        );

    \I__5538\ : InMux
    port map (
            O => \N__30396\,
            I => \N__30387\
        );

    \I__5537\ : Span4Mux_h
    port map (
            O => \N__30393\,
            I => \N__30384\
        );

    \I__5536\ : Span4Mux_v
    port map (
            O => \N__30390\,
            I => \N__30379\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__30387\,
            I => \N__30379\
        );

    \I__5534\ : Odrv4
    port map (
            O => \N__30384\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__5533\ : Odrv4
    port map (
            O => \N__30379\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__5532\ : InMux
    port map (
            O => \N__30374\,
            I => \N__30371\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__30371\,
            I => \N__30366\
        );

    \I__5530\ : InMux
    port map (
            O => \N__30370\,
            I => \N__30363\
        );

    \I__5529\ : InMux
    port map (
            O => \N__30369\,
            I => \N__30360\
        );

    \I__5528\ : Odrv4
    port map (
            O => \N__30366\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__30363\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__30360\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__5525\ : CascadeMux
    port map (
            O => \N__30353\,
            I => \N__30350\
        );

    \I__5524\ : InMux
    port map (
            O => \N__30350\,
            I => \N__30347\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__30347\,
            I => \N__30344\
        );

    \I__5522\ : Span4Mux_v
    port map (
            O => \N__30344\,
            I => \N__30341\
        );

    \I__5521\ : Odrv4
    port map (
            O => \N__30341\,
            I => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\
        );

    \I__5520\ : CascadeMux
    port map (
            O => \N__30338\,
            I => \N__30334\
        );

    \I__5519\ : CascadeMux
    port map (
            O => \N__30337\,
            I => \N__30331\
        );

    \I__5518\ : InMux
    port map (
            O => \N__30334\,
            I => \N__30328\
        );

    \I__5517\ : InMux
    port map (
            O => \N__30331\,
            I => \N__30324\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__30328\,
            I => \N__30321\
        );

    \I__5515\ : InMux
    port map (
            O => \N__30327\,
            I => \N__30318\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__30324\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__5513\ : Odrv4
    port map (
            O => \N__30321\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__30318\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__5511\ : InMux
    port map (
            O => \N__30311\,
            I => \N__30307\
        );

    \I__5510\ : InMux
    port map (
            O => \N__30310\,
            I => \N__30304\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__30307\,
            I => \N__30300\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__30304\,
            I => \N__30297\
        );

    \I__5507\ : InMux
    port map (
            O => \N__30303\,
            I => \N__30294\
        );

    \I__5506\ : Span4Mux_v
    port map (
            O => \N__30300\,
            I => \N__30287\
        );

    \I__5505\ : Span4Mux_h
    port map (
            O => \N__30297\,
            I => \N__30287\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__30294\,
            I => \N__30287\
        );

    \I__5503\ : Span4Mux_h
    port map (
            O => \N__30287\,
            I => \N__30283\
        );

    \I__5502\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30280\
        );

    \I__5501\ : Odrv4
    port map (
            O => \N__30283\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__30280\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__5499\ : CascadeMux
    port map (
            O => \N__30275\,
            I => \N__30272\
        );

    \I__5498\ : InMux
    port map (
            O => \N__30272\,
            I => \N__30269\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__30269\,
            I => \N__30266\
        );

    \I__5496\ : Span4Mux_v
    port map (
            O => \N__30266\,
            I => \N__30263\
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__30263\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__5494\ : CascadeMux
    port map (
            O => \N__30260\,
            I => \N__30256\
        );

    \I__5493\ : InMux
    port map (
            O => \N__30259\,
            I => \N__30253\
        );

    \I__5492\ : InMux
    port map (
            O => \N__30256\,
            I => \N__30250\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__30253\,
            I => \N__30246\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__30250\,
            I => \N__30243\
        );

    \I__5489\ : InMux
    port map (
            O => \N__30249\,
            I => \N__30240\
        );

    \I__5488\ : Span4Mux_v
    port map (
            O => \N__30246\,
            I => \N__30237\
        );

    \I__5487\ : Span4Mux_h
    port map (
            O => \N__30243\,
            I => \N__30231\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__30240\,
            I => \N__30231\
        );

    \I__5485\ : Span4Mux_v
    port map (
            O => \N__30237\,
            I => \N__30228\
        );

    \I__5484\ : InMux
    port map (
            O => \N__30236\,
            I => \N__30225\
        );

    \I__5483\ : Span4Mux_h
    port map (
            O => \N__30231\,
            I => \N__30222\
        );

    \I__5482\ : Span4Mux_v
    port map (
            O => \N__30228\,
            I => \N__30217\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__30225\,
            I => \N__30217\
        );

    \I__5480\ : Odrv4
    port map (
            O => \N__30222\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__5479\ : Odrv4
    port map (
            O => \N__30217\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__5478\ : InMux
    port map (
            O => \N__30212\,
            I => \N__30209\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__30209\,
            I => \N__30206\
        );

    \I__5476\ : Span4Mux_h
    port map (
            O => \N__30206\,
            I => \N__30203\
        );

    \I__5475\ : Span4Mux_v
    port map (
            O => \N__30203\,
            I => \N__30199\
        );

    \I__5474\ : InMux
    port map (
            O => \N__30202\,
            I => \N__30196\
        );

    \I__5473\ : Span4Mux_v
    port map (
            O => \N__30199\,
            I => \N__30190\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__30196\,
            I => \N__30190\
        );

    \I__5471\ : InMux
    port map (
            O => \N__30195\,
            I => \N__30187\
        );

    \I__5470\ : Odrv4
    port map (
            O => \N__30190\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__30187\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__5468\ : InMux
    port map (
            O => \N__30182\,
            I => \N__30179\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__30179\,
            I => \N__30176\
        );

    \I__5466\ : Span4Mux_v
    port map (
            O => \N__30176\,
            I => \N__30173\
        );

    \I__5465\ : Odrv4
    port map (
            O => \N__30173\,
            I => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\
        );

    \I__5464\ : CascadeMux
    port map (
            O => \N__30170\,
            I => \N__30165\
        );

    \I__5463\ : InMux
    port map (
            O => \N__30169\,
            I => \N__30160\
        );

    \I__5462\ : InMux
    port map (
            O => \N__30168\,
            I => \N__30160\
        );

    \I__5461\ : InMux
    port map (
            O => \N__30165\,
            I => \N__30156\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__30160\,
            I => \N__30153\
        );

    \I__5459\ : InMux
    port map (
            O => \N__30159\,
            I => \N__30150\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__30156\,
            I => \N__30147\
        );

    \I__5457\ : Span4Mux_v
    port map (
            O => \N__30153\,
            I => \N__30142\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__30150\,
            I => \N__30142\
        );

    \I__5455\ : Span12Mux_h
    port map (
            O => \N__30147\,
            I => \N__30139\
        );

    \I__5454\ : Span4Mux_h
    port map (
            O => \N__30142\,
            I => \N__30136\
        );

    \I__5453\ : Odrv12
    port map (
            O => \N__30139\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__30136\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__5451\ : InMux
    port map (
            O => \N__30131\,
            I => \N__30127\
        );

    \I__5450\ : InMux
    port map (
            O => \N__30130\,
            I => \N__30123\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__30127\,
            I => \N__30120\
        );

    \I__5448\ : InMux
    port map (
            O => \N__30126\,
            I => \N__30117\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__30123\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__5446\ : Odrv4
    port map (
            O => \N__30120\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__30117\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__5444\ : CascadeMux
    port map (
            O => \N__30110\,
            I => \N__30107\
        );

    \I__5443\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30104\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__30104\,
            I => \N__30101\
        );

    \I__5441\ : Span4Mux_v
    port map (
            O => \N__30101\,
            I => \N__30098\
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__30098\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__5439\ : InMux
    port map (
            O => \N__30095\,
            I => \N__30091\
        );

    \I__5438\ : InMux
    port map (
            O => \N__30094\,
            I => \N__30087\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__30091\,
            I => \N__30084\
        );

    \I__5436\ : InMux
    port map (
            O => \N__30090\,
            I => \N__30081\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__30087\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__5434\ : Odrv4
    port map (
            O => \N__30084\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__30081\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__5432\ : InMux
    port map (
            O => \N__30074\,
            I => \N__30070\
        );

    \I__5431\ : CascadeMux
    port map (
            O => \N__30073\,
            I => \N__30066\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__30070\,
            I => \N__30063\
        );

    \I__5429\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30060\
        );

    \I__5428\ : InMux
    port map (
            O => \N__30066\,
            I => \N__30057\
        );

    \I__5427\ : Span4Mux_h
    port map (
            O => \N__30063\,
            I => \N__30053\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__30060\,
            I => \N__30050\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__30057\,
            I => \N__30047\
        );

    \I__5424\ : InMux
    port map (
            O => \N__30056\,
            I => \N__30044\
        );

    \I__5423\ : Span4Mux_h
    port map (
            O => \N__30053\,
            I => \N__30041\
        );

    \I__5422\ : Span4Mux_h
    port map (
            O => \N__30050\,
            I => \N__30038\
        );

    \I__5421\ : Span4Mux_v
    port map (
            O => \N__30047\,
            I => \N__30033\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__30044\,
            I => \N__30033\
        );

    \I__5419\ : Odrv4
    port map (
            O => \N__30041\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__5418\ : Odrv4
    port map (
            O => \N__30038\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__5417\ : Odrv4
    port map (
            O => \N__30033\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__5416\ : InMux
    port map (
            O => \N__30026\,
            I => \N__30023\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__30023\,
            I => \N__30020\
        );

    \I__5414\ : Span4Mux_v
    port map (
            O => \N__30020\,
            I => \N__30017\
        );

    \I__5413\ : Odrv4
    port map (
            O => \N__30017\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__5412\ : CascadeMux
    port map (
            O => \N__30014\,
            I => \N__30011\
        );

    \I__5411\ : InMux
    port map (
            O => \N__30011\,
            I => \N__30008\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__30008\,
            I => \N__30002\
        );

    \I__5409\ : InMux
    port map (
            O => \N__30007\,
            I => \N__29999\
        );

    \I__5408\ : InMux
    port map (
            O => \N__30006\,
            I => \N__29996\
        );

    \I__5407\ : InMux
    port map (
            O => \N__30005\,
            I => \N__29993\
        );

    \I__5406\ : Span4Mux_v
    port map (
            O => \N__30002\,
            I => \N__29990\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__29999\,
            I => \N__29987\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__29996\,
            I => \N__29982\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__29993\,
            I => \N__29982\
        );

    \I__5402\ : Span4Mux_h
    port map (
            O => \N__29990\,
            I => \N__29977\
        );

    \I__5401\ : Span4Mux_v
    port map (
            O => \N__29987\,
            I => \N__29977\
        );

    \I__5400\ : Span4Mux_v
    port map (
            O => \N__29982\,
            I => \N__29974\
        );

    \I__5399\ : Odrv4
    port map (
            O => \N__29977\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__5398\ : Odrv4
    port map (
            O => \N__29974\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__5397\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29966\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__29966\,
            I => \N__29961\
        );

    \I__5395\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29958\
        );

    \I__5394\ : InMux
    port map (
            O => \N__29964\,
            I => \N__29955\
        );

    \I__5393\ : Odrv4
    port map (
            O => \N__29961\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__29958\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__29955\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__5390\ : CascadeMux
    port map (
            O => \N__29948\,
            I => \N__29945\
        );

    \I__5389\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29942\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__29942\,
            I => \N__29939\
        );

    \I__5387\ : Span4Mux_v
    port map (
            O => \N__29939\,
            I => \N__29936\
        );

    \I__5386\ : Odrv4
    port map (
            O => \N__29936\,
            I => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\
        );

    \I__5385\ : CascadeMux
    port map (
            O => \N__29933\,
            I => \N__29930\
        );

    \I__5384\ : InMux
    port map (
            O => \N__29930\,
            I => \N__29918\
        );

    \I__5383\ : InMux
    port map (
            O => \N__29929\,
            I => \N__29918\
        );

    \I__5382\ : InMux
    port map (
            O => \N__29928\,
            I => \N__29918\
        );

    \I__5381\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29918\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__29918\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5379\ : CascadeMux
    port map (
            O => \N__29915\,
            I => \N__29911\
        );

    \I__5378\ : InMux
    port map (
            O => \N__29914\,
            I => \N__29903\
        );

    \I__5377\ : InMux
    port map (
            O => \N__29911\,
            I => \N__29903\
        );

    \I__5376\ : InMux
    port map (
            O => \N__29910\,
            I => \N__29903\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__29903\,
            I => \N__29900\
        );

    \I__5374\ : Span4Mux_v
    port map (
            O => \N__29900\,
            I => \N__29897\
        );

    \I__5373\ : Span4Mux_h
    port map (
            O => \N__29897\,
            I => \N__29894\
        );

    \I__5372\ : Span4Mux_h
    port map (
            O => \N__29894\,
            I => \N__29891\
        );

    \I__5371\ : Odrv4
    port map (
            O => \N__29891\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__5370\ : CEMux
    port map (
            O => \N__29888\,
            I => \N__29883\
        );

    \I__5369\ : CEMux
    port map (
            O => \N__29887\,
            I => \N__29879\
        );

    \I__5368\ : CEMux
    port map (
            O => \N__29886\,
            I => \N__29876\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__29883\,
            I => \N__29872\
        );

    \I__5366\ : CEMux
    port map (
            O => \N__29882\,
            I => \N__29869\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__29879\,
            I => \N__29866\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__29876\,
            I => \N__29863\
        );

    \I__5363\ : CEMux
    port map (
            O => \N__29875\,
            I => \N__29860\
        );

    \I__5362\ : Span4Mux_h
    port map (
            O => \N__29872\,
            I => \N__29857\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__29869\,
            I => \N__29854\
        );

    \I__5360\ : Span4Mux_v
    port map (
            O => \N__29866\,
            I => \N__29847\
        );

    \I__5359\ : Span4Mux_v
    port map (
            O => \N__29863\,
            I => \N__29847\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__29860\,
            I => \N__29847\
        );

    \I__5357\ : Span4Mux_v
    port map (
            O => \N__29857\,
            I => \N__29844\
        );

    \I__5356\ : Span4Mux_v
    port map (
            O => \N__29854\,
            I => \N__29841\
        );

    \I__5355\ : Span4Mux_h
    port map (
            O => \N__29847\,
            I => \N__29838\
        );

    \I__5354\ : Span4Mux_v
    port map (
            O => \N__29844\,
            I => \N__29835\
        );

    \I__5353\ : Span4Mux_h
    port map (
            O => \N__29841\,
            I => \N__29830\
        );

    \I__5352\ : Span4Mux_h
    port map (
            O => \N__29838\,
            I => \N__29830\
        );

    \I__5351\ : Odrv4
    port map (
            O => \N__29835\,
            I => \delay_measurement_inst.delay_hc_timer.N_198_i\
        );

    \I__5350\ : Odrv4
    port map (
            O => \N__29830\,
            I => \delay_measurement_inst.delay_hc_timer.N_198_i\
        );

    \I__5349\ : CascadeMux
    port map (
            O => \N__29825\,
            I => \N__29822\
        );

    \I__5348\ : InMux
    port map (
            O => \N__29822\,
            I => \N__29819\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__29819\,
            I => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\
        );

    \I__5346\ : CascadeMux
    port map (
            O => \N__29816\,
            I => \N__29812\
        );

    \I__5345\ : CascadeMux
    port map (
            O => \N__29815\,
            I => \N__29809\
        );

    \I__5344\ : InMux
    port map (
            O => \N__29812\,
            I => \N__29806\
        );

    \I__5343\ : InMux
    port map (
            O => \N__29809\,
            I => \N__29803\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__29806\,
            I => \N__29799\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__29803\,
            I => \N__29796\
        );

    \I__5340\ : InMux
    port map (
            O => \N__29802\,
            I => \N__29793\
        );

    \I__5339\ : Span4Mux_v
    port map (
            O => \N__29799\,
            I => \N__29788\
        );

    \I__5338\ : Span4Mux_h
    port map (
            O => \N__29796\,
            I => \N__29788\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__29793\,
            I => \N__29785\
        );

    \I__5336\ : Span4Mux_h
    port map (
            O => \N__29788\,
            I => \N__29781\
        );

    \I__5335\ : Span4Mux_h
    port map (
            O => \N__29785\,
            I => \N__29778\
        );

    \I__5334\ : InMux
    port map (
            O => \N__29784\,
            I => \N__29775\
        );

    \I__5333\ : Odrv4
    port map (
            O => \N__29781\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__5332\ : Odrv4
    port map (
            O => \N__29778\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__29775\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__5330\ : InMux
    port map (
            O => \N__29768\,
            I => \N__29764\
        );

    \I__5329\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29761\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__29764\,
            I => \N__29757\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__29761\,
            I => \N__29754\
        );

    \I__5326\ : InMux
    port map (
            O => \N__29760\,
            I => \N__29751\
        );

    \I__5325\ : Odrv4
    port map (
            O => \N__29757\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__5324\ : Odrv4
    port map (
            O => \N__29754\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__29751\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__5322\ : InMux
    port map (
            O => \N__29744\,
            I => \N__29741\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__29741\,
            I => \N__29738\
        );

    \I__5320\ : Odrv12
    port map (
            O => \N__29738\,
            I => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\
        );

    \I__5319\ : CascadeMux
    port map (
            O => \N__29735\,
            I => \N__29732\
        );

    \I__5318\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29729\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__29729\,
            I => \N__29726\
        );

    \I__5316\ : Span4Mux_v
    port map (
            O => \N__29726\,
            I => \N__29723\
        );

    \I__5315\ : Odrv4
    port map (
            O => \N__29723\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__5314\ : CascadeMux
    port map (
            O => \N__29720\,
            I => \N__29716\
        );

    \I__5313\ : InMux
    port map (
            O => \N__29719\,
            I => \N__29713\
        );

    \I__5312\ : InMux
    port map (
            O => \N__29716\,
            I => \N__29710\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__29713\,
            I => \N__29706\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__29710\,
            I => \N__29703\
        );

    \I__5309\ : InMux
    port map (
            O => \N__29709\,
            I => \N__29700\
        );

    \I__5308\ : Odrv4
    port map (
            O => \N__29706\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__5307\ : Odrv4
    port map (
            O => \N__29703\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__29700\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__29693\,
            I => \N__29688\
        );

    \I__5304\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29685\
        );

    \I__5303\ : InMux
    port map (
            O => \N__29691\,
            I => \N__29682\
        );

    \I__5302\ : InMux
    port map (
            O => \N__29688\,
            I => \N__29679\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__29685\,
            I => \N__29676\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__29682\,
            I => \N__29672\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__29679\,
            I => \N__29669\
        );

    \I__5298\ : Span4Mux_v
    port map (
            O => \N__29676\,
            I => \N__29666\
        );

    \I__5297\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29663\
        );

    \I__5296\ : Span4Mux_v
    port map (
            O => \N__29672\,
            I => \N__29660\
        );

    \I__5295\ : Span4Mux_h
    port map (
            O => \N__29669\,
            I => \N__29653\
        );

    \I__5294\ : Span4Mux_h
    port map (
            O => \N__29666\,
            I => \N__29653\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__29663\,
            I => \N__29653\
        );

    \I__5292\ : Odrv4
    port map (
            O => \N__29660\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__5291\ : Odrv4
    port map (
            O => \N__29653\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__5290\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29645\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__29645\,
            I => \N__29642\
        );

    \I__5288\ : Span12Mux_v
    port map (
            O => \N__29642\,
            I => \N__29639\
        );

    \I__5287\ : Odrv12
    port map (
            O => \N__29639\,
            I => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\
        );

    \I__5286\ : CascadeMux
    port map (
            O => \N__29636\,
            I => \N__29632\
        );

    \I__5285\ : CascadeMux
    port map (
            O => \N__29635\,
            I => \N__29629\
        );

    \I__5284\ : InMux
    port map (
            O => \N__29632\,
            I => \N__29625\
        );

    \I__5283\ : InMux
    port map (
            O => \N__29629\,
            I => \N__29622\
        );

    \I__5282\ : InMux
    port map (
            O => \N__29628\,
            I => \N__29619\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__29625\,
            I => \N__29616\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__29622\,
            I => \N__29613\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__29619\,
            I => \N__29610\
        );

    \I__5278\ : Span4Mux_h
    port map (
            O => \N__29616\,
            I => \N__29607\
        );

    \I__5277\ : Span4Mux_h
    port map (
            O => \N__29613\,
            I => \N__29604\
        );

    \I__5276\ : Span4Mux_h
    port map (
            O => \N__29610\,
            I => \N__29601\
        );

    \I__5275\ : Span4Mux_v
    port map (
            O => \N__29607\,
            I => \N__29595\
        );

    \I__5274\ : Span4Mux_h
    port map (
            O => \N__29604\,
            I => \N__29595\
        );

    \I__5273\ : Span4Mux_v
    port map (
            O => \N__29601\,
            I => \N__29592\
        );

    \I__5272\ : InMux
    port map (
            O => \N__29600\,
            I => \N__29589\
        );

    \I__5271\ : Odrv4
    port map (
            O => \N__29595\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__5270\ : Odrv4
    port map (
            O => \N__29592\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__29589\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__5268\ : InMux
    port map (
            O => \N__29582\,
            I => \N__29579\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__29579\,
            I => \N__29576\
        );

    \I__5266\ : Span4Mux_h
    port map (
            O => \N__29576\,
            I => \N__29571\
        );

    \I__5265\ : InMux
    port map (
            O => \N__29575\,
            I => \N__29568\
        );

    \I__5264\ : InMux
    port map (
            O => \N__29574\,
            I => \N__29565\
        );

    \I__5263\ : Span4Mux_v
    port map (
            O => \N__29571\,
            I => \N__29560\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__29568\,
            I => \N__29560\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__29565\,
            I => \N__29557\
        );

    \I__5260\ : Odrv4
    port map (
            O => \N__29560\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__5259\ : Odrv4
    port map (
            O => \N__29557\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__5258\ : CascadeMux
    port map (
            O => \N__29552\,
            I => \N__29549\
        );

    \I__5257\ : InMux
    port map (
            O => \N__29549\,
            I => \N__29546\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__29546\,
            I => \N__29543\
        );

    \I__5255\ : Sp12to4
    port map (
            O => \N__29543\,
            I => \N__29540\
        );

    \I__5254\ : Odrv12
    port map (
            O => \N__29540\,
            I => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\
        );

    \I__5253\ : CascadeMux
    port map (
            O => \N__29537\,
            I => \N__29534\
        );

    \I__5252\ : InMux
    port map (
            O => \N__29534\,
            I => \N__29529\
        );

    \I__5251\ : InMux
    port map (
            O => \N__29533\,
            I => \N__29526\
        );

    \I__5250\ : InMux
    port map (
            O => \N__29532\,
            I => \N__29523\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__29529\,
            I => \N__29520\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__29526\,
            I => \N__29516\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__29523\,
            I => \N__29513\
        );

    \I__5246\ : Span4Mux_h
    port map (
            O => \N__29520\,
            I => \N__29510\
        );

    \I__5245\ : InMux
    port map (
            O => \N__29519\,
            I => \N__29507\
        );

    \I__5244\ : Span4Mux_h
    port map (
            O => \N__29516\,
            I => \N__29504\
        );

    \I__5243\ : Span4Mux_v
    port map (
            O => \N__29513\,
            I => \N__29501\
        );

    \I__5242\ : Span4Mux_h
    port map (
            O => \N__29510\,
            I => \N__29496\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__29507\,
            I => \N__29496\
        );

    \I__5240\ : Odrv4
    port map (
            O => \N__29504\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__29501\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__5238\ : Odrv4
    port map (
            O => \N__29496\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__5237\ : InMux
    port map (
            O => \N__29489\,
            I => \N__29485\
        );

    \I__5236\ : CascadeMux
    port map (
            O => \N__29488\,
            I => \N__29482\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__29485\,
            I => \N__29479\
        );

    \I__5234\ : InMux
    port map (
            O => \N__29482\,
            I => \N__29475\
        );

    \I__5233\ : Span4Mux_h
    port map (
            O => \N__29479\,
            I => \N__29472\
        );

    \I__5232\ : InMux
    port map (
            O => \N__29478\,
            I => \N__29469\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__29475\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__5230\ : Odrv4
    port map (
            O => \N__29472\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__29469\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__5228\ : CascadeMux
    port map (
            O => \N__29462\,
            I => \N__29459\
        );

    \I__5227\ : InMux
    port map (
            O => \N__29459\,
            I => \N__29456\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__29456\,
            I => \N__29453\
        );

    \I__5225\ : Span4Mux_h
    port map (
            O => \N__29453\,
            I => \N__29450\
        );

    \I__5224\ : Odrv4
    port map (
            O => \N__29450\,
            I => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\
        );

    \I__5223\ : CascadeMux
    port map (
            O => \N__29447\,
            I => \N__29443\
        );

    \I__5222\ : InMux
    port map (
            O => \N__29446\,
            I => \N__29440\
        );

    \I__5221\ : InMux
    port map (
            O => \N__29443\,
            I => \N__29437\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__29440\,
            I => \N__29434\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__29437\,
            I => \N__29431\
        );

    \I__5218\ : Span4Mux_v
    port map (
            O => \N__29434\,
            I => \N__29428\
        );

    \I__5217\ : Span4Mux_v
    port map (
            O => \N__29431\,
            I => \N__29425\
        );

    \I__5216\ : Odrv4
    port map (
            O => \N__29428\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__5215\ : Odrv4
    port map (
            O => \N__29425\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__5214\ : InMux
    port map (
            O => \N__29420\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__5213\ : InMux
    port map (
            O => \N__29417\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__5212\ : InMux
    port map (
            O => \N__29414\,
            I => \N__29411\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__29411\,
            I => \N__29408\
        );

    \I__5210\ : Span4Mux_h
    port map (
            O => \N__29408\,
            I => \N__29405\
        );

    \I__5209\ : Odrv4
    port map (
            O => \N__29405\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__5208\ : InMux
    port map (
            O => \N__29402\,
            I => \N__29399\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__29399\,
            I => \N__29396\
        );

    \I__5206\ : Odrv4
    port map (
            O => \N__29396\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__5205\ : InMux
    port map (
            O => \N__29393\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__5204\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29387\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__29387\,
            I => \N__29384\
        );

    \I__5202\ : Span4Mux_v
    port map (
            O => \N__29384\,
            I => \N__29381\
        );

    \I__5201\ : Odrv4
    port map (
            O => \N__29381\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__5200\ : InMux
    port map (
            O => \N__29378\,
            I => \N__29375\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__29375\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__5198\ : InMux
    port map (
            O => \N__29372\,
            I => \N__29369\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__29369\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__5196\ : InMux
    port map (
            O => \N__29366\,
            I => \N__29363\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__29363\,
            I => \N__29360\
        );

    \I__5194\ : Span4Mux_h
    port map (
            O => \N__29360\,
            I => \N__29357\
        );

    \I__5193\ : Odrv4
    port map (
            O => \N__29357\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__5192\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29351\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__29351\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__5190\ : InMux
    port map (
            O => \N__29348\,
            I => \N__29345\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__29345\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__5188\ : InMux
    port map (
            O => \N__29342\,
            I => \N__29339\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__29339\,
            I => \N__29336\
        );

    \I__5186\ : Span4Mux_h
    port map (
            O => \N__29336\,
            I => \N__29333\
        );

    \I__5185\ : Odrv4
    port map (
            O => \N__29333\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__5184\ : InMux
    port map (
            O => \N__29330\,
            I => \N__29327\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__29327\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__5182\ : InMux
    port map (
            O => \N__29324\,
            I => \N__29321\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__29321\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__5180\ : CascadeMux
    port map (
            O => \N__29318\,
            I => \N__29315\
        );

    \I__5179\ : InMux
    port map (
            O => \N__29315\,
            I => \N__29298\
        );

    \I__5178\ : InMux
    port map (
            O => \N__29314\,
            I => \N__29291\
        );

    \I__5177\ : InMux
    port map (
            O => \N__29313\,
            I => \N__29291\
        );

    \I__5176\ : InMux
    port map (
            O => \N__29312\,
            I => \N__29291\
        );

    \I__5175\ : InMux
    port map (
            O => \N__29311\,
            I => \N__29278\
        );

    \I__5174\ : InMux
    port map (
            O => \N__29310\,
            I => \N__29278\
        );

    \I__5173\ : InMux
    port map (
            O => \N__29309\,
            I => \N__29278\
        );

    \I__5172\ : InMux
    port map (
            O => \N__29308\,
            I => \N__29278\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29307\,
            I => \N__29278\
        );

    \I__5170\ : InMux
    port map (
            O => \N__29306\,
            I => \N__29278\
        );

    \I__5169\ : InMux
    port map (
            O => \N__29305\,
            I => \N__29271\
        );

    \I__5168\ : InMux
    port map (
            O => \N__29304\,
            I => \N__29271\
        );

    \I__5167\ : InMux
    port map (
            O => \N__29303\,
            I => \N__29271\
        );

    \I__5166\ : InMux
    port map (
            O => \N__29302\,
            I => \N__29266\
        );

    \I__5165\ : InMux
    port map (
            O => \N__29301\,
            I => \N__29266\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__29298\,
            I => \N__29263\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__29291\,
            I => \N__29260\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__29278\,
            I => \N__29257\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__29271\,
            I => \N__29252\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__29266\,
            I => \N__29252\
        );

    \I__5159\ : Span4Mux_h
    port map (
            O => \N__29263\,
            I => \N__29249\
        );

    \I__5158\ : Span4Mux_h
    port map (
            O => \N__29260\,
            I => \N__29246\
        );

    \I__5157\ : Span4Mux_v
    port map (
            O => \N__29257\,
            I => \N__29243\
        );

    \I__5156\ : Span4Mux_v
    port map (
            O => \N__29252\,
            I => \N__29240\
        );

    \I__5155\ : Odrv4
    port map (
            O => \N__29249\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__5154\ : Odrv4
    port map (
            O => \N__29246\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__29243\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__5152\ : Odrv4
    port map (
            O => \N__29240\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__5151\ : InMux
    port map (
            O => \N__29231\,
            I => \N__29228\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__29228\,
            I => \N__29225\
        );

    \I__5149\ : Span4Mux_v
    port map (
            O => \N__29225\,
            I => \N__29222\
        );

    \I__5148\ : Odrv4
    port map (
            O => \N__29222\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__5147\ : CEMux
    port map (
            O => \N__29219\,
            I => \N__29214\
        );

    \I__5146\ : CEMux
    port map (
            O => \N__29218\,
            I => \N__29211\
        );

    \I__5145\ : CEMux
    port map (
            O => \N__29217\,
            I => \N__29207\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__29214\,
            I => \N__29204\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__29211\,
            I => \N__29201\
        );

    \I__5142\ : CEMux
    port map (
            O => \N__29210\,
            I => \N__29198\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__29207\,
            I => \N__29195\
        );

    \I__5140\ : Span4Mux_v
    port map (
            O => \N__29204\,
            I => \N__29192\
        );

    \I__5139\ : Span4Mux_v
    port map (
            O => \N__29201\,
            I => \N__29189\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__29198\,
            I => \N__29186\
        );

    \I__5137\ : Span4Mux_h
    port map (
            O => \N__29195\,
            I => \N__29183\
        );

    \I__5136\ : Span4Mux_h
    port map (
            O => \N__29192\,
            I => \N__29180\
        );

    \I__5135\ : Span4Mux_h
    port map (
            O => \N__29189\,
            I => \N__29177\
        );

    \I__5134\ : Span4Mux_h
    port map (
            O => \N__29186\,
            I => \N__29174\
        );

    \I__5133\ : Span4Mux_v
    port map (
            O => \N__29183\,
            I => \N__29171\
        );

    \I__5132\ : Span4Mux_v
    port map (
            O => \N__29180\,
            I => \N__29164\
        );

    \I__5131\ : Span4Mux_v
    port map (
            O => \N__29177\,
            I => \N__29164\
        );

    \I__5130\ : Span4Mux_v
    port map (
            O => \N__29174\,
            I => \N__29164\
        );

    \I__5129\ : Odrv4
    port map (
            O => \N__29171\,
            I => \delay_measurement_inst.delay_hc_timer.N_199_i\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__29164\,
            I => \delay_measurement_inst.delay_hc_timer.N_199_i\
        );

    \I__5127\ : InMux
    port map (
            O => \N__29159\,
            I => \N__29153\
        );

    \I__5126\ : InMux
    port map (
            O => \N__29158\,
            I => \N__29153\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__29153\,
            I => \N__29150\
        );

    \I__5124\ : Span4Mux_h
    port map (
            O => \N__29150\,
            I => \N__29147\
        );

    \I__5123\ : Span4Mux_h
    port map (
            O => \N__29147\,
            I => \N__29144\
        );

    \I__5122\ : Span4Mux_h
    port map (
            O => \N__29144\,
            I => \N__29139\
        );

    \I__5121\ : InMux
    port map (
            O => \N__29143\,
            I => \N__29136\
        );

    \I__5120\ : InMux
    port map (
            O => \N__29142\,
            I => \N__29133\
        );

    \I__5119\ : Span4Mux_v
    port map (
            O => \N__29139\,
            I => \N__29130\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__29136\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__29133\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__29130\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__5115\ : InMux
    port map (
            O => \N__29123\,
            I => \N__29091\
        );

    \I__5114\ : InMux
    port map (
            O => \N__29122\,
            I => \N__29091\
        );

    \I__5113\ : InMux
    port map (
            O => \N__29121\,
            I => \N__29091\
        );

    \I__5112\ : InMux
    port map (
            O => \N__29120\,
            I => \N__29091\
        );

    \I__5111\ : InMux
    port map (
            O => \N__29119\,
            I => \N__29082\
        );

    \I__5110\ : InMux
    port map (
            O => \N__29118\,
            I => \N__29082\
        );

    \I__5109\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29082\
        );

    \I__5108\ : InMux
    port map (
            O => \N__29116\,
            I => \N__29082\
        );

    \I__5107\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29073\
        );

    \I__5106\ : InMux
    port map (
            O => \N__29114\,
            I => \N__29073\
        );

    \I__5105\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29073\
        );

    \I__5104\ : InMux
    port map (
            O => \N__29112\,
            I => \N__29073\
        );

    \I__5103\ : InMux
    port map (
            O => \N__29111\,
            I => \N__29064\
        );

    \I__5102\ : InMux
    port map (
            O => \N__29110\,
            I => \N__29064\
        );

    \I__5101\ : InMux
    port map (
            O => \N__29109\,
            I => \N__29064\
        );

    \I__5100\ : InMux
    port map (
            O => \N__29108\,
            I => \N__29064\
        );

    \I__5099\ : InMux
    port map (
            O => \N__29107\,
            I => \N__29049\
        );

    \I__5098\ : InMux
    port map (
            O => \N__29106\,
            I => \N__29049\
        );

    \I__5097\ : InMux
    port map (
            O => \N__29105\,
            I => \N__29049\
        );

    \I__5096\ : InMux
    port map (
            O => \N__29104\,
            I => \N__29049\
        );

    \I__5095\ : InMux
    port map (
            O => \N__29103\,
            I => \N__29040\
        );

    \I__5094\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29040\
        );

    \I__5093\ : InMux
    port map (
            O => \N__29101\,
            I => \N__29040\
        );

    \I__5092\ : InMux
    port map (
            O => \N__29100\,
            I => \N__29040\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__29091\,
            I => \N__29031\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__29082\,
            I => \N__29031\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__29073\,
            I => \N__29031\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__29064\,
            I => \N__29031\
        );

    \I__5087\ : InMux
    port map (
            O => \N__29063\,
            I => \N__29026\
        );

    \I__5086\ : InMux
    port map (
            O => \N__29062\,
            I => \N__29026\
        );

    \I__5085\ : InMux
    port map (
            O => \N__29061\,
            I => \N__29017\
        );

    \I__5084\ : InMux
    port map (
            O => \N__29060\,
            I => \N__29017\
        );

    \I__5083\ : InMux
    port map (
            O => \N__29059\,
            I => \N__29017\
        );

    \I__5082\ : InMux
    port map (
            O => \N__29058\,
            I => \N__29017\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__29049\,
            I => \N__29010\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__29040\,
            I => \N__29010\
        );

    \I__5079\ : Span4Mux_v
    port map (
            O => \N__29031\,
            I => \N__29010\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__29026\,
            I => \N__29005\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__29017\,
            I => \N__29005\
        );

    \I__5076\ : Span4Mux_h
    port map (
            O => \N__29010\,
            I => \N__29002\
        );

    \I__5075\ : Span12Mux_h
    port map (
            O => \N__29005\,
            I => \N__28999\
        );

    \I__5074\ : Span4Mux_v
    port map (
            O => \N__29002\,
            I => \N__28996\
        );

    \I__5073\ : Odrv12
    port map (
            O => \N__28999\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5072\ : Odrv4
    port map (
            O => \N__28996\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5071\ : InMux
    port map (
            O => \N__28991\,
            I => \N__28988\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__28988\,
            I => \N__28985\
        );

    \I__5069\ : Span4Mux_h
    port map (
            O => \N__28985\,
            I => \N__28982\
        );

    \I__5068\ : Odrv4
    port map (
            O => \N__28982\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__5067\ : InMux
    port map (
            O => \N__28979\,
            I => \N__28976\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__28976\,
            I => \N__28973\
        );

    \I__5065\ : Odrv4
    port map (
            O => \N__28973\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__5064\ : InMux
    port map (
            O => \N__28970\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__5063\ : InMux
    port map (
            O => \N__28967\,
            I => \N__28964\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__28964\,
            I => \N__28961\
        );

    \I__5061\ : Odrv12
    port map (
            O => \N__28961\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__5060\ : InMux
    port map (
            O => \N__28958\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__5059\ : InMux
    port map (
            O => \N__28955\,
            I => \N__28952\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__28952\,
            I => \N__28949\
        );

    \I__5057\ : Odrv4
    port map (
            O => \N__28949\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__5056\ : InMux
    port map (
            O => \N__28946\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__5055\ : CascadeMux
    port map (
            O => \N__28943\,
            I => \N__28940\
        );

    \I__5054\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28937\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__28937\,
            I => \N__28934\
        );

    \I__5052\ : Span4Mux_v
    port map (
            O => \N__28934\,
            I => \N__28931\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__28931\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__5050\ : InMux
    port map (
            O => \N__28928\,
            I => \N__28925\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__28925\,
            I => \N__28922\
        );

    \I__5048\ : Span4Mux_v
    port map (
            O => \N__28922\,
            I => \N__28919\
        );

    \I__5047\ : Span4Mux_h
    port map (
            O => \N__28919\,
            I => \N__28916\
        );

    \I__5046\ : Odrv4
    port map (
            O => \N__28916\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__5045\ : InMux
    port map (
            O => \N__28913\,
            I => \bfn_12_16_0_\
        );

    \I__5044\ : InMux
    port map (
            O => \N__28910\,
            I => \N__28907\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__28907\,
            I => \N__28904\
        );

    \I__5042\ : Span4Mux_v
    port map (
            O => \N__28904\,
            I => \N__28901\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__28901\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__5040\ : InMux
    port map (
            O => \N__28898\,
            I => \N__28895\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__28895\,
            I => \N__28892\
        );

    \I__5038\ : Span4Mux_v
    port map (
            O => \N__28892\,
            I => \N__28889\
        );

    \I__5037\ : Span4Mux_h
    port map (
            O => \N__28889\,
            I => \N__28886\
        );

    \I__5036\ : Odrv4
    port map (
            O => \N__28886\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__5035\ : InMux
    port map (
            O => \N__28883\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__5034\ : CascadeMux
    port map (
            O => \N__28880\,
            I => \N__28877\
        );

    \I__5033\ : InMux
    port map (
            O => \N__28877\,
            I => \N__28874\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__28874\,
            I => \N__28871\
        );

    \I__5031\ : Span4Mux_v
    port map (
            O => \N__28871\,
            I => \N__28868\
        );

    \I__5030\ : Odrv4
    port map (
            O => \N__28868\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__5029\ : InMux
    port map (
            O => \N__28865\,
            I => \N__28862\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__28862\,
            I => \N__28859\
        );

    \I__5027\ : Span4Mux_h
    port map (
            O => \N__28859\,
            I => \N__28856\
        );

    \I__5026\ : Odrv4
    port map (
            O => \N__28856\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__5025\ : InMux
    port map (
            O => \N__28853\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__5024\ : InMux
    port map (
            O => \N__28850\,
            I => \N__28847\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__28847\,
            I => \N__28844\
        );

    \I__5022\ : Span4Mux_v
    port map (
            O => \N__28844\,
            I => \N__28841\
        );

    \I__5021\ : Odrv4
    port map (
            O => \N__28841\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__5020\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28835\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__28835\,
            I => \N__28832\
        );

    \I__5018\ : Span4Mux_h
    port map (
            O => \N__28832\,
            I => \N__28829\
        );

    \I__5017\ : Odrv4
    port map (
            O => \N__28829\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__5016\ : InMux
    port map (
            O => \N__28826\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__5015\ : CascadeMux
    port map (
            O => \N__28823\,
            I => \N__28820\
        );

    \I__5014\ : InMux
    port map (
            O => \N__28820\,
            I => \N__28817\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__28817\,
            I => \N__28814\
        );

    \I__5012\ : Span4Mux_v
    port map (
            O => \N__28814\,
            I => \N__28811\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__28811\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__5010\ : InMux
    port map (
            O => \N__28808\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__5009\ : InMux
    port map (
            O => \N__28805\,
            I => \N__28802\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__28802\,
            I => \N__28799\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__28799\,
            I => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\
        );

    \I__5006\ : InMux
    port map (
            O => \N__28796\,
            I => \N__28793\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__28793\,
            I => \N__28790\
        );

    \I__5004\ : Odrv4
    port map (
            O => \N__28790\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__5003\ : InMux
    port map (
            O => \N__28787\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__5002\ : InMux
    port map (
            O => \N__28784\,
            I => \N__28781\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__28781\,
            I => \N__28778\
        );

    \I__5000\ : Span4Mux_h
    port map (
            O => \N__28778\,
            I => \N__28775\
        );

    \I__4999\ : Odrv4
    port map (
            O => \N__28775\,
            I => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\
        );

    \I__4998\ : CascadeMux
    port map (
            O => \N__28772\,
            I => \N__28769\
        );

    \I__4997\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28766\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__28766\,
            I => \N__28763\
        );

    \I__4995\ : Span4Mux_v
    port map (
            O => \N__28763\,
            I => \N__28760\
        );

    \I__4994\ : Span4Mux_h
    port map (
            O => \N__28760\,
            I => \N__28757\
        );

    \I__4993\ : Odrv4
    port map (
            O => \N__28757\,
            I => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\
        );

    \I__4992\ : InMux
    port map (
            O => \N__28754\,
            I => \N__28751\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__28751\,
            I => \N__28748\
        );

    \I__4990\ : Odrv4
    port map (
            O => \N__28748\,
            I => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\
        );

    \I__4989\ : InMux
    port map (
            O => \N__28745\,
            I => \N__28740\
        );

    \I__4988\ : InMux
    port map (
            O => \N__28744\,
            I => \N__28736\
        );

    \I__4987\ : InMux
    port map (
            O => \N__28743\,
            I => \N__28733\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__28740\,
            I => \N__28730\
        );

    \I__4985\ : CascadeMux
    port map (
            O => \N__28739\,
            I => \N__28727\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__28736\,
            I => \N__28724\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__28733\,
            I => \N__28721\
        );

    \I__4982\ : Span4Mux_h
    port map (
            O => \N__28730\,
            I => \N__28718\
        );

    \I__4981\ : InMux
    port map (
            O => \N__28727\,
            I => \N__28715\
        );

    \I__4980\ : Odrv4
    port map (
            O => \N__28724\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__4979\ : Odrv12
    port map (
            O => \N__28721\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__4978\ : Odrv4
    port map (
            O => \N__28718\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__28715\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__4976\ : InMux
    port map (
            O => \N__28706\,
            I => \N__28702\
        );

    \I__4975\ : InMux
    port map (
            O => \N__28705\,
            I => \N__28698\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__28702\,
            I => \N__28695\
        );

    \I__4973\ : InMux
    port map (
            O => \N__28701\,
            I => \N__28692\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__28698\,
            I => \N__28689\
        );

    \I__4971\ : Span4Mux_h
    port map (
            O => \N__28695\,
            I => \N__28686\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__28692\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__4969\ : Odrv4
    port map (
            O => \N__28689\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__4968\ : Odrv4
    port map (
            O => \N__28686\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__4967\ : CascadeMux
    port map (
            O => \N__28679\,
            I => \N__28676\
        );

    \I__4966\ : InMux
    port map (
            O => \N__28676\,
            I => \N__28673\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__28673\,
            I => \N__28670\
        );

    \I__4964\ : Odrv4
    port map (
            O => \N__28670\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__4963\ : InMux
    port map (
            O => \N__28667\,
            I => \N__28663\
        );

    \I__4962\ : InMux
    port map (
            O => \N__28666\,
            I => \N__28659\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__28663\,
            I => \N__28656\
        );

    \I__4960\ : InMux
    port map (
            O => \N__28662\,
            I => \N__28653\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__28659\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__4958\ : Odrv4
    port map (
            O => \N__28656\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__28653\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__4956\ : InMux
    port map (
            O => \N__28646\,
            I => \N__28642\
        );

    \I__4955\ : InMux
    port map (
            O => \N__28645\,
            I => \N__28637\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__28642\,
            I => \N__28634\
        );

    \I__4953\ : InMux
    port map (
            O => \N__28641\,
            I => \N__28631\
        );

    \I__4952\ : InMux
    port map (
            O => \N__28640\,
            I => \N__28628\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__28637\,
            I => \N__28625\
        );

    \I__4950\ : Span4Mux_v
    port map (
            O => \N__28634\,
            I => \N__28620\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__28631\,
            I => \N__28620\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__28628\,
            I => \N__28617\
        );

    \I__4947\ : Span12Mux_v
    port map (
            O => \N__28625\,
            I => \N__28614\
        );

    \I__4946\ : Span4Mux_h
    port map (
            O => \N__28620\,
            I => \N__28609\
        );

    \I__4945\ : Span4Mux_v
    port map (
            O => \N__28617\,
            I => \N__28609\
        );

    \I__4944\ : Odrv12
    port map (
            O => \N__28614\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__4943\ : Odrv4
    port map (
            O => \N__28609\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__4942\ : CascadeMux
    port map (
            O => \N__28604\,
            I => \N__28601\
        );

    \I__4941\ : InMux
    port map (
            O => \N__28601\,
            I => \N__28595\
        );

    \I__4940\ : InMux
    port map (
            O => \N__28600\,
            I => \N__28595\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__28595\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\
        );

    \I__4938\ : InMux
    port map (
            O => \N__28592\,
            I => \N__28588\
        );

    \I__4937\ : InMux
    port map (
            O => \N__28591\,
            I => \N__28585\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__28588\,
            I => \N__28581\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__28585\,
            I => \N__28578\
        );

    \I__4934\ : InMux
    port map (
            O => \N__28584\,
            I => \N__28574\
        );

    \I__4933\ : Span4Mux_h
    port map (
            O => \N__28581\,
            I => \N__28571\
        );

    \I__4932\ : Span4Mux_v
    port map (
            O => \N__28578\,
            I => \N__28568\
        );

    \I__4931\ : InMux
    port map (
            O => \N__28577\,
            I => \N__28565\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__28574\,
            I => \N__28562\
        );

    \I__4929\ : Span4Mux_v
    port map (
            O => \N__28571\,
            I => \N__28559\
        );

    \I__4928\ : Span4Mux_h
    port map (
            O => \N__28568\,
            I => \N__28554\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__28565\,
            I => \N__28554\
        );

    \I__4926\ : Span4Mux_h
    port map (
            O => \N__28562\,
            I => \N__28551\
        );

    \I__4925\ : Span4Mux_v
    port map (
            O => \N__28559\,
            I => \N__28548\
        );

    \I__4924\ : Span4Mux_v
    port map (
            O => \N__28554\,
            I => \N__28545\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__28551\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__4922\ : Odrv4
    port map (
            O => \N__28548\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__28545\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__4920\ : InMux
    port map (
            O => \N__28538\,
            I => \N__28535\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__28535\,
            I => \N__28531\
        );

    \I__4918\ : InMux
    port map (
            O => \N__28534\,
            I => \N__28527\
        );

    \I__4917\ : Span4Mux_v
    port map (
            O => \N__28531\,
            I => \N__28524\
        );

    \I__4916\ : InMux
    port map (
            O => \N__28530\,
            I => \N__28521\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__28527\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__4914\ : Odrv4
    port map (
            O => \N__28524\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__28521\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__4912\ : CEMux
    port map (
            O => \N__28514\,
            I => \N__28475\
        );

    \I__4911\ : CEMux
    port map (
            O => \N__28513\,
            I => \N__28475\
        );

    \I__4910\ : CEMux
    port map (
            O => \N__28512\,
            I => \N__28475\
        );

    \I__4909\ : CEMux
    port map (
            O => \N__28511\,
            I => \N__28475\
        );

    \I__4908\ : CEMux
    port map (
            O => \N__28510\,
            I => \N__28475\
        );

    \I__4907\ : CEMux
    port map (
            O => \N__28509\,
            I => \N__28475\
        );

    \I__4906\ : CEMux
    port map (
            O => \N__28508\,
            I => \N__28475\
        );

    \I__4905\ : CEMux
    port map (
            O => \N__28507\,
            I => \N__28475\
        );

    \I__4904\ : CEMux
    port map (
            O => \N__28506\,
            I => \N__28475\
        );

    \I__4903\ : CEMux
    port map (
            O => \N__28505\,
            I => \N__28475\
        );

    \I__4902\ : CEMux
    port map (
            O => \N__28504\,
            I => \N__28475\
        );

    \I__4901\ : CEMux
    port map (
            O => \N__28503\,
            I => \N__28475\
        );

    \I__4900\ : CEMux
    port map (
            O => \N__28502\,
            I => \N__28475\
        );

    \I__4899\ : GlobalMux
    port map (
            O => \N__28475\,
            I => \N__28472\
        );

    \I__4898\ : gio2CtrlBuf
    port map (
            O => \N__28472\,
            I => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \I__4897\ : InMux
    port map (
            O => \N__28469\,
            I => \N__28466\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__28466\,
            I => \N__28463\
        );

    \I__4895\ : Span4Mux_h
    port map (
            O => \N__28463\,
            I => \N__28459\
        );

    \I__4894\ : InMux
    port map (
            O => \N__28462\,
            I => \N__28456\
        );

    \I__4893\ : Odrv4
    port map (
            O => \N__28459\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__28456\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\
        );

    \I__4891\ : InMux
    port map (
            O => \N__28451\,
            I => \N__28446\
        );

    \I__4890\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28443\
        );

    \I__4889\ : InMux
    port map (
            O => \N__28449\,
            I => \N__28440\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__28446\,
            I => \N__28437\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__28443\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__28440\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__4885\ : Odrv4
    port map (
            O => \N__28437\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__28430\,
            I => \N__28427\
        );

    \I__4883\ : InMux
    port map (
            O => \N__28427\,
            I => \N__28423\
        );

    \I__4882\ : CascadeMux
    port map (
            O => \N__28426\,
            I => \N__28419\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__28423\,
            I => \N__28416\
        );

    \I__4880\ : InMux
    port map (
            O => \N__28422\,
            I => \N__28413\
        );

    \I__4879\ : InMux
    port map (
            O => \N__28419\,
            I => \N__28410\
        );

    \I__4878\ : Span4Mux_h
    port map (
            O => \N__28416\,
            I => \N__28407\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__28413\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__28410\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__4875\ : Odrv4
    port map (
            O => \N__28407\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__4874\ : InMux
    port map (
            O => \N__28400\,
            I => \N__28397\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__28397\,
            I => \N__28394\
        );

    \I__4872\ : Span4Mux_v
    port map (
            O => \N__28394\,
            I => \N__28390\
        );

    \I__4871\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28387\
        );

    \I__4870\ : Odrv4
    port map (
            O => \N__28390\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__28387\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\
        );

    \I__4868\ : CascadeMux
    port map (
            O => \N__28382\,
            I => \N__28379\
        );

    \I__4867\ : InMux
    port map (
            O => \N__28379\,
            I => \N__28376\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__28376\,
            I => \N__28373\
        );

    \I__4865\ : Span4Mux_h
    port map (
            O => \N__28373\,
            I => \N__28370\
        );

    \I__4864\ : Odrv4
    port map (
            O => \N__28370\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\
        );

    \I__4863\ : InMux
    port map (
            O => \N__28367\,
            I => \N__28363\
        );

    \I__4862\ : InMux
    port map (
            O => \N__28366\,
            I => \N__28360\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__28363\,
            I => \N__28357\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__28360\,
            I => \N__28354\
        );

    \I__4859\ : Span4Mux_h
    port map (
            O => \N__28357\,
            I => \N__28351\
        );

    \I__4858\ : Span4Mux_v
    port map (
            O => \N__28354\,
            I => \N__28348\
        );

    \I__4857\ : Odrv4
    port map (
            O => \N__28351\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__4856\ : Odrv4
    port map (
            O => \N__28348\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__4855\ : CascadeMux
    port map (
            O => \N__28343\,
            I => \N__28340\
        );

    \I__4854\ : InMux
    port map (
            O => \N__28340\,
            I => \N__28337\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__28337\,
            I => \N__28334\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__28334\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\
        );

    \I__4851\ : CascadeMux
    port map (
            O => \N__28331\,
            I => \N__28327\
        );

    \I__4850\ : InMux
    port map (
            O => \N__28330\,
            I => \N__28321\
        );

    \I__4849\ : InMux
    port map (
            O => \N__28327\,
            I => \N__28321\
        );

    \I__4848\ : InMux
    port map (
            O => \N__28326\,
            I => \N__28318\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__28321\,
            I => \N__28314\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__28318\,
            I => \N__28311\
        );

    \I__4845\ : InMux
    port map (
            O => \N__28317\,
            I => \N__28308\
        );

    \I__4844\ : Odrv4
    port map (
            O => \N__28314\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__4843\ : Odrv4
    port map (
            O => \N__28311\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__28308\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__4841\ : InMux
    port map (
            O => \N__28301\,
            I => \N__28298\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__28298\,
            I => \N__28294\
        );

    \I__4839\ : InMux
    port map (
            O => \N__28297\,
            I => \N__28291\
        );

    \I__4838\ : Span4Mux_h
    port map (
            O => \N__28294\,
            I => \N__28288\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__28291\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__28288\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__4835\ : InMux
    port map (
            O => \N__28283\,
            I => \N__28280\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__28280\,
            I => \N__28274\
        );

    \I__4833\ : InMux
    port map (
            O => \N__28279\,
            I => \N__28267\
        );

    \I__4832\ : InMux
    port map (
            O => \N__28278\,
            I => \N__28267\
        );

    \I__4831\ : InMux
    port map (
            O => \N__28277\,
            I => \N__28267\
        );

    \I__4830\ : Odrv12
    port map (
            O => \N__28274\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__28267\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__4828\ : CascadeMux
    port map (
            O => \N__28262\,
            I => \N__28258\
        );

    \I__4827\ : InMux
    port map (
            O => \N__28261\,
            I => \N__28247\
        );

    \I__4826\ : InMux
    port map (
            O => \N__28258\,
            I => \N__28247\
        );

    \I__4825\ : InMux
    port map (
            O => \N__28257\,
            I => \N__28247\
        );

    \I__4824\ : InMux
    port map (
            O => \N__28256\,
            I => \N__28247\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__28247\,
            I => \N__28244\
        );

    \I__4822\ : Span4Mux_h
    port map (
            O => \N__28244\,
            I => \N__28241\
        );

    \I__4821\ : Odrv4
    port map (
            O => \N__28241\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__4820\ : InMux
    port map (
            O => \N__28238\,
            I => \N__28234\
        );

    \I__4819\ : InMux
    port map (
            O => \N__28237\,
            I => \N__28231\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__28234\,
            I => \N__28228\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__28231\,
            I => \N__28225\
        );

    \I__4816\ : Span4Mux_h
    port map (
            O => \N__28228\,
            I => \N__28222\
        );

    \I__4815\ : Span4Mux_h
    port map (
            O => \N__28225\,
            I => \N__28219\
        );

    \I__4814\ : Odrv4
    port map (
            O => \N__28222\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__4813\ : Odrv4
    port map (
            O => \N__28219\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__4812\ : CascadeMux
    port map (
            O => \N__28214\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\
        );

    \I__4811\ : InMux
    port map (
            O => \N__28211\,
            I => \N__28204\
        );

    \I__4810\ : InMux
    port map (
            O => \N__28210\,
            I => \N__28204\
        );

    \I__4809\ : InMux
    port map (
            O => \N__28209\,
            I => \N__28201\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__28204\,
            I => \N__28198\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__28201\,
            I => \N__28193\
        );

    \I__4806\ : Span4Mux_v
    port map (
            O => \N__28198\,
            I => \N__28190\
        );

    \I__4805\ : InMux
    port map (
            O => \N__28197\,
            I => \N__28185\
        );

    \I__4804\ : InMux
    port map (
            O => \N__28196\,
            I => \N__28185\
        );

    \I__4803\ : Odrv12
    port map (
            O => \N__28193\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__4802\ : Odrv4
    port map (
            O => \N__28190\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__28185\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__4800\ : InMux
    port map (
            O => \N__28178\,
            I => \N__28175\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__28175\,
            I => \N__28170\
        );

    \I__4798\ : InMux
    port map (
            O => \N__28174\,
            I => \N__28167\
        );

    \I__4797\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28163\
        );

    \I__4796\ : Span4Mux_v
    port map (
            O => \N__28170\,
            I => \N__28158\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__28167\,
            I => \N__28158\
        );

    \I__4794\ : InMux
    port map (
            O => \N__28166\,
            I => \N__28155\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__28163\,
            I => \N__28152\
        );

    \I__4792\ : Span4Mux_h
    port map (
            O => \N__28158\,
            I => \N__28149\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__28155\,
            I => \N__28146\
        );

    \I__4790\ : Span4Mux_v
    port map (
            O => \N__28152\,
            I => \N__28143\
        );

    \I__4789\ : Span4Mux_v
    port map (
            O => \N__28149\,
            I => \N__28140\
        );

    \I__4788\ : Span4Mux_v
    port map (
            O => \N__28146\,
            I => \N__28137\
        );

    \I__4787\ : Odrv4
    port map (
            O => \N__28143\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__4786\ : Odrv4
    port map (
            O => \N__28140\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__28137\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__4784\ : InMux
    port map (
            O => \N__28130\,
            I => \N__28127\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__28127\,
            I => \N__28122\
        );

    \I__4782\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28119\
        );

    \I__4781\ : InMux
    port map (
            O => \N__28125\,
            I => \N__28116\
        );

    \I__4780\ : Span4Mux_v
    port map (
            O => \N__28122\,
            I => \N__28113\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__28119\,
            I => \N__28110\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__28116\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__4777\ : Odrv4
    port map (
            O => \N__28113\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__28110\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__4775\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28100\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__28100\,
            I => \N__28097\
        );

    \I__4773\ : Span4Mux_v
    port map (
            O => \N__28097\,
            I => \N__28094\
        );

    \I__4772\ : Odrv4
    port map (
            O => \N__28094\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\
        );

    \I__4771\ : InMux
    port map (
            O => \N__28091\,
            I => \N__28084\
        );

    \I__4770\ : InMux
    port map (
            O => \N__28090\,
            I => \N__28084\
        );

    \I__4769\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28081\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__28084\,
            I => \N__28078\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__28081\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__4766\ : Odrv4
    port map (
            O => \N__28078\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__28073\,
            I => \N__28070\
        );

    \I__4764\ : InMux
    port map (
            O => \N__28070\,
            I => \N__28064\
        );

    \I__4763\ : InMux
    port map (
            O => \N__28069\,
            I => \N__28064\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__28064\,
            I => \N__28061\
        );

    \I__4761\ : Span4Mux_h
    port map (
            O => \N__28061\,
            I => \N__28058\
        );

    \I__4760\ : Span4Mux_h
    port map (
            O => \N__28058\,
            I => \N__28055\
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__28055\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\
        );

    \I__4758\ : CascadeMux
    port map (
            O => \N__28052\,
            I => \N__28048\
        );

    \I__4757\ : InMux
    port map (
            O => \N__28051\,
            I => \N__28043\
        );

    \I__4756\ : InMux
    port map (
            O => \N__28048\,
            I => \N__28043\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__28043\,
            I => \N__28039\
        );

    \I__4754\ : InMux
    port map (
            O => \N__28042\,
            I => \N__28036\
        );

    \I__4753\ : Span4Mux_h
    port map (
            O => \N__28039\,
            I => \N__28033\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__28036\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__4751\ : Odrv4
    port map (
            O => \N__28033\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__4750\ : InMux
    port map (
            O => \N__28028\,
            I => \N__28022\
        );

    \I__4749\ : InMux
    port map (
            O => \N__28027\,
            I => \N__28022\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__28022\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__28019\,
            I => \N__28016\
        );

    \I__4746\ : InMux
    port map (
            O => \N__28016\,
            I => \N__28013\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__28013\,
            I => \N__28010\
        );

    \I__4744\ : Span4Mux_h
    port map (
            O => \N__28010\,
            I => \N__28007\
        );

    \I__4743\ : Odrv4
    port map (
            O => \N__28007\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt28\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__28004\,
            I => \N__28001\
        );

    \I__4741\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27998\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__27998\,
            I => \N__27995\
        );

    \I__4739\ : Span4Mux_h
    port map (
            O => \N__27995\,
            I => \N__27992\
        );

    \I__4738\ : Odrv4
    port map (
            O => \N__27992\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt24\
        );

    \I__4737\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27984\
        );

    \I__4736\ : InMux
    port map (
            O => \N__27988\,
            I => \N__27979\
        );

    \I__4735\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27979\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__27984\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__27979\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__27974\,
            I => \N__27971\
        );

    \I__4731\ : InMux
    port map (
            O => \N__27971\,
            I => \N__27964\
        );

    \I__4730\ : InMux
    port map (
            O => \N__27970\,
            I => \N__27964\
        );

    \I__4729\ : InMux
    port map (
            O => \N__27969\,
            I => \N__27961\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__27964\,
            I => \N__27958\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__27961\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__4726\ : Odrv4
    port map (
            O => \N__27958\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__4725\ : InMux
    port map (
            O => \N__27953\,
            I => \N__27950\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__27950\,
            I => \N__27947\
        );

    \I__4723\ : Span4Mux_h
    port map (
            O => \N__27947\,
            I => \N__27944\
        );

    \I__4722\ : Odrv4
    port map (
            O => \N__27944\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\
        );

    \I__4721\ : InMux
    port map (
            O => \N__27941\,
            I => \N__27935\
        );

    \I__4720\ : InMux
    port map (
            O => \N__27940\,
            I => \N__27935\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__27935\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\
        );

    \I__4718\ : CascadeMux
    port map (
            O => \N__27932\,
            I => \N__27928\
        );

    \I__4717\ : InMux
    port map (
            O => \N__27931\,
            I => \N__27923\
        );

    \I__4716\ : InMux
    port map (
            O => \N__27928\,
            I => \N__27923\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__27923\,
            I => \N__27919\
        );

    \I__4714\ : InMux
    port map (
            O => \N__27922\,
            I => \N__27916\
        );

    \I__4713\ : Span4Mux_h
    port map (
            O => \N__27919\,
            I => \N__27913\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__27916\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__27913\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__4710\ : InMux
    port map (
            O => \N__27908\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__4709\ : InMux
    port map (
            O => \N__27905\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__4708\ : InMux
    port map (
            O => \N__27902\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__4707\ : InMux
    port map (
            O => \N__27899\,
            I => \N__27889\
        );

    \I__4706\ : InMux
    port map (
            O => \N__27898\,
            I => \N__27889\
        );

    \I__4705\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27889\
        );

    \I__4704\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27886\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__27889\,
            I => \N__27883\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__27886\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__4701\ : Odrv4
    port map (
            O => \N__27883\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__4700\ : InMux
    port map (
            O => \N__27878\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__4699\ : InMux
    port map (
            O => \N__27875\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__4698\ : CascadeMux
    port map (
            O => \N__27872\,
            I => \N__27867\
        );

    \I__4697\ : CascadeMux
    port map (
            O => \N__27871\,
            I => \N__27864\
        );

    \I__4696\ : InMux
    port map (
            O => \N__27870\,
            I => \N__27857\
        );

    \I__4695\ : InMux
    port map (
            O => \N__27867\,
            I => \N__27857\
        );

    \I__4694\ : InMux
    port map (
            O => \N__27864\,
            I => \N__27857\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__27857\,
            I => \N__27853\
        );

    \I__4692\ : InMux
    port map (
            O => \N__27856\,
            I => \N__27850\
        );

    \I__4691\ : Span4Mux_h
    port map (
            O => \N__27853\,
            I => \N__27847\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__27850\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__4689\ : Odrv4
    port map (
            O => \N__27847\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__4688\ : InMux
    port map (
            O => \N__27842\,
            I => \N__27839\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__27839\,
            I => \N__27836\
        );

    \I__4686\ : Span4Mux_v
    port map (
            O => \N__27836\,
            I => \N__27831\
        );

    \I__4685\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27828\
        );

    \I__4684\ : InMux
    port map (
            O => \N__27834\,
            I => \N__27825\
        );

    \I__4683\ : Odrv4
    port map (
            O => \N__27831\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__27828\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__27825\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__4680\ : InMux
    port map (
            O => \N__27818\,
            I => \N__27815\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__27815\,
            I => \N__27810\
        );

    \I__4678\ : InMux
    port map (
            O => \N__27814\,
            I => \N__27807\
        );

    \I__4677\ : InMux
    port map (
            O => \N__27813\,
            I => \N__27804\
        );

    \I__4676\ : Span4Mux_h
    port map (
            O => \N__27810\,
            I => \N__27799\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__27807\,
            I => \N__27799\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__27804\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__27799\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4672\ : InMux
    port map (
            O => \N__27794\,
            I => \N__27790\
        );

    \I__4671\ : InMux
    port map (
            O => \N__27793\,
            I => \N__27787\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__27790\,
            I => \N__27784\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__27787\,
            I => \N__27781\
        );

    \I__4668\ : Odrv12
    port map (
            O => \N__27784\,
            I => \phase_controller_inst2.state_RNIG7JFZ0Z_2\
        );

    \I__4667\ : Odrv12
    port map (
            O => \N__27781\,
            I => \phase_controller_inst2.state_RNIG7JFZ0Z_2\
        );

    \I__4666\ : InMux
    port map (
            O => \N__27776\,
            I => \N__27769\
        );

    \I__4665\ : InMux
    port map (
            O => \N__27775\,
            I => \N__27769\
        );

    \I__4664\ : InMux
    port map (
            O => \N__27774\,
            I => \N__27766\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__27769\,
            I => \N__27763\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__27766\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4661\ : Odrv4
    port map (
            O => \N__27763\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4660\ : InMux
    port map (
            O => \N__27758\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__4659\ : InMux
    port map (
            O => \N__27755\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__4658\ : InMux
    port map (
            O => \N__27752\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__4657\ : InMux
    port map (
            O => \N__27749\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__4656\ : InMux
    port map (
            O => \N__27746\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__27743\,
            I => \N__27740\
        );

    \I__4654\ : InMux
    port map (
            O => \N__27740\,
            I => \N__27736\
        );

    \I__4653\ : InMux
    port map (
            O => \N__27739\,
            I => \N__27732\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__27736\,
            I => \N__27729\
        );

    \I__4651\ : InMux
    port map (
            O => \N__27735\,
            I => \N__27726\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__27732\,
            I => \N__27723\
        );

    \I__4649\ : Span4Mux_h
    port map (
            O => \N__27729\,
            I => \N__27720\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__27726\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__27723\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__4646\ : Odrv4
    port map (
            O => \N__27720\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__4645\ : InMux
    port map (
            O => \N__27713\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__4644\ : InMux
    port map (
            O => \N__27710\,
            I => \N__27706\
        );

    \I__4643\ : InMux
    port map (
            O => \N__27709\,
            I => \N__27703\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__27706\,
            I => \N__27699\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__27703\,
            I => \N__27696\
        );

    \I__4640\ : InMux
    port map (
            O => \N__27702\,
            I => \N__27693\
        );

    \I__4639\ : Span4Mux_v
    port map (
            O => \N__27699\,
            I => \N__27690\
        );

    \I__4638\ : Span4Mux_h
    port map (
            O => \N__27696\,
            I => \N__27687\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__27693\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__27690\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__4635\ : Odrv4
    port map (
            O => \N__27687\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__4634\ : InMux
    port map (
            O => \N__27680\,
            I => \bfn_12_9_0_\
        );

    \I__4633\ : CascadeMux
    port map (
            O => \N__27677\,
            I => \N__27673\
        );

    \I__4632\ : InMux
    port map (
            O => \N__27676\,
            I => \N__27668\
        );

    \I__4631\ : InMux
    port map (
            O => \N__27673\,
            I => \N__27668\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__27668\,
            I => \N__27664\
        );

    \I__4629\ : InMux
    port map (
            O => \N__27667\,
            I => \N__27661\
        );

    \I__4628\ : Span4Mux_h
    port map (
            O => \N__27664\,
            I => \N__27658\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__27661\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__4626\ : Odrv4
    port map (
            O => \N__27658\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__4625\ : InMux
    port map (
            O => \N__27653\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__4624\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27646\
        );

    \I__4623\ : InMux
    port map (
            O => \N__27649\,
            I => \N__27643\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__27646\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__27643\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4620\ : InMux
    port map (
            O => \N__27638\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__4619\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27631\
        );

    \I__4618\ : InMux
    port map (
            O => \N__27634\,
            I => \N__27628\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__27631\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__27628\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4615\ : InMux
    port map (
            O => \N__27623\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__4614\ : InMux
    port map (
            O => \N__27620\,
            I => \N__27616\
        );

    \I__4613\ : InMux
    port map (
            O => \N__27619\,
            I => \N__27613\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__27616\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__27613\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__4610\ : InMux
    port map (
            O => \N__27608\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__4609\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27601\
        );

    \I__4608\ : InMux
    port map (
            O => \N__27604\,
            I => \N__27598\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__27601\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__27598\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__4605\ : InMux
    port map (
            O => \N__27593\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__4604\ : InMux
    port map (
            O => \N__27590\,
            I => \N__27586\
        );

    \I__4603\ : InMux
    port map (
            O => \N__27589\,
            I => \N__27583\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__27586\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__27583\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__4600\ : InMux
    port map (
            O => \N__27578\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__4599\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27571\
        );

    \I__4598\ : InMux
    port map (
            O => \N__27574\,
            I => \N__27568\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__27571\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__27568\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__4595\ : InMux
    port map (
            O => \N__27563\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__4594\ : InMux
    port map (
            O => \N__27560\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__4593\ : InMux
    port map (
            O => \N__27557\,
            I => \bfn_12_8_0_\
        );

    \I__4592\ : CascadeMux
    port map (
            O => \N__27554\,
            I => \N__27550\
        );

    \I__4591\ : InMux
    port map (
            O => \N__27553\,
            I => \N__27544\
        );

    \I__4590\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27544\
        );

    \I__4589\ : InMux
    port map (
            O => \N__27549\,
            I => \N__27541\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__27544\,
            I => \N__27538\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__27541\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4586\ : Odrv4
    port map (
            O => \N__27538\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4585\ : InMux
    port map (
            O => \N__27533\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__4584\ : InMux
    port map (
            O => \N__27530\,
            I => \N__27526\
        );

    \I__4583\ : InMux
    port map (
            O => \N__27529\,
            I => \N__27523\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__27526\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__27523\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4580\ : InMux
    port map (
            O => \N__27518\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__4579\ : CascadeMux
    port map (
            O => \N__27515\,
            I => \N__27512\
        );

    \I__4578\ : InMux
    port map (
            O => \N__27512\,
            I => \N__27509\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__27509\,
            I => \N__27506\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__27506\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28\
        );

    \I__4575\ : InMux
    port map (
            O => \N__27503\,
            I => \N__27499\
        );

    \I__4574\ : InMux
    port map (
            O => \N__27502\,
            I => \N__27496\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__27499\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__27496\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4571\ : InMux
    port map (
            O => \N__27491\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__4570\ : InMux
    port map (
            O => \N__27488\,
            I => \N__27484\
        );

    \I__4569\ : InMux
    port map (
            O => \N__27487\,
            I => \N__27481\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__27484\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__27481\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__4566\ : InMux
    port map (
            O => \N__27476\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__4565\ : InMux
    port map (
            O => \N__27473\,
            I => \N__27469\
        );

    \I__4564\ : InMux
    port map (
            O => \N__27472\,
            I => \N__27466\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__27469\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__27466\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__4561\ : InMux
    port map (
            O => \N__27461\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__4560\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27454\
        );

    \I__4559\ : InMux
    port map (
            O => \N__27457\,
            I => \N__27451\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__27454\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__27451\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__4556\ : InMux
    port map (
            O => \N__27446\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__4555\ : InMux
    port map (
            O => \N__27443\,
            I => \N__27439\
        );

    \I__4554\ : InMux
    port map (
            O => \N__27442\,
            I => \N__27436\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__27439\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__27436\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__4551\ : InMux
    port map (
            O => \N__27431\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__4550\ : InMux
    port map (
            O => \N__27428\,
            I => \N__27424\
        );

    \I__4549\ : InMux
    port map (
            O => \N__27427\,
            I => \N__27421\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__27424\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__27421\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__4546\ : InMux
    port map (
            O => \N__27416\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__4545\ : InMux
    port map (
            O => \N__27413\,
            I => \N__27409\
        );

    \I__4544\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27406\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__27409\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__27406\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__4541\ : InMux
    port map (
            O => \N__27401\,
            I => \bfn_12_7_0_\
        );

    \I__4540\ : InMux
    port map (
            O => \N__27398\,
            I => \N__27395\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__27395\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__4538\ : InMux
    port map (
            O => \N__27392\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__4537\ : IoInMux
    port map (
            O => \N__27389\,
            I => \N__27386\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__27386\,
            I => \N__27383\
        );

    \I__4535\ : IoSpan4Mux
    port map (
            O => \N__27383\,
            I => \N__27380\
        );

    \I__4534\ : Sp12to4
    port map (
            O => \N__27380\,
            I => \N__27377\
        );

    \I__4533\ : Span12Mux_s9_v
    port map (
            O => \N__27377\,
            I => \N__27374\
        );

    \I__4532\ : Span12Mux_h
    port map (
            O => \N__27374\,
            I => \N__27371\
        );

    \I__4531\ : Span12Mux_v
    port map (
            O => \N__27371\,
            I => \N__27368\
        );

    \I__4530\ : Odrv12
    port map (
            O => \N__27368\,
            I => pwm_output_c
        );

    \I__4529\ : IoInMux
    port map (
            O => \N__27365\,
            I => \N__27362\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__27362\,
            I => \N__27359\
        );

    \I__4527\ : Span12Mux_s3_v
    port map (
            O => \N__27359\,
            I => \N__27356\
        );

    \I__4526\ : Odrv12
    port map (
            O => \N__27356\,
            I => s3_phy_c
        );

    \I__4525\ : InMux
    port map (
            O => \N__27353\,
            I => \N__27350\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__27350\,
            I => \N__27347\
        );

    \I__4523\ : Span4Mux_v
    port map (
            O => \N__27347\,
            I => \N__27344\
        );

    \I__4522\ : Odrv4
    port map (
            O => \N__27344\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__4521\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27335\
        );

    \I__4520\ : InMux
    port map (
            O => \N__27340\,
            I => \N__27335\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__27335\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\
        );

    \I__4518\ : InMux
    port map (
            O => \N__27332\,
            I => \N__27329\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__27329\,
            I => \N__27324\
        );

    \I__4516\ : InMux
    port map (
            O => \N__27328\,
            I => \N__27321\
        );

    \I__4515\ : InMux
    port map (
            O => \N__27327\,
            I => \N__27318\
        );

    \I__4514\ : Span4Mux_h
    port map (
            O => \N__27324\,
            I => \N__27315\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__27321\,
            I => \N__27312\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__27318\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__4511\ : Odrv4
    port map (
            O => \N__27315\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__27312\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__4509\ : InMux
    port map (
            O => \N__27305\,
            I => \N__27302\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__27302\,
            I => \N__27298\
        );

    \I__4507\ : InMux
    port map (
            O => \N__27301\,
            I => \N__27293\
        );

    \I__4506\ : Span4Mux_h
    port map (
            O => \N__27298\,
            I => \N__27290\
        );

    \I__4505\ : InMux
    port map (
            O => \N__27297\,
            I => \N__27285\
        );

    \I__4504\ : InMux
    port map (
            O => \N__27296\,
            I => \N__27285\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__27293\,
            I => \N__27282\
        );

    \I__4502\ : Span4Mux_v
    port map (
            O => \N__27290\,
            I => \N__27277\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__27285\,
            I => \N__27277\
        );

    \I__4500\ : Span4Mux_v
    port map (
            O => \N__27282\,
            I => \N__27274\
        );

    \I__4499\ : Span4Mux_h
    port map (
            O => \N__27277\,
            I => \N__27271\
        );

    \I__4498\ : Odrv4
    port map (
            O => \N__27274\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__4497\ : Odrv4
    port map (
            O => \N__27271\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__27266\,
            I => \N__27263\
        );

    \I__4495\ : InMux
    port map (
            O => \N__27263\,
            I => \N__27260\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__27260\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\
        );

    \I__4493\ : InMux
    port map (
            O => \N__27257\,
            I => \N__27254\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__27254\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__4491\ : InMux
    port map (
            O => \N__27251\,
            I => \N__27248\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__27248\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__4489\ : InMux
    port map (
            O => \N__27245\,
            I => \N__27242\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__27242\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__4487\ : InMux
    port map (
            O => \N__27239\,
            I => \N__27236\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__27236\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__4485\ : InMux
    port map (
            O => \N__27233\,
            I => \N__27230\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__27230\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__4483\ : InMux
    port map (
            O => \N__27227\,
            I => \N__27224\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__27224\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__4481\ : InMux
    port map (
            O => \N__27221\,
            I => \N__27218\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__27218\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__4479\ : InMux
    port map (
            O => \N__27215\,
            I => \N__27212\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__27212\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__4477\ : InMux
    port map (
            O => \N__27209\,
            I => \N__27206\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__27206\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__4475\ : CascadeMux
    port map (
            O => \N__27203\,
            I => \N__27200\
        );

    \I__4474\ : InMux
    port map (
            O => \N__27200\,
            I => \N__27197\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__27197\,
            I => \N__27194\
        );

    \I__4472\ : Odrv4
    port map (
            O => \N__27194\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__4471\ : InMux
    port map (
            O => \N__27191\,
            I => \N__27184\
        );

    \I__4470\ : InMux
    port map (
            O => \N__27190\,
            I => \N__27184\
        );

    \I__4469\ : InMux
    port map (
            O => \N__27189\,
            I => \N__27181\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__27184\,
            I => \N__27177\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__27181\,
            I => \N__27174\
        );

    \I__4466\ : InMux
    port map (
            O => \N__27180\,
            I => \N__27171\
        );

    \I__4465\ : Span4Mux_h
    port map (
            O => \N__27177\,
            I => \N__27168\
        );

    \I__4464\ : Span4Mux_v
    port map (
            O => \N__27174\,
            I => \N__27163\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__27171\,
            I => \N__27163\
        );

    \I__4462\ : Odrv4
    port map (
            O => \N__27168\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__27163\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__4460\ : CascadeMux
    port map (
            O => \N__27158\,
            I => \N__27155\
        );

    \I__4459\ : InMux
    port map (
            O => \N__27155\,
            I => \N__27149\
        );

    \I__4458\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27149\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__27149\,
            I => \N__27145\
        );

    \I__4456\ : InMux
    port map (
            O => \N__27148\,
            I => \N__27142\
        );

    \I__4455\ : Odrv4
    port map (
            O => \N__27145\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__27142\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__4453\ : InMux
    port map (
            O => \N__27137\,
            I => \N__27134\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__27134\,
            I => \N__27131\
        );

    \I__4451\ : Odrv4
    port map (
            O => \N__27131\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__4450\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27123\
        );

    \I__4449\ : InMux
    port map (
            O => \N__27127\,
            I => \N__27120\
        );

    \I__4448\ : InMux
    port map (
            O => \N__27126\,
            I => \N__27116\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__27123\,
            I => \N__27113\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__27120\,
            I => \N__27110\
        );

    \I__4445\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27107\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__27116\,
            I => \N__27104\
        );

    \I__4443\ : Span4Mux_v
    port map (
            O => \N__27113\,
            I => \N__27097\
        );

    \I__4442\ : Span4Mux_v
    port map (
            O => \N__27110\,
            I => \N__27097\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__27107\,
            I => \N__27097\
        );

    \I__4440\ : Span4Mux_v
    port map (
            O => \N__27104\,
            I => \N__27094\
        );

    \I__4439\ : Span4Mux_h
    port map (
            O => \N__27097\,
            I => \N__27091\
        );

    \I__4438\ : Odrv4
    port map (
            O => \N__27094\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__4437\ : Odrv4
    port map (
            O => \N__27091\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__4436\ : InMux
    port map (
            O => \N__27086\,
            I => \N__27081\
        );

    \I__4435\ : CascadeMux
    port map (
            O => \N__27085\,
            I => \N__27078\
        );

    \I__4434\ : CascadeMux
    port map (
            O => \N__27084\,
            I => \N__27075\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__27081\,
            I => \N__27072\
        );

    \I__4432\ : InMux
    port map (
            O => \N__27078\,
            I => \N__27069\
        );

    \I__4431\ : InMux
    port map (
            O => \N__27075\,
            I => \N__27066\
        );

    \I__4430\ : Span4Mux_h
    port map (
            O => \N__27072\,
            I => \N__27063\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__27069\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__27066\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__27063\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__4426\ : CascadeMux
    port map (
            O => \N__27056\,
            I => \N__27052\
        );

    \I__4425\ : InMux
    port map (
            O => \N__27055\,
            I => \N__27048\
        );

    \I__4424\ : InMux
    port map (
            O => \N__27052\,
            I => \N__27045\
        );

    \I__4423\ : InMux
    port map (
            O => \N__27051\,
            I => \N__27041\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__27048\,
            I => \N__27038\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__27045\,
            I => \N__27035\
        );

    \I__4420\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27032\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__27041\,
            I => \N__27029\
        );

    \I__4418\ : Span4Mux_v
    port map (
            O => \N__27038\,
            I => \N__27022\
        );

    \I__4417\ : Span4Mux_h
    port map (
            O => \N__27035\,
            I => \N__27022\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__27032\,
            I => \N__27022\
        );

    \I__4415\ : Span4Mux_h
    port map (
            O => \N__27029\,
            I => \N__27019\
        );

    \I__4414\ : Span4Mux_h
    port map (
            O => \N__27022\,
            I => \N__27016\
        );

    \I__4413\ : Odrv4
    port map (
            O => \N__27019\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__4412\ : Odrv4
    port map (
            O => \N__27016\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__4411\ : InMux
    port map (
            O => \N__27011\,
            I => \N__27006\
        );

    \I__4410\ : InMux
    port map (
            O => \N__27010\,
            I => \N__27003\
        );

    \I__4409\ : InMux
    port map (
            O => \N__27009\,
            I => \N__27000\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__27006\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__27003\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__27000\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__4405\ : InMux
    port map (
            O => \N__26993\,
            I => \N__26989\
        );

    \I__4404\ : InMux
    port map (
            O => \N__26992\,
            I => \N__26978\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__26989\,
            I => \N__26973\
        );

    \I__4402\ : InMux
    port map (
            O => \N__26988\,
            I => \N__26966\
        );

    \I__4401\ : InMux
    port map (
            O => \N__26987\,
            I => \N__26966\
        );

    \I__4400\ : InMux
    port map (
            O => \N__26986\,
            I => \N__26966\
        );

    \I__4399\ : InMux
    port map (
            O => \N__26985\,
            I => \N__26961\
        );

    \I__4398\ : InMux
    port map (
            O => \N__26984\,
            I => \N__26958\
        );

    \I__4397\ : InMux
    port map (
            O => \N__26983\,
            I => \N__26951\
        );

    \I__4396\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26951\
        );

    \I__4395\ : InMux
    port map (
            O => \N__26981\,
            I => \N__26951\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__26978\,
            I => \N__26948\
        );

    \I__4393\ : InMux
    port map (
            O => \N__26977\,
            I => \N__26943\
        );

    \I__4392\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26943\
        );

    \I__4391\ : Span4Mux_v
    port map (
            O => \N__26973\,
            I => \N__26931\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__26966\,
            I => \N__26931\
        );

    \I__4389\ : InMux
    port map (
            O => \N__26965\,
            I => \N__26926\
        );

    \I__4388\ : InMux
    port map (
            O => \N__26964\,
            I => \N__26926\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__26961\,
            I => \N__26923\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__26958\,
            I => \N__26912\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__26951\,
            I => \N__26912\
        );

    \I__4384\ : Span4Mux_h
    port map (
            O => \N__26948\,
            I => \N__26912\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__26943\,
            I => \N__26912\
        );

    \I__4382\ : InMux
    port map (
            O => \N__26942\,
            I => \N__26895\
        );

    \I__4381\ : InMux
    port map (
            O => \N__26941\,
            I => \N__26895\
        );

    \I__4380\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26895\
        );

    \I__4379\ : InMux
    port map (
            O => \N__26939\,
            I => \N__26895\
        );

    \I__4378\ : InMux
    port map (
            O => \N__26938\,
            I => \N__26895\
        );

    \I__4377\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26895\
        );

    \I__4376\ : InMux
    port map (
            O => \N__26936\,
            I => \N__26895\
        );

    \I__4375\ : Span4Mux_v
    port map (
            O => \N__26931\,
            I => \N__26890\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__26926\,
            I => \N__26890\
        );

    \I__4373\ : Span4Mux_h
    port map (
            O => \N__26923\,
            I => \N__26887\
        );

    \I__4372\ : InMux
    port map (
            O => \N__26922\,
            I => \N__26884\
        );

    \I__4371\ : InMux
    port map (
            O => \N__26921\,
            I => \N__26881\
        );

    \I__4370\ : Span4Mux_v
    port map (
            O => \N__26912\,
            I => \N__26878\
        );

    \I__4369\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26873\
        );

    \I__4368\ : InMux
    port map (
            O => \N__26910\,
            I => \N__26873\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__26895\,
            I => \N__26866\
        );

    \I__4366\ : Span4Mux_v
    port map (
            O => \N__26890\,
            I => \N__26866\
        );

    \I__4365\ : Span4Mux_v
    port map (
            O => \N__26887\,
            I => \N__26866\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__26884\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__26881\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__4362\ : Odrv4
    port map (
            O => \N__26878\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__26873\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__4360\ : Odrv4
    port map (
            O => \N__26866\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__4359\ : InMux
    port map (
            O => \N__26855\,
            I => \N__26852\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__26852\,
            I => \N__26849\
        );

    \I__4357\ : Span4Mux_v
    port map (
            O => \N__26849\,
            I => \N__26846\
        );

    \I__4356\ : Odrv4
    port map (
            O => \N__26846\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__4355\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26840\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__26840\,
            I => \N__26837\
        );

    \I__4353\ : Odrv12
    port map (
            O => \N__26837\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__4352\ : InMux
    port map (
            O => \N__26834\,
            I => \N__26801\
        );

    \I__4351\ : InMux
    port map (
            O => \N__26833\,
            I => \N__26801\
        );

    \I__4350\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26801\
        );

    \I__4349\ : InMux
    port map (
            O => \N__26831\,
            I => \N__26801\
        );

    \I__4348\ : InMux
    port map (
            O => \N__26830\,
            I => \N__26801\
        );

    \I__4347\ : InMux
    port map (
            O => \N__26829\,
            I => \N__26801\
        );

    \I__4346\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26801\
        );

    \I__4345\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26801\
        );

    \I__4344\ : InMux
    port map (
            O => \N__26826\,
            I => \N__26784\
        );

    \I__4343\ : InMux
    port map (
            O => \N__26825\,
            I => \N__26784\
        );

    \I__4342\ : InMux
    port map (
            O => \N__26824\,
            I => \N__26784\
        );

    \I__4341\ : InMux
    port map (
            O => \N__26823\,
            I => \N__26784\
        );

    \I__4340\ : InMux
    port map (
            O => \N__26822\,
            I => \N__26784\
        );

    \I__4339\ : InMux
    port map (
            O => \N__26821\,
            I => \N__26784\
        );

    \I__4338\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26784\
        );

    \I__4337\ : InMux
    port map (
            O => \N__26819\,
            I => \N__26784\
        );

    \I__4336\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26781\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__26801\,
            I => \N__26775\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__26784\,
            I => \N__26775\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__26781\,
            I => \N__26772\
        );

    \I__4332\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26769\
        );

    \I__4331\ : Span4Mux_s3_h
    port map (
            O => \N__26775\,
            I => \N__26766\
        );

    \I__4330\ : Span4Mux_v
    port map (
            O => \N__26772\,
            I => \N__26763\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__26769\,
            I => \N__26760\
        );

    \I__4328\ : Span4Mux_v
    port map (
            O => \N__26766\,
            I => \N__26757\
        );

    \I__4327\ : Span4Mux_h
    port map (
            O => \N__26763\,
            I => \N__26754\
        );

    \I__4326\ : Span4Mux_s3_h
    port map (
            O => \N__26760\,
            I => \N__26751\
        );

    \I__4325\ : Span4Mux_h
    port map (
            O => \N__26757\,
            I => \N__26748\
        );

    \I__4324\ : Span4Mux_v
    port map (
            O => \N__26754\,
            I => \N__26743\
        );

    \I__4323\ : Span4Mux_h
    port map (
            O => \N__26751\,
            I => \N__26743\
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__26748\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__4321\ : Odrv4
    port map (
            O => \N__26743\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__4320\ : InMux
    port map (
            O => \N__26738\,
            I => \N__26735\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__26735\,
            I => \N__26732\
        );

    \I__4318\ : Odrv4
    port map (
            O => \N__26732\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__4317\ : InMux
    port map (
            O => \N__26729\,
            I => \N__26726\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__26726\,
            I => \N__26723\
        );

    \I__4315\ : Odrv4
    port map (
            O => \N__26723\,
            I => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\
        );

    \I__4314\ : InMux
    port map (
            O => \N__26720\,
            I => \N__26717\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__26717\,
            I => \N__26714\
        );

    \I__4312\ : Odrv4
    port map (
            O => \N__26714\,
            I => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\
        );

    \I__4311\ : InMux
    port map (
            O => \N__26711\,
            I => \N__26708\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__26708\,
            I => \N__26705\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__26705\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__26702\,
            I => \N__26699\
        );

    \I__4307\ : InMux
    port map (
            O => \N__26699\,
            I => \N__26696\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__26696\,
            I => \N__26693\
        );

    \I__4305\ : Span4Mux_v
    port map (
            O => \N__26693\,
            I => \N__26690\
        );

    \I__4304\ : Odrv4
    port map (
            O => \N__26690\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__4303\ : CascadeMux
    port map (
            O => \N__26687\,
            I => \N__26684\
        );

    \I__4302\ : InMux
    port map (
            O => \N__26684\,
            I => \N__26681\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__26681\,
            I => \N__26678\
        );

    \I__4300\ : Span4Mux_v
    port map (
            O => \N__26678\,
            I => \N__26675\
        );

    \I__4299\ : Odrv4
    port map (
            O => \N__26675\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__4298\ : CascadeMux
    port map (
            O => \N__26672\,
            I => \N__26669\
        );

    \I__4297\ : InMux
    port map (
            O => \N__26669\,
            I => \N__26666\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__26666\,
            I => \N__26663\
        );

    \I__4295\ : Odrv4
    port map (
            O => \N__26663\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__4294\ : InMux
    port map (
            O => \N__26660\,
            I => \N__26657\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__26657\,
            I => \N__26654\
        );

    \I__4292\ : Span4Mux_h
    port map (
            O => \N__26654\,
            I => \N__26651\
        );

    \I__4291\ : Odrv4
    port map (
            O => \N__26651\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__4290\ : CascadeMux
    port map (
            O => \N__26648\,
            I => \N__26644\
        );

    \I__4289\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26639\
        );

    \I__4288\ : InMux
    port map (
            O => \N__26644\,
            I => \N__26636\
        );

    \I__4287\ : InMux
    port map (
            O => \N__26643\,
            I => \N__26633\
        );

    \I__4286\ : InMux
    port map (
            O => \N__26642\,
            I => \N__26630\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__26639\,
            I => \N__26625\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__26636\,
            I => \N__26625\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__26633\,
            I => \N__26620\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__26630\,
            I => \N__26620\
        );

    \I__4281\ : Span4Mux_v
    port map (
            O => \N__26625\,
            I => \N__26617\
        );

    \I__4280\ : Span4Mux_v
    port map (
            O => \N__26620\,
            I => \N__26614\
        );

    \I__4279\ : Odrv4
    port map (
            O => \N__26617\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__4278\ : Odrv4
    port map (
            O => \N__26614\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__4277\ : CascadeMux
    port map (
            O => \N__26609\,
            I => \N__26606\
        );

    \I__4276\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26599\
        );

    \I__4275\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26599\
        );

    \I__4274\ : InMux
    port map (
            O => \N__26604\,
            I => \N__26596\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__26599\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__26596\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__4271\ : InMux
    port map (
            O => \N__26591\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__4270\ : CascadeMux
    port map (
            O => \N__26588\,
            I => \N__26585\
        );

    \I__4269\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26582\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__26582\,
            I => \N__26579\
        );

    \I__4267\ : Span4Mux_h
    port map (
            O => \N__26579\,
            I => \N__26576\
        );

    \I__4266\ : Odrv4
    port map (
            O => \N__26576\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__4265\ : InMux
    port map (
            O => \N__26573\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__4264\ : InMux
    port map (
            O => \N__26570\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__4263\ : CascadeMux
    port map (
            O => \N__26567\,
            I => \N__26563\
        );

    \I__4262\ : CascadeMux
    port map (
            O => \N__26566\,
            I => \N__26560\
        );

    \I__4261\ : InMux
    port map (
            O => \N__26563\,
            I => \N__26557\
        );

    \I__4260\ : InMux
    port map (
            O => \N__26560\,
            I => \N__26554\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__26557\,
            I => \N__26551\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__26554\,
            I => \N__26546\
        );

    \I__4257\ : Span4Mux_v
    port map (
            O => \N__26551\,
            I => \N__26543\
        );

    \I__4256\ : InMux
    port map (
            O => \N__26550\,
            I => \N__26538\
        );

    \I__4255\ : InMux
    port map (
            O => \N__26549\,
            I => \N__26538\
        );

    \I__4254\ : Span4Mux_h
    port map (
            O => \N__26546\,
            I => \N__26531\
        );

    \I__4253\ : Span4Mux_h
    port map (
            O => \N__26543\,
            I => \N__26531\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__26538\,
            I => \N__26531\
        );

    \I__4251\ : Odrv4
    port map (
            O => \N__26531\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__4250\ : InMux
    port map (
            O => \N__26528\,
            I => \N__26523\
        );

    \I__4249\ : InMux
    port map (
            O => \N__26527\,
            I => \N__26520\
        );

    \I__4248\ : InMux
    port map (
            O => \N__26526\,
            I => \N__26517\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__26523\,
            I => \N__26514\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__26520\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__26517\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__26514\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__4243\ : CascadeMux
    port map (
            O => \N__26507\,
            I => \N__26504\
        );

    \I__4242\ : InMux
    port map (
            O => \N__26504\,
            I => \N__26501\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__26501\,
            I => \N__26498\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__26498\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__4239\ : InMux
    port map (
            O => \N__26495\,
            I => \N__26492\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__26492\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__4237\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26486\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__26486\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__4235\ : CascadeMux
    port map (
            O => \N__26483\,
            I => \N__26480\
        );

    \I__4234\ : InMux
    port map (
            O => \N__26480\,
            I => \N__26477\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__26477\,
            I => \N__26474\
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__26474\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__4231\ : InMux
    port map (
            O => \N__26471\,
            I => \N__26468\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__26468\,
            I => \N__26465\
        );

    \I__4229\ : Odrv4
    port map (
            O => \N__26465\,
            I => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\
        );

    \I__4228\ : CascadeMux
    port map (
            O => \N__26462\,
            I => \N__26459\
        );

    \I__4227\ : InMux
    port map (
            O => \N__26459\,
            I => \N__26456\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__26456\,
            I => \N__26453\
        );

    \I__4225\ : Odrv12
    port map (
            O => \N__26453\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__4224\ : InMux
    port map (
            O => \N__26450\,
            I => \N__26447\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__26447\,
            I => \N__26444\
        );

    \I__4222\ : Span4Mux_h
    port map (
            O => \N__26444\,
            I => \N__26441\
        );

    \I__4221\ : Odrv4
    port map (
            O => \N__26441\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__4220\ : InMux
    port map (
            O => \N__26438\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__4219\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26432\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__26432\,
            I => \N__26429\
        );

    \I__4217\ : Span4Mux_v
    port map (
            O => \N__26429\,
            I => \N__26426\
        );

    \I__4216\ : Odrv4
    port map (
            O => \N__26426\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__4215\ : InMux
    port map (
            O => \N__26423\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__4214\ : InMux
    port map (
            O => \N__26420\,
            I => \N__26417\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__26417\,
            I => \N__26414\
        );

    \I__4212\ : Span4Mux_h
    port map (
            O => \N__26414\,
            I => \N__26411\
        );

    \I__4211\ : Odrv4
    port map (
            O => \N__26411\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__4210\ : InMux
    port map (
            O => \N__26408\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__4209\ : InMux
    port map (
            O => \N__26405\,
            I => \N__26402\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__26402\,
            I => \N__26399\
        );

    \I__4207\ : Span4Mux_h
    port map (
            O => \N__26399\,
            I => \N__26396\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__26396\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__4205\ : InMux
    port map (
            O => \N__26393\,
            I => \bfn_11_18_0_\
        );

    \I__4204\ : InMux
    port map (
            O => \N__26390\,
            I => \N__26387\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__26387\,
            I => \N__26384\
        );

    \I__4202\ : Span4Mux_h
    port map (
            O => \N__26384\,
            I => \N__26381\
        );

    \I__4201\ : Odrv4
    port map (
            O => \N__26381\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__4200\ : InMux
    port map (
            O => \N__26378\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__4199\ : InMux
    port map (
            O => \N__26375\,
            I => \N__26372\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__26372\,
            I => \N__26369\
        );

    \I__4197\ : Span4Mux_h
    port map (
            O => \N__26369\,
            I => \N__26366\
        );

    \I__4196\ : Odrv4
    port map (
            O => \N__26366\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__4195\ : InMux
    port map (
            O => \N__26363\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__4194\ : InMux
    port map (
            O => \N__26360\,
            I => \N__26357\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__26357\,
            I => \N__26354\
        );

    \I__4192\ : Span4Mux_h
    port map (
            O => \N__26354\,
            I => \N__26351\
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__26351\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__4190\ : InMux
    port map (
            O => \N__26348\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__4189\ : InMux
    port map (
            O => \N__26345\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__4188\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26339\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__26339\,
            I => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__26336\,
            I => \N__26333\
        );

    \I__4185\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26330\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__26330\,
            I => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__26327\,
            I => \N__26324\
        );

    \I__4182\ : InMux
    port map (
            O => \N__26324\,
            I => \N__26321\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__26321\,
            I => \N__26318\
        );

    \I__4180\ : Span4Mux_v
    port map (
            O => \N__26318\,
            I => \N__26315\
        );

    \I__4179\ : Odrv4
    port map (
            O => \N__26315\,
            I => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\
        );

    \I__4178\ : InMux
    port map (
            O => \N__26312\,
            I => \N__26309\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__26309\,
            I => \N__26306\
        );

    \I__4176\ : Odrv4
    port map (
            O => \N__26306\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__4175\ : InMux
    port map (
            O => \N__26303\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__4174\ : InMux
    port map (
            O => \N__26300\,
            I => \N__26297\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__26297\,
            I => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__26294\,
            I => \N__26291\
        );

    \I__4171\ : InMux
    port map (
            O => \N__26291\,
            I => \N__26288\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__26288\,
            I => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\
        );

    \I__4169\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26282\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__26282\,
            I => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\
        );

    \I__4167\ : CascadeMux
    port map (
            O => \N__26279\,
            I => \N__26276\
        );

    \I__4166\ : InMux
    port map (
            O => \N__26276\,
            I => \N__26273\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__26273\,
            I => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26270\,
            I => \N__26267\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__26267\,
            I => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\
        );

    \I__4162\ : CascadeMux
    port map (
            O => \N__26264\,
            I => \N__26261\
        );

    \I__4161\ : InMux
    port map (
            O => \N__26261\,
            I => \N__26258\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__26258\,
            I => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__26255\,
            I => \N__26252\
        );

    \I__4158\ : InMux
    port map (
            O => \N__26252\,
            I => \N__26249\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__26249\,
            I => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\
        );

    \I__4156\ : InMux
    port map (
            O => \N__26246\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__4155\ : InMux
    port map (
            O => \N__26243\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__4154\ : InMux
    port map (
            O => \N__26240\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__4153\ : CascadeMux
    port map (
            O => \N__26237\,
            I => \N__26233\
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__26236\,
            I => \N__26229\
        );

    \I__4151\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26222\
        );

    \I__4150\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26222\
        );

    \I__4149\ : InMux
    port map (
            O => \N__26229\,
            I => \N__26222\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__26222\,
            I => \N__26218\
        );

    \I__4147\ : InMux
    port map (
            O => \N__26221\,
            I => \N__26215\
        );

    \I__4146\ : Sp12to4
    port map (
            O => \N__26218\,
            I => \N__26212\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__26215\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__4144\ : Odrv12
    port map (
            O => \N__26212\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__4143\ : InMux
    port map (
            O => \N__26207\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__4142\ : IoInMux
    port map (
            O => \N__26204\,
            I => \N__26189\
        );

    \I__4141\ : InMux
    port map (
            O => \N__26203\,
            I => \N__26186\
        );

    \I__4140\ : InMux
    port map (
            O => \N__26202\,
            I => \N__26177\
        );

    \I__4139\ : InMux
    port map (
            O => \N__26201\,
            I => \N__26177\
        );

    \I__4138\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26177\
        );

    \I__4137\ : InMux
    port map (
            O => \N__26199\,
            I => \N__26177\
        );

    \I__4136\ : InMux
    port map (
            O => \N__26198\,
            I => \N__26170\
        );

    \I__4135\ : InMux
    port map (
            O => \N__26197\,
            I => \N__26170\
        );

    \I__4134\ : InMux
    port map (
            O => \N__26196\,
            I => \N__26170\
        );

    \I__4133\ : InMux
    port map (
            O => \N__26195\,
            I => \N__26161\
        );

    \I__4132\ : InMux
    port map (
            O => \N__26194\,
            I => \N__26161\
        );

    \I__4131\ : InMux
    port map (
            O => \N__26193\,
            I => \N__26161\
        );

    \I__4130\ : InMux
    port map (
            O => \N__26192\,
            I => \N__26161\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__26189\,
            I => \N__26139\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__26186\,
            I => \N__26130\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__26177\,
            I => \N__26130\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__26170\,
            I => \N__26130\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__26161\,
            I => \N__26130\
        );

    \I__4124\ : InMux
    port map (
            O => \N__26160\,
            I => \N__26121\
        );

    \I__4123\ : InMux
    port map (
            O => \N__26159\,
            I => \N__26121\
        );

    \I__4122\ : InMux
    port map (
            O => \N__26158\,
            I => \N__26121\
        );

    \I__4121\ : InMux
    port map (
            O => \N__26157\,
            I => \N__26121\
        );

    \I__4120\ : InMux
    port map (
            O => \N__26156\,
            I => \N__26112\
        );

    \I__4119\ : InMux
    port map (
            O => \N__26155\,
            I => \N__26112\
        );

    \I__4118\ : InMux
    port map (
            O => \N__26154\,
            I => \N__26112\
        );

    \I__4117\ : InMux
    port map (
            O => \N__26153\,
            I => \N__26112\
        );

    \I__4116\ : InMux
    port map (
            O => \N__26152\,
            I => \N__26103\
        );

    \I__4115\ : InMux
    port map (
            O => \N__26151\,
            I => \N__26103\
        );

    \I__4114\ : InMux
    port map (
            O => \N__26150\,
            I => \N__26103\
        );

    \I__4113\ : InMux
    port map (
            O => \N__26149\,
            I => \N__26103\
        );

    \I__4112\ : InMux
    port map (
            O => \N__26148\,
            I => \N__26094\
        );

    \I__4111\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26094\
        );

    \I__4110\ : InMux
    port map (
            O => \N__26146\,
            I => \N__26094\
        );

    \I__4109\ : InMux
    port map (
            O => \N__26145\,
            I => \N__26094\
        );

    \I__4108\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26087\
        );

    \I__4107\ : InMux
    port map (
            O => \N__26143\,
            I => \N__26087\
        );

    \I__4106\ : InMux
    port map (
            O => \N__26142\,
            I => \N__26087\
        );

    \I__4105\ : Span4Mux_s0_v
    port map (
            O => \N__26139\,
            I => \N__26084\
        );

    \I__4104\ : Span4Mux_v
    port map (
            O => \N__26130\,
            I => \N__26081\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__26121\,
            I => \N__26070\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__26112\,
            I => \N__26070\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__26103\,
            I => \N__26070\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__26094\,
            I => \N__26070\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__26087\,
            I => \N__26070\
        );

    \I__4098\ : Sp12to4
    port map (
            O => \N__26084\,
            I => \N__26067\
        );

    \I__4097\ : Span4Mux_h
    port map (
            O => \N__26081\,
            I => \N__26062\
        );

    \I__4096\ : Span4Mux_v
    port map (
            O => \N__26070\,
            I => \N__26062\
        );

    \I__4095\ : Span12Mux_s5_h
    port map (
            O => \N__26067\,
            I => \N__26059\
        );

    \I__4094\ : Span4Mux_h
    port map (
            O => \N__26062\,
            I => \N__26056\
        );

    \I__4093\ : Span12Mux_v
    port map (
            O => \N__26059\,
            I => \N__26053\
        );

    \I__4092\ : Odrv4
    port map (
            O => \N__26056\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4091\ : Odrv12
    port map (
            O => \N__26053\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__4090\ : InMux
    port map (
            O => \N__26048\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__4089\ : CascadeMux
    port map (
            O => \N__26045\,
            I => \N__26041\
        );

    \I__4088\ : InMux
    port map (
            O => \N__26044\,
            I => \N__26033\
        );

    \I__4087\ : InMux
    port map (
            O => \N__26041\,
            I => \N__26033\
        );

    \I__4086\ : InMux
    port map (
            O => \N__26040\,
            I => \N__26033\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__26033\,
            I => \N__26029\
        );

    \I__4084\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26026\
        );

    \I__4083\ : Span4Mux_h
    port map (
            O => \N__26029\,
            I => \N__26023\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__26026\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__4081\ : Odrv4
    port map (
            O => \N__26023\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__26018\,
            I => \N__26015\
        );

    \I__4079\ : InMux
    port map (
            O => \N__26015\,
            I => \N__26012\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__26012\,
            I => \N__26009\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__26009\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__4076\ : CascadeMux
    port map (
            O => \N__26006\,
            I => \N__26003\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26003\,
            I => \N__26000\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__26000\,
            I => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\
        );

    \I__4073\ : CascadeMux
    port map (
            O => \N__25997\,
            I => \N__25993\
        );

    \I__4072\ : CascadeMux
    port map (
            O => \N__25996\,
            I => \N__25990\
        );

    \I__4071\ : InMux
    port map (
            O => \N__25993\,
            I => \N__25987\
        );

    \I__4070\ : InMux
    port map (
            O => \N__25990\,
            I => \N__25984\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__25987\,
            I => \N__25978\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__25984\,
            I => \N__25978\
        );

    \I__4067\ : InMux
    port map (
            O => \N__25983\,
            I => \N__25975\
        );

    \I__4066\ : Span4Mux_h
    port map (
            O => \N__25978\,
            I => \N__25972\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__25975\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4064\ : Odrv4
    port map (
            O => \N__25972\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4063\ : InMux
    port map (
            O => \N__25967\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__4062\ : InMux
    port map (
            O => \N__25964\,
            I => \N__25960\
        );

    \I__4061\ : InMux
    port map (
            O => \N__25963\,
            I => \N__25957\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__25960\,
            I => \N__25951\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__25957\,
            I => \N__25951\
        );

    \I__4058\ : InMux
    port map (
            O => \N__25956\,
            I => \N__25948\
        );

    \I__4057\ : Span4Mux_h
    port map (
            O => \N__25951\,
            I => \N__25945\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__25948\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__25945\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4054\ : InMux
    port map (
            O => \N__25940\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__4053\ : InMux
    port map (
            O => \N__25937\,
            I => \N__25931\
        );

    \I__4052\ : InMux
    port map (
            O => \N__25936\,
            I => \N__25931\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__25931\,
            I => \N__25927\
        );

    \I__4050\ : InMux
    port map (
            O => \N__25930\,
            I => \N__25924\
        );

    \I__4049\ : Span4Mux_h
    port map (
            O => \N__25927\,
            I => \N__25921\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__25924\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__25921\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__4046\ : InMux
    port map (
            O => \N__25916\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__4045\ : CascadeMux
    port map (
            O => \N__25913\,
            I => \N__25909\
        );

    \I__4044\ : InMux
    port map (
            O => \N__25912\,
            I => \N__25904\
        );

    \I__4043\ : InMux
    port map (
            O => \N__25909\,
            I => \N__25904\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__25904\,
            I => \N__25900\
        );

    \I__4041\ : InMux
    port map (
            O => \N__25903\,
            I => \N__25897\
        );

    \I__4040\ : Span4Mux_v
    port map (
            O => \N__25900\,
            I => \N__25894\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__25897\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__4038\ : Odrv4
    port map (
            O => \N__25894\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__4037\ : InMux
    port map (
            O => \N__25889\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__4036\ : CascadeMux
    port map (
            O => \N__25886\,
            I => \N__25882\
        );

    \I__4035\ : InMux
    port map (
            O => \N__25885\,
            I => \N__25877\
        );

    \I__4034\ : InMux
    port map (
            O => \N__25882\,
            I => \N__25877\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__25877\,
            I => \N__25873\
        );

    \I__4032\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25870\
        );

    \I__4031\ : Span4Mux_h
    port map (
            O => \N__25873\,
            I => \N__25867\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__25870\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__4029\ : Odrv4
    port map (
            O => \N__25867\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__4028\ : InMux
    port map (
            O => \N__25862\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__4027\ : InMux
    port map (
            O => \N__25859\,
            I => \N__25853\
        );

    \I__4026\ : InMux
    port map (
            O => \N__25858\,
            I => \N__25853\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__25853\,
            I => \N__25849\
        );

    \I__4024\ : InMux
    port map (
            O => \N__25852\,
            I => \N__25846\
        );

    \I__4023\ : Span4Mux_v
    port map (
            O => \N__25849\,
            I => \N__25843\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__25846\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__25843\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__4020\ : InMux
    port map (
            O => \N__25838\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__4019\ : InMux
    port map (
            O => \N__25835\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__4018\ : InMux
    port map (
            O => \N__25832\,
            I => \bfn_11_14_0_\
        );

    \I__4017\ : InMux
    port map (
            O => \N__25829\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__4016\ : InMux
    port map (
            O => \N__25826\,
            I => \N__25822\
        );

    \I__4015\ : InMux
    port map (
            O => \N__25825\,
            I => \N__25819\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__25822\,
            I => \N__25816\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__25819\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4012\ : Odrv4
    port map (
            O => \N__25816\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__4011\ : InMux
    port map (
            O => \N__25811\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__4010\ : InMux
    port map (
            O => \N__25808\,
            I => \N__25804\
        );

    \I__4009\ : InMux
    port map (
            O => \N__25807\,
            I => \N__25801\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__25804\,
            I => \N__25798\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__25801\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4006\ : Odrv12
    port map (
            O => \N__25798\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__4005\ : InMux
    port map (
            O => \N__25793\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__4004\ : InMux
    port map (
            O => \N__25790\,
            I => \N__25786\
        );

    \I__4003\ : InMux
    port map (
            O => \N__25789\,
            I => \N__25783\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__25786\,
            I => \N__25780\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__25783\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__4000\ : Odrv4
    port map (
            O => \N__25780\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3999\ : InMux
    port map (
            O => \N__25775\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__3998\ : InMux
    port map (
            O => \N__25772\,
            I => \N__25768\
        );

    \I__3997\ : InMux
    port map (
            O => \N__25771\,
            I => \N__25765\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__25768\,
            I => \N__25762\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__25765\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3994\ : Odrv12
    port map (
            O => \N__25762\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3993\ : InMux
    port map (
            O => \N__25757\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__3992\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25750\
        );

    \I__3991\ : InMux
    port map (
            O => \N__25753\,
            I => \N__25747\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__25750\,
            I => \N__25744\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__25747\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3988\ : Odrv12
    port map (
            O => \N__25744\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3987\ : InMux
    port map (
            O => \N__25739\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__3986\ : InMux
    port map (
            O => \N__25736\,
            I => \N__25732\
        );

    \I__3985\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25729\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__25732\,
            I => \N__25726\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__25729\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3982\ : Odrv4
    port map (
            O => \N__25726\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3981\ : InMux
    port map (
            O => \N__25721\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__3980\ : InMux
    port map (
            O => \N__25718\,
            I => \N__25713\
        );

    \I__3979\ : InMux
    port map (
            O => \N__25717\,
            I => \N__25708\
        );

    \I__3978\ : InMux
    port map (
            O => \N__25716\,
            I => \N__25708\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__25713\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__25708\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3975\ : InMux
    port map (
            O => \N__25703\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__3974\ : InMux
    port map (
            O => \N__25700\,
            I => \N__25695\
        );

    \I__3973\ : InMux
    port map (
            O => \N__25699\,
            I => \N__25690\
        );

    \I__3972\ : InMux
    port map (
            O => \N__25698\,
            I => \N__25690\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__25695\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__25690\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3969\ : InMux
    port map (
            O => \N__25685\,
            I => \bfn_11_13_0_\
        );

    \I__3968\ : InMux
    port map (
            O => \N__25682\,
            I => \N__25678\
        );

    \I__3967\ : InMux
    port map (
            O => \N__25681\,
            I => \N__25675\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__25678\,
            I => \N__25672\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__25675\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3964\ : Odrv4
    port map (
            O => \N__25672\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3963\ : InMux
    port map (
            O => \N__25667\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__25664\,
            I => \N__25661\
        );

    \I__3961\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25658\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__25658\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28\
        );

    \I__3959\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25651\
        );

    \I__3958\ : InMux
    port map (
            O => \N__25654\,
            I => \N__25648\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__25651\,
            I => \N__25645\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__25648\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3955\ : Odrv4
    port map (
            O => \N__25645\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3954\ : InMux
    port map (
            O => \N__25640\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__3953\ : InMux
    port map (
            O => \N__25637\,
            I => \N__25634\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__25634\,
            I => \N__25630\
        );

    \I__3951\ : InMux
    port map (
            O => \N__25633\,
            I => \N__25627\
        );

    \I__3950\ : Span4Mux_h
    port map (
            O => \N__25630\,
            I => \N__25624\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__25627\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3948\ : Odrv4
    port map (
            O => \N__25624\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3947\ : InMux
    port map (
            O => \N__25619\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__3946\ : InMux
    port map (
            O => \N__25616\,
            I => \N__25612\
        );

    \I__3945\ : InMux
    port map (
            O => \N__25615\,
            I => \N__25609\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__25612\,
            I => \N__25606\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__25609\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3942\ : Odrv4
    port map (
            O => \N__25606\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3941\ : InMux
    port map (
            O => \N__25601\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__3940\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25594\
        );

    \I__3939\ : InMux
    port map (
            O => \N__25597\,
            I => \N__25591\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__25594\,
            I => \N__25588\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__25591\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3936\ : Odrv12
    port map (
            O => \N__25588\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3935\ : InMux
    port map (
            O => \N__25583\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__3934\ : InMux
    port map (
            O => \N__25580\,
            I => \N__25577\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__25577\,
            I => \N__25573\
        );

    \I__3932\ : InMux
    port map (
            O => \N__25576\,
            I => \N__25570\
        );

    \I__3931\ : Span4Mux_h
    port map (
            O => \N__25573\,
            I => \N__25567\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__25570\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__25567\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3928\ : InMux
    port map (
            O => \N__25562\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__3927\ : InMux
    port map (
            O => \N__25559\,
            I => \N__25555\
        );

    \I__3926\ : InMux
    port map (
            O => \N__25558\,
            I => \N__25552\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__25555\,
            I => \N__25549\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__25552\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3923\ : Odrv4
    port map (
            O => \N__25549\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3922\ : InMux
    port map (
            O => \N__25544\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__3921\ : InMux
    port map (
            O => \N__25541\,
            I => \N__25537\
        );

    \I__3920\ : InMux
    port map (
            O => \N__25540\,
            I => \N__25534\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__25537\,
            I => \N__25531\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__25534\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__25531\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3916\ : InMux
    port map (
            O => \N__25526\,
            I => \bfn_11_12_0_\
        );

    \I__3915\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25520\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__25520\,
            I => \N__25517\
        );

    \I__3913\ : Span4Mux_v
    port map (
            O => \N__25517\,
            I => \N__25514\
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__25514\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__25511\,
            I => \N__25508\
        );

    \I__3910\ : InMux
    port map (
            O => \N__25508\,
            I => \N__25505\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__25505\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt24\
        );

    \I__3908\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25499\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__25499\,
            I => \N__25496\
        );

    \I__3906\ : Odrv12
    port map (
            O => \N__25496\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt26\
        );

    \I__3905\ : CascadeMux
    port map (
            O => \N__25493\,
            I => \N__25490\
        );

    \I__3904\ : InMux
    port map (
            O => \N__25490\,
            I => \N__25487\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__25487\,
            I => \N__25484\
        );

    \I__3902\ : Span4Mux_v
    port map (
            O => \N__25484\,
            I => \N__25481\
        );

    \I__3901\ : Odrv4
    port map (
            O => \N__25481\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\
        );

    \I__3900\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25475\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__25475\,
            I => \N__25472\
        );

    \I__3898\ : Odrv4
    port map (
            O => \N__25472\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\
        );

    \I__3897\ : CascadeMux
    port map (
            O => \N__25469\,
            I => \N__25466\
        );

    \I__3896\ : InMux
    port map (
            O => \N__25466\,
            I => \N__25463\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__25463\,
            I => \N__25460\
        );

    \I__3894\ : Span4Mux_v
    port map (
            O => \N__25460\,
            I => \N__25456\
        );

    \I__3893\ : InMux
    port map (
            O => \N__25459\,
            I => \N__25453\
        );

    \I__3892\ : Odrv4
    port map (
            O => \N__25456\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt30\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__25453\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt30\
        );

    \I__3890\ : InMux
    port map (
            O => \N__25448\,
            I => \N__25445\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__25445\,
            I => \N__25442\
        );

    \I__3888\ : Odrv12
    port map (
            O => \N__25442\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\
        );

    \I__3887\ : InMux
    port map (
            O => \N__25439\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_28\
        );

    \I__3886\ : InMux
    port map (
            O => \N__25436\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30\
        );

    \I__3885\ : InMux
    port map (
            O => \N__25433\,
            I => \N__25430\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__25430\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt28\
        );

    \I__3883\ : InMux
    port map (
            O => \N__25427\,
            I => \N__25424\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__25424\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__25421\,
            I => \N__25417\
        );

    \I__3880\ : InMux
    port map (
            O => \N__25420\,
            I => \N__25413\
        );

    \I__3879\ : InMux
    port map (
            O => \N__25417\,
            I => \N__25410\
        );

    \I__3878\ : InMux
    port map (
            O => \N__25416\,
            I => \N__25407\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__25413\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__25410\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__25407\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3874\ : InMux
    port map (
            O => \N__25400\,
            I => \N__25397\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__25397\,
            I => \N__25394\
        );

    \I__3872\ : Span4Mux_h
    port map (
            O => \N__25394\,
            I => \N__25391\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__25391\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__25388\,
            I => \N__25385\
        );

    \I__3869\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25382\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__25382\,
            I => \N__25379\
        );

    \I__3867\ : Odrv4
    port map (
            O => \N__25379\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__3866\ : InMux
    port map (
            O => \N__25376\,
            I => \N__25373\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__25373\,
            I => \N__25370\
        );

    \I__3864\ : Span4Mux_h
    port map (
            O => \N__25370\,
            I => \N__25367\
        );

    \I__3863\ : Odrv4
    port map (
            O => \N__25367\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__25364\,
            I => \N__25361\
        );

    \I__3861\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25358\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__25358\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__3859\ : CascadeMux
    port map (
            O => \N__25355\,
            I => \N__25352\
        );

    \I__3858\ : InMux
    port map (
            O => \N__25352\,
            I => \N__25349\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__25349\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__3856\ : CascadeMux
    port map (
            O => \N__25346\,
            I => \N__25343\
        );

    \I__3855\ : InMux
    port map (
            O => \N__25343\,
            I => \N__25340\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__25340\,
            I => \N__25337\
        );

    \I__3853\ : Span4Mux_v
    port map (
            O => \N__25337\,
            I => \N__25334\
        );

    \I__3852\ : Odrv4
    port map (
            O => \N__25334\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__3851\ : InMux
    port map (
            O => \N__25331\,
            I => \N__25328\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__25328\,
            I => \N__25325\
        );

    \I__3849\ : Odrv4
    port map (
            O => \N__25325\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__3848\ : InMux
    port map (
            O => \N__25322\,
            I => \N__25319\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__25319\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\
        );

    \I__3846\ : CascadeMux
    port map (
            O => \N__25316\,
            I => \N__25313\
        );

    \I__3845\ : InMux
    port map (
            O => \N__25313\,
            I => \N__25310\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__25310\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt18\
        );

    \I__3843\ : InMux
    port map (
            O => \N__25307\,
            I => \N__25304\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__25304\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__25301\,
            I => \N__25298\
        );

    \I__3840\ : InMux
    port map (
            O => \N__25298\,
            I => \N__25295\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__25295\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__3838\ : CascadeMux
    port map (
            O => \N__25292\,
            I => \N__25289\
        );

    \I__3837\ : InMux
    port map (
            O => \N__25289\,
            I => \N__25286\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__25286\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__3835\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25280\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__25280\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__3833\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25274\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__25274\,
            I => \N__25271\
        );

    \I__3831\ : Odrv4
    port map (
            O => \N__25271\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__25268\,
            I => \N__25265\
        );

    \I__3829\ : InMux
    port map (
            O => \N__25265\,
            I => \N__25262\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__25262\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__3827\ : InMux
    port map (
            O => \N__25259\,
            I => \N__25256\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__25256\,
            I => \N__25253\
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__25253\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__3824\ : CascadeMux
    port map (
            O => \N__25250\,
            I => \N__25247\
        );

    \I__3823\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25244\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__25244\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__25241\,
            I => \N__25238\
        );

    \I__3820\ : InMux
    port map (
            O => \N__25238\,
            I => \N__25235\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__25235\,
            I => \N__25232\
        );

    \I__3818\ : Odrv4
    port map (
            O => \N__25232\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__3817\ : InMux
    port map (
            O => \N__25229\,
            I => \N__25226\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__25226\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__3815\ : InMux
    port map (
            O => \N__25223\,
            I => \N__25220\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__25220\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__3813\ : CascadeMux
    port map (
            O => \N__25217\,
            I => \N__25214\
        );

    \I__3812\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25211\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__25211\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__3810\ : InMux
    port map (
            O => \N__25208\,
            I => \N__25205\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__25205\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__25202\,
            I => \N__25199\
        );

    \I__3807\ : InMux
    port map (
            O => \N__25199\,
            I => \N__25196\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__25196\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__3805\ : InMux
    port map (
            O => \N__25193\,
            I => \N__25190\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__25190\,
            I => \N__25187\
        );

    \I__3803\ : Odrv12
    port map (
            O => \N__25187\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__3802\ : CascadeMux
    port map (
            O => \N__25184\,
            I => \N__25181\
        );

    \I__3801\ : InMux
    port map (
            O => \N__25181\,
            I => \N__25178\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__25178\,
            I => \N__25175\
        );

    \I__3799\ : Odrv4
    port map (
            O => \N__25175\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__3798\ : InMux
    port map (
            O => \N__25172\,
            I => \N__25169\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__25169\,
            I => \N__25166\
        );

    \I__3796\ : Span4Mux_v
    port map (
            O => \N__25166\,
            I => \N__25161\
        );

    \I__3795\ : InMux
    port map (
            O => \N__25165\,
            I => \N__25158\
        );

    \I__3794\ : InMux
    port map (
            O => \N__25164\,
            I => \N__25155\
        );

    \I__3793\ : Span4Mux_v
    port map (
            O => \N__25161\,
            I => \N__25149\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__25158\,
            I => \N__25149\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__25155\,
            I => \N__25146\
        );

    \I__3790\ : InMux
    port map (
            O => \N__25154\,
            I => \N__25143\
        );

    \I__3789\ : Span4Mux_h
    port map (
            O => \N__25149\,
            I => \N__25140\
        );

    \I__3788\ : Span12Mux_h
    port map (
            O => \N__25146\,
            I => \N__25137\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__25143\,
            I => \N__25134\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__25140\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__3785\ : Odrv12
    port map (
            O => \N__25137\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__3784\ : Odrv12
    port map (
            O => \N__25134\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__3783\ : InMux
    port map (
            O => \N__25127\,
            I => \N__25124\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__25124\,
            I => \N__25119\
        );

    \I__3781\ : InMux
    port map (
            O => \N__25123\,
            I => \N__25116\
        );

    \I__3780\ : InMux
    port map (
            O => \N__25122\,
            I => \N__25113\
        );

    \I__3779\ : Span4Mux_v
    port map (
            O => \N__25119\,
            I => \N__25108\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__25116\,
            I => \N__25108\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__25113\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__3776\ : Odrv4
    port map (
            O => \N__25108\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__3775\ : CascadeMux
    port map (
            O => \N__25103\,
            I => \N__25098\
        );

    \I__3774\ : InMux
    port map (
            O => \N__25102\,
            I => \N__25095\
        );

    \I__3773\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25092\
        );

    \I__3772\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25089\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__25095\,
            I => \N__25084\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__25092\,
            I => \N__25084\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__25089\,
            I => \N__25081\
        );

    \I__3768\ : Span4Mux_h
    port map (
            O => \N__25084\,
            I => \N__25077\
        );

    \I__3767\ : Span4Mux_v
    port map (
            O => \N__25081\,
            I => \N__25074\
        );

    \I__3766\ : InMux
    port map (
            O => \N__25080\,
            I => \N__25071\
        );

    \I__3765\ : Span4Mux_v
    port map (
            O => \N__25077\,
            I => \N__25068\
        );

    \I__3764\ : Span4Mux_h
    port map (
            O => \N__25074\,
            I => \N__25063\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__25071\,
            I => \N__25063\
        );

    \I__3762\ : Odrv4
    port map (
            O => \N__25068\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__25063\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__3760\ : InMux
    port map (
            O => \N__25058\,
            I => \N__25054\
        );

    \I__3759\ : InMux
    port map (
            O => \N__25057\,
            I => \N__25050\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__25054\,
            I => \N__25047\
        );

    \I__3757\ : InMux
    port map (
            O => \N__25053\,
            I => \N__25044\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__25050\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__3755\ : Odrv12
    port map (
            O => \N__25047\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__25044\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__3753\ : InMux
    port map (
            O => \N__25037\,
            I => \N__25028\
        );

    \I__3752\ : InMux
    port map (
            O => \N__25036\,
            I => \N__25028\
        );

    \I__3751\ : InMux
    port map (
            O => \N__25035\,
            I => \N__25028\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__25028\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__25025\,
            I => \N__25022\
        );

    \I__3748\ : InMux
    port map (
            O => \N__25022\,
            I => \N__25013\
        );

    \I__3747\ : InMux
    port map (
            O => \N__25021\,
            I => \N__25013\
        );

    \I__3746\ : InMux
    port map (
            O => \N__25020\,
            I => \N__25013\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__25013\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\
        );

    \I__3744\ : CascadeMux
    port map (
            O => \N__25010\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_\
        );

    \I__3743\ : InMux
    port map (
            O => \N__25007\,
            I => \N__25004\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__25004\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__25001\,
            I => \N__24998\
        );

    \I__3740\ : InMux
    port map (
            O => \N__24998\,
            I => \N__24995\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__24995\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__3738\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24989\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__24989\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__3736\ : CascadeMux
    port map (
            O => \N__24986\,
            I => \N__24983\
        );

    \I__3735\ : InMux
    port map (
            O => \N__24983\,
            I => \N__24980\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__24980\,
            I => \N__24977\
        );

    \I__3733\ : Odrv4
    port map (
            O => \N__24977\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__3732\ : InMux
    port map (
            O => \N__24974\,
            I => \N__24971\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__24971\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__24968\,
            I => \N__24965\
        );

    \I__3729\ : InMux
    port map (
            O => \N__24965\,
            I => \N__24962\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__24962\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__3727\ : InMux
    port map (
            O => \N__24959\,
            I => \N__24956\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__24956\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__3725\ : InMux
    port map (
            O => \N__24953\,
            I => \N__24947\
        );

    \I__3724\ : InMux
    port map (
            O => \N__24952\,
            I => \N__24947\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__24947\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\
        );

    \I__3722\ : InMux
    port map (
            O => \N__24944\,
            I => \N__24941\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__24941\,
            I => \N__24938\
        );

    \I__3720\ : Span12Mux_s11_h
    port map (
            O => \N__24938\,
            I => \N__24934\
        );

    \I__3719\ : InMux
    port map (
            O => \N__24937\,
            I => \N__24931\
        );

    \I__3718\ : Odrv12
    port map (
            O => \N__24934\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__24931\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__3716\ : CascadeMux
    port map (
            O => \N__24926\,
            I => \elapsed_time_ns_1_RNII43T9_0_6_cascade_\
        );

    \I__3715\ : InMux
    port map (
            O => \N__24923\,
            I => \N__24917\
        );

    \I__3714\ : InMux
    port map (
            O => \N__24922\,
            I => \N__24917\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__24917\,
            I => \N__24913\
        );

    \I__3712\ : InMux
    port map (
            O => \N__24916\,
            I => \N__24910\
        );

    \I__3711\ : Span4Mux_v
    port map (
            O => \N__24913\,
            I => \N__24906\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__24910\,
            I => \N__24903\
        );

    \I__3709\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24900\
        );

    \I__3708\ : Span4Mux_v
    port map (
            O => \N__24906\,
            I => \N__24895\
        );

    \I__3707\ : Span4Mux_v
    port map (
            O => \N__24903\,
            I => \N__24895\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__24900\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__3705\ : Odrv4
    port map (
            O => \N__24895\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__3704\ : InMux
    port map (
            O => \N__24890\,
            I => \N__24887\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__24887\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__3702\ : InMux
    port map (
            O => \N__24884\,
            I => \bfn_10_21_0_\
        );

    \I__3701\ : InMux
    port map (
            O => \N__24881\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__3700\ : InMux
    port map (
            O => \N__24878\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__3699\ : InMux
    port map (
            O => \N__24875\,
            I => \N__24872\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__24872\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__3697\ : InMux
    port map (
            O => \N__24869\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__3696\ : InMux
    port map (
            O => \N__24866\,
            I => \N__24863\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__24863\,
            I => \N__24860\
        );

    \I__3694\ : Span4Mux_h
    port map (
            O => \N__24860\,
            I => \N__24857\
        );

    \I__3693\ : Odrv4
    port map (
            O => \N__24857\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__3692\ : InMux
    port map (
            O => \N__24854\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__3691\ : InMux
    port map (
            O => \N__24851\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__3690\ : CascadeMux
    port map (
            O => \N__24848\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\
        );

    \I__3689\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24842\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__24842\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__3687\ : InMux
    port map (
            O => \N__24839\,
            I => \N__24836\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__24836\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__3685\ : InMux
    port map (
            O => \N__24833\,
            I => \N__24830\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__24830\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__3683\ : InMux
    port map (
            O => \N__24827\,
            I => \bfn_10_20_0_\
        );

    \I__3682\ : InMux
    port map (
            O => \N__24824\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__3681\ : CascadeMux
    port map (
            O => \N__24821\,
            I => \N__24818\
        );

    \I__3680\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24815\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__24815\,
            I => \N__24812\
        );

    \I__3678\ : Odrv4
    port map (
            O => \N__24812\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__3677\ : InMux
    port map (
            O => \N__24809\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__3676\ : InMux
    port map (
            O => \N__24806\,
            I => \N__24803\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__24803\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__3674\ : InMux
    port map (
            O => \N__24800\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__3673\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24794\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__24794\,
            I => \N__24791\
        );

    \I__3671\ : Odrv4
    port map (
            O => \N__24791\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__3670\ : InMux
    port map (
            O => \N__24788\,
            I => \N__24783\
        );

    \I__3669\ : InMux
    port map (
            O => \N__24787\,
            I => \N__24780\
        );

    \I__3668\ : InMux
    port map (
            O => \N__24786\,
            I => \N__24777\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__24783\,
            I => \N__24774\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__24780\,
            I => \N__24769\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__24777\,
            I => \N__24769\
        );

    \I__3664\ : Sp12to4
    port map (
            O => \N__24774\,
            I => \N__24766\
        );

    \I__3663\ : Span4Mux_v
    port map (
            O => \N__24769\,
            I => \N__24763\
        );

    \I__3662\ : Odrv12
    port map (
            O => \N__24766\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__3661\ : Odrv4
    port map (
            O => \N__24763\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__3660\ : InMux
    port map (
            O => \N__24758\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__3659\ : InMux
    port map (
            O => \N__24755\,
            I => \N__24752\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__24752\,
            I => \N__24749\
        );

    \I__3657\ : Span4Mux_h
    port map (
            O => \N__24749\,
            I => \N__24746\
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__24746\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__3655\ : InMux
    port map (
            O => \N__24743\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__3654\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24737\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__24737\,
            I => \N__24734\
        );

    \I__3652\ : Odrv4
    port map (
            O => \N__24734\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__3651\ : InMux
    port map (
            O => \N__24731\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__3650\ : InMux
    port map (
            O => \N__24728\,
            I => \N__24725\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__24725\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__3648\ : InMux
    port map (
            O => \N__24722\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__3647\ : InMux
    port map (
            O => \N__24719\,
            I => \N__24716\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__24716\,
            I => \N__24713\
        );

    \I__3645\ : Odrv4
    port map (
            O => \N__24713\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__3644\ : InMux
    port map (
            O => \N__24710\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__3643\ : InMux
    port map (
            O => \N__24707\,
            I => \N__24704\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__24704\,
            I => \N__24701\
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__24701\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__3640\ : InMux
    port map (
            O => \N__24698\,
            I => \N__24693\
        );

    \I__3639\ : InMux
    port map (
            O => \N__24697\,
            I => \N__24690\
        );

    \I__3638\ : InMux
    port map (
            O => \N__24696\,
            I => \N__24687\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__24693\,
            I => \N__24684\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__24690\,
            I => \N__24679\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__24687\,
            I => \N__24679\
        );

    \I__3634\ : Odrv12
    port map (
            O => \N__24684\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__3633\ : Odrv12
    port map (
            O => \N__24679\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__3632\ : InMux
    port map (
            O => \N__24674\,
            I => \bfn_10_19_0_\
        );

    \I__3631\ : InMux
    port map (
            O => \N__24671\,
            I => \N__24668\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__24668\,
            I => \N__24665\
        );

    \I__3629\ : Odrv4
    port map (
            O => \N__24665\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__3628\ : InMux
    port map (
            O => \N__24662\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__3627\ : InMux
    port map (
            O => \N__24659\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__3626\ : InMux
    port map (
            O => \N__24656\,
            I => \N__24653\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__24653\,
            I => \N__24650\
        );

    \I__3624\ : Odrv12
    port map (
            O => \N__24650\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__3623\ : InMux
    port map (
            O => \N__24647\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__3622\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24641\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__24641\,
            I => \N__24638\
        );

    \I__3620\ : Odrv4
    port map (
            O => \N__24638\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__3619\ : InMux
    port map (
            O => \N__24635\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__3618\ : InMux
    port map (
            O => \N__24632\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__3617\ : InMux
    port map (
            O => \N__24629\,
            I => \N__24626\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__24626\,
            I => \N__24623\
        );

    \I__3615\ : Odrv12
    port map (
            O => \N__24623\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__3614\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24615\
        );

    \I__3613\ : InMux
    port map (
            O => \N__24619\,
            I => \N__24610\
        );

    \I__3612\ : InMux
    port map (
            O => \N__24618\,
            I => \N__24610\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__24615\,
            I => \N__24605\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__24610\,
            I => \N__24605\
        );

    \I__3609\ : Odrv12
    port map (
            O => \N__24605\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__3608\ : InMux
    port map (
            O => \N__24602\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__3607\ : InMux
    port map (
            O => \N__24599\,
            I => \N__24596\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__24596\,
            I => \N__24593\
        );

    \I__3605\ : Odrv12
    port map (
            O => \N__24593\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__3604\ : InMux
    port map (
            O => \N__24590\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__24587\,
            I => \N__24584\
        );

    \I__3602\ : InMux
    port map (
            O => \N__24584\,
            I => \N__24581\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__24581\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__3600\ : InMux
    port map (
            O => \N__24578\,
            I => \N__24575\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__24575\,
            I => \N__24572\
        );

    \I__3598\ : Odrv12
    port map (
            O => \N__24572\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__3597\ : InMux
    port map (
            O => \N__24569\,
            I => \N__24560\
        );

    \I__3596\ : InMux
    port map (
            O => \N__24568\,
            I => \N__24560\
        );

    \I__3595\ : InMux
    port map (
            O => \N__24567\,
            I => \N__24560\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__24560\,
            I => \N__24557\
        );

    \I__3593\ : Odrv12
    port map (
            O => \N__24557\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__3592\ : InMux
    port map (
            O => \N__24554\,
            I => \N__24551\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__24551\,
            I => \N__24548\
        );

    \I__3590\ : Span4Mux_h
    port map (
            O => \N__24548\,
            I => \N__24545\
        );

    \I__3589\ : Odrv4
    port map (
            O => \N__24545\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__3588\ : InMux
    port map (
            O => \N__24542\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__3587\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__24536\,
            I => \N__24533\
        );

    \I__3585\ : Span4Mux_h
    port map (
            O => \N__24533\,
            I => \N__24530\
        );

    \I__3584\ : Odrv4
    port map (
            O => \N__24530\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__3583\ : InMux
    port map (
            O => \N__24527\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__3582\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24521\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__24521\,
            I => \N__24518\
        );

    \I__3580\ : Span4Mux_v
    port map (
            O => \N__24518\,
            I => \N__24515\
        );

    \I__3579\ : Odrv4
    port map (
            O => \N__24515\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__3578\ : InMux
    port map (
            O => \N__24512\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__3577\ : InMux
    port map (
            O => \N__24509\,
            I => \N__24506\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__24506\,
            I => \N__24503\
        );

    \I__3575\ : Odrv12
    port map (
            O => \N__24503\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__24500\,
            I => \N__24496\
        );

    \I__3573\ : CascadeMux
    port map (
            O => \N__24499\,
            I => \N__24493\
        );

    \I__3572\ : InMux
    port map (
            O => \N__24496\,
            I => \N__24490\
        );

    \I__3571\ : InMux
    port map (
            O => \N__24493\,
            I => \N__24487\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__24490\,
            I => \N__24484\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__24487\,
            I => \N__24478\
        );

    \I__3568\ : Span4Mux_v
    port map (
            O => \N__24484\,
            I => \N__24478\
        );

    \I__3567\ : InMux
    port map (
            O => \N__24483\,
            I => \N__24475\
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__24478\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__24475\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__3564\ : InMux
    port map (
            O => \N__24470\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__3563\ : InMux
    port map (
            O => \N__24467\,
            I => \N__24464\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__24464\,
            I => \N__24461\
        );

    \I__3561\ : Span4Mux_h
    port map (
            O => \N__24461\,
            I => \N__24458\
        );

    \I__3560\ : Odrv4
    port map (
            O => \N__24458\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__3559\ : InMux
    port map (
            O => \N__24455\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__3558\ : InMux
    port map (
            O => \N__24452\,
            I => \N__24449\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__24449\,
            I => \N__24446\
        );

    \I__3556\ : Odrv12
    port map (
            O => \N__24446\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__3555\ : InMux
    port map (
            O => \N__24443\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__3554\ : InMux
    port map (
            O => \N__24440\,
            I => \N__24437\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__24437\,
            I => \N__24432\
        );

    \I__3552\ : InMux
    port map (
            O => \N__24436\,
            I => \N__24427\
        );

    \I__3551\ : InMux
    port map (
            O => \N__24435\,
            I => \N__24427\
        );

    \I__3550\ : Span4Mux_v
    port map (
            O => \N__24432\,
            I => \N__24422\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__24427\,
            I => \N__24422\
        );

    \I__3548\ : Span4Mux_h
    port map (
            O => \N__24422\,
            I => \N__24418\
        );

    \I__3547\ : InMux
    port map (
            O => \N__24421\,
            I => \N__24415\
        );

    \I__3546\ : Span4Mux_v
    port map (
            O => \N__24418\,
            I => \N__24412\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__24415\,
            I => \N__24409\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__24412\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__24409\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__24404\,
            I => \N__24401\
        );

    \I__3541\ : InMux
    port map (
            O => \N__24401\,
            I => \N__24398\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__24398\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__3539\ : InMux
    port map (
            O => \N__24395\,
            I => \N__24391\
        );

    \I__3538\ : InMux
    port map (
            O => \N__24394\,
            I => \N__24388\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__24391\,
            I => \N__24382\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__24388\,
            I => \N__24382\
        );

    \I__3535\ : InMux
    port map (
            O => \N__24387\,
            I => \N__24379\
        );

    \I__3534\ : Span4Mux_v
    port map (
            O => \N__24382\,
            I => \N__24375\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__24379\,
            I => \N__24372\
        );

    \I__3532\ : InMux
    port map (
            O => \N__24378\,
            I => \N__24369\
        );

    \I__3531\ : Span4Mux_h
    port map (
            O => \N__24375\,
            I => \N__24366\
        );

    \I__3530\ : Span4Mux_h
    port map (
            O => \N__24372\,
            I => \N__24361\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__24369\,
            I => \N__24361\
        );

    \I__3528\ : Odrv4
    port map (
            O => \N__24366\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__3527\ : Odrv4
    port map (
            O => \N__24361\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__24356\,
            I => \N__24353\
        );

    \I__3525\ : InMux
    port map (
            O => \N__24353\,
            I => \N__24350\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__24350\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__24347\,
            I => \N__24344\
        );

    \I__3522\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24341\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__24341\,
            I => \N__24338\
        );

    \I__3520\ : Odrv4
    port map (
            O => \N__24338\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__3519\ : CascadeMux
    port map (
            O => \N__24335\,
            I => \N__24332\
        );

    \I__3518\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24329\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__24329\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__3516\ : InMux
    port map (
            O => \N__24326\,
            I => \N__24323\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__24323\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__3514\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24317\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__24317\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__3512\ : InMux
    port map (
            O => \N__24314\,
            I => \N__24311\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__24311\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__3510\ : CascadeMux
    port map (
            O => \N__24308\,
            I => \N__24305\
        );

    \I__3509\ : InMux
    port map (
            O => \N__24305\,
            I => \N__24302\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__24302\,
            I => \N__24299\
        );

    \I__3507\ : Span4Mux_v
    port map (
            O => \N__24299\,
            I => \N__24296\
        );

    \I__3506\ : Odrv4
    port map (
            O => \N__24296\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__3505\ : InMux
    port map (
            O => \N__24293\,
            I => \N__24290\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__24290\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__24287\,
            I => \current_shift_inst.control_input_axb_0_cascade_\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__24284\,
            I => \N__24279\
        );

    \I__3501\ : InMux
    port map (
            O => \N__24283\,
            I => \N__24276\
        );

    \I__3500\ : InMux
    port map (
            O => \N__24282\,
            I => \N__24273\
        );

    \I__3499\ : InMux
    port map (
            O => \N__24279\,
            I => \N__24270\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__24276\,
            I => \current_shift_inst.N_1288_i\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__24273\,
            I => \current_shift_inst.N_1288_i\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__24270\,
            I => \current_shift_inst.N_1288_i\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__24263\,
            I => \N__24259\
        );

    \I__3494\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24256\
        );

    \I__3493\ : InMux
    port map (
            O => \N__24259\,
            I => \N__24253\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__24256\,
            I => \N__24250\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__24253\,
            I => \N__24246\
        );

    \I__3490\ : Span4Mux_v
    port map (
            O => \N__24250\,
            I => \N__24243\
        );

    \I__3489\ : InMux
    port map (
            O => \N__24249\,
            I => \N__24240\
        );

    \I__3488\ : Span4Mux_h
    port map (
            O => \N__24246\,
            I => \N__24237\
        );

    \I__3487\ : Sp12to4
    port map (
            O => \N__24243\,
            I => \N__24232\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__24240\,
            I => \N__24232\
        );

    \I__3485\ : Span4Mux_v
    port map (
            O => \N__24237\,
            I => \N__24228\
        );

    \I__3484\ : Span12Mux_h
    port map (
            O => \N__24232\,
            I => \N__24225\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24231\,
            I => \N__24222\
        );

    \I__3482\ : Odrv4
    port map (
            O => \N__24228\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__3481\ : Odrv12
    port map (
            O => \N__24225\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__24222\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__3479\ : CascadeMux
    port map (
            O => \N__24215\,
            I => \N__24212\
        );

    \I__3478\ : InMux
    port map (
            O => \N__24212\,
            I => \N__24209\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__24209\,
            I => \N__24206\
        );

    \I__3476\ : Span4Mux_v
    port map (
            O => \N__24206\,
            I => \N__24203\
        );

    \I__3475\ : Span4Mux_h
    port map (
            O => \N__24203\,
            I => \N__24200\
        );

    \I__3474\ : Odrv4
    port map (
            O => \N__24200\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__3473\ : InMux
    port map (
            O => \N__24197\,
            I => \N__24194\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__24194\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt26\
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__24191\,
            I => \N__24188\
        );

    \I__3470\ : InMux
    port map (
            O => \N__24188\,
            I => \N__24178\
        );

    \I__3469\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24178\
        );

    \I__3468\ : InMux
    port map (
            O => \N__24186\,
            I => \N__24178\
        );

    \I__3467\ : InMux
    port map (
            O => \N__24185\,
            I => \N__24175\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__24178\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__24175\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__3464\ : InMux
    port map (
            O => \N__24170\,
            I => \N__24167\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__24167\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__3462\ : CascadeMux
    port map (
            O => \N__24164\,
            I => \N__24161\
        );

    \I__3461\ : InMux
    port map (
            O => \N__24161\,
            I => \N__24158\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__24158\,
            I => \N__24155\
        );

    \I__3459\ : Odrv4
    port map (
            O => \N__24155\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt16\
        );

    \I__3458\ : InMux
    port map (
            O => \N__24152\,
            I => \N__24149\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__24149\,
            I => \N__24144\
        );

    \I__3456\ : InMux
    port map (
            O => \N__24148\,
            I => \N__24139\
        );

    \I__3455\ : InMux
    port map (
            O => \N__24147\,
            I => \N__24139\
        );

    \I__3454\ : Span4Mux_v
    port map (
            O => \N__24144\,
            I => \N__24136\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__24139\,
            I => \N__24132\
        );

    \I__3452\ : Span4Mux_v
    port map (
            O => \N__24136\,
            I => \N__24129\
        );

    \I__3451\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24126\
        );

    \I__3450\ : Span4Mux_v
    port map (
            O => \N__24132\,
            I => \N__24123\
        );

    \I__3449\ : Span4Mux_v
    port map (
            O => \N__24129\,
            I => \N__24118\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__24126\,
            I => \N__24118\
        );

    \I__3447\ : Odrv4
    port map (
            O => \N__24123\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__24118\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__3445\ : InMux
    port map (
            O => \N__24113\,
            I => \N__24110\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__24110\,
            I => \N__24107\
        );

    \I__3443\ : Span4Mux_v
    port map (
            O => \N__24107\,
            I => \N__24104\
        );

    \I__3442\ : Span4Mux_v
    port map (
            O => \N__24104\,
            I => \N__24101\
        );

    \I__3441\ : Odrv4
    port map (
            O => \N__24101\,
            I => \il_min_comp1_D1\
        );

    \I__3440\ : InMux
    port map (
            O => \N__24098\,
            I => \N__24092\
        );

    \I__3439\ : InMux
    port map (
            O => \N__24097\,
            I => \N__24092\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__24092\,
            I => \N__24089\
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__24089\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__24086\,
            I => \N__24082\
        );

    \I__3435\ : CascadeMux
    port map (
            O => \N__24085\,
            I => \N__24079\
        );

    \I__3434\ : InMux
    port map (
            O => \N__24082\,
            I => \N__24074\
        );

    \I__3433\ : InMux
    port map (
            O => \N__24079\,
            I => \N__24074\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__24074\,
            I => \N__24071\
        );

    \I__3431\ : Odrv4
    port map (
            O => \N__24071\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__3430\ : InMux
    port map (
            O => \N__24068\,
            I => \N__24065\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__24065\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\
        );

    \I__3428\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24059\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__24059\,
            I => \N__24054\
        );

    \I__3426\ : InMux
    port map (
            O => \N__24058\,
            I => \N__24051\
        );

    \I__3425\ : InMux
    port map (
            O => \N__24057\,
            I => \N__24048\
        );

    \I__3424\ : Span4Mux_v
    port map (
            O => \N__24054\,
            I => \N__24043\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__24051\,
            I => \N__24043\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__24048\,
            I => \N__24037\
        );

    \I__3421\ : Span4Mux_h
    port map (
            O => \N__24043\,
            I => \N__24037\
        );

    \I__3420\ : InMux
    port map (
            O => \N__24042\,
            I => \N__24034\
        );

    \I__3419\ : Span4Mux_v
    port map (
            O => \N__24037\,
            I => \N__24029\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__24034\,
            I => \N__24029\
        );

    \I__3417\ : Span4Mux_v
    port map (
            O => \N__24029\,
            I => \N__24026\
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__24026\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__3415\ : InMux
    port map (
            O => \N__24023\,
            I => \N__24018\
        );

    \I__3414\ : InMux
    port map (
            O => \N__24022\,
            I => \N__24015\
        );

    \I__3413\ : InMux
    port map (
            O => \N__24021\,
            I => \N__24012\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__24018\,
            I => \N__24009\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__24015\,
            I => \N__24006\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__24012\,
            I => \N__24000\
        );

    \I__3409\ : Span4Mux_h
    port map (
            O => \N__24009\,
            I => \N__24000\
        );

    \I__3408\ : Span4Mux_v
    port map (
            O => \N__24006\,
            I => \N__23997\
        );

    \I__3407\ : InMux
    port map (
            O => \N__24005\,
            I => \N__23994\
        );

    \I__3406\ : Span4Mux_v
    port map (
            O => \N__24000\,
            I => \N__23991\
        );

    \I__3405\ : Span4Mux_v
    port map (
            O => \N__23997\,
            I => \N__23986\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__23994\,
            I => \N__23986\
        );

    \I__3403\ : Odrv4
    port map (
            O => \N__23991\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__23986\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__3401\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23978\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__23978\,
            I => \N__23975\
        );

    \I__3399\ : Span4Mux_h
    port map (
            O => \N__23975\,
            I => \N__23972\
        );

    \I__3398\ : Span4Mux_v
    port map (
            O => \N__23972\,
            I => \N__23969\
        );

    \I__3397\ : Odrv4
    port map (
            O => \N__23969\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\
        );

    \I__3396\ : InMux
    port map (
            O => \N__23966\,
            I => \N__23963\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__23963\,
            I => \N__23960\
        );

    \I__3394\ : Span4Mux_v
    port map (
            O => \N__23960\,
            I => \N__23957\
        );

    \I__3393\ : Span4Mux_v
    port map (
            O => \N__23957\,
            I => \N__23952\
        );

    \I__3392\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23949\
        );

    \I__3391\ : InMux
    port map (
            O => \N__23955\,
            I => \N__23946\
        );

    \I__3390\ : Odrv4
    port map (
            O => \N__23952\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__23949\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__23946\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__3387\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23934\
        );

    \I__3386\ : InMux
    port map (
            O => \N__23938\,
            I => \N__23930\
        );

    \I__3385\ : InMux
    port map (
            O => \N__23937\,
            I => \N__23927\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__23934\,
            I => \N__23924\
        );

    \I__3383\ : InMux
    port map (
            O => \N__23933\,
            I => \N__23921\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__23930\,
            I => \N__23918\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__23927\,
            I => \N__23915\
        );

    \I__3380\ : Span4Mux_h
    port map (
            O => \N__23924\,
            I => \N__23912\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__23921\,
            I => \N__23909\
        );

    \I__3378\ : Span4Mux_v
    port map (
            O => \N__23918\,
            I => \N__23904\
        );

    \I__3377\ : Span4Mux_h
    port map (
            O => \N__23915\,
            I => \N__23904\
        );

    \I__3376\ : Span4Mux_v
    port map (
            O => \N__23912\,
            I => \N__23899\
        );

    \I__3375\ : Span4Mux_h
    port map (
            O => \N__23909\,
            I => \N__23899\
        );

    \I__3374\ : Span4Mux_v
    port map (
            O => \N__23904\,
            I => \N__23896\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__23899\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__3372\ : Odrv4
    port map (
            O => \N__23896\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__3371\ : InMux
    port map (
            O => \N__23891\,
            I => \N__23888\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__23888\,
            I => \N__23885\
        );

    \I__3369\ : Span4Mux_v
    port map (
            O => \N__23885\,
            I => \N__23880\
        );

    \I__3368\ : InMux
    port map (
            O => \N__23884\,
            I => \N__23877\
        );

    \I__3367\ : InMux
    port map (
            O => \N__23883\,
            I => \N__23874\
        );

    \I__3366\ : Sp12to4
    port map (
            O => \N__23880\,
            I => \N__23869\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__23877\,
            I => \N__23869\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__23874\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__3363\ : Odrv12
    port map (
            O => \N__23869\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__3362\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23860\
        );

    \I__3361\ : InMux
    port map (
            O => \N__23863\,
            I => \N__23857\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__23860\,
            I => \N__23853\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__23857\,
            I => \N__23849\
        );

    \I__3358\ : InMux
    port map (
            O => \N__23856\,
            I => \N__23846\
        );

    \I__3357\ : Span4Mux_v
    port map (
            O => \N__23853\,
            I => \N__23843\
        );

    \I__3356\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23840\
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__23849\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__23846\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__23843\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__23840\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__3351\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23828\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__23828\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__3349\ : CascadeMux
    port map (
            O => \N__23825\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df30_cascade_\
        );

    \I__3348\ : InMux
    port map (
            O => \N__23822\,
            I => \N__23819\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__23819\,
            I => \N__23816\
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__23816\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__23813\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__23810\,
            I => \N__23807\
        );

    \I__3343\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23804\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__23804\,
            I => \N__23801\
        );

    \I__3341\ : Span4Mux_v
    port map (
            O => \N__23801\,
            I => \N__23797\
        );

    \I__3340\ : InMux
    port map (
            O => \N__23800\,
            I => \N__23794\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__23797\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt30\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__23794\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt30\
        );

    \I__3337\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23780\
        );

    \I__3336\ : InMux
    port map (
            O => \N__23788\,
            I => \N__23780\
        );

    \I__3335\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23780\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__23780\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\
        );

    \I__3333\ : InMux
    port map (
            O => \N__23777\,
            I => \N__23768\
        );

    \I__3332\ : InMux
    port map (
            O => \N__23776\,
            I => \N__23768\
        );

    \I__3331\ : InMux
    port map (
            O => \N__23775\,
            I => \N__23768\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__23768\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\
        );

    \I__3329\ : InMux
    port map (
            O => \N__23765\,
            I => \N__23762\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__23762\,
            I => \N__23759\
        );

    \I__3327\ : Odrv4
    port map (
            O => \N__23759\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\
        );

    \I__3326\ : CascadeMux
    port map (
            O => \N__23756\,
            I => \N__23753\
        );

    \I__3325\ : InMux
    port map (
            O => \N__23753\,
            I => \N__23749\
        );

    \I__3324\ : InMux
    port map (
            O => \N__23752\,
            I => \N__23746\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__23749\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__23746\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__3321\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23738\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__23738\,
            I => \N__23733\
        );

    \I__3319\ : InMux
    port map (
            O => \N__23737\,
            I => \N__23730\
        );

    \I__3318\ : InMux
    port map (
            O => \N__23736\,
            I => \N__23727\
        );

    \I__3317\ : Span4Mux_v
    port map (
            O => \N__23733\,
            I => \N__23724\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__23730\,
            I => \N__23721\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__23727\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__3314\ : Odrv4
    port map (
            O => \N__23724\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__3313\ : Odrv12
    port map (
            O => \N__23721\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__3312\ : InMux
    port map (
            O => \N__23714\,
            I => \N__23710\
        );

    \I__3311\ : InMux
    port map (
            O => \N__23713\,
            I => \N__23707\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__23710\,
            I => \N__23704\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__23707\,
            I => \N__23700\
        );

    \I__3308\ : Span4Mux_h
    port map (
            O => \N__23704\,
            I => \N__23696\
        );

    \I__3307\ : InMux
    port map (
            O => \N__23703\,
            I => \N__23693\
        );

    \I__3306\ : Span4Mux_h
    port map (
            O => \N__23700\,
            I => \N__23690\
        );

    \I__3305\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23687\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__23696\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__23693\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__3302\ : Odrv4
    port map (
            O => \N__23690\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__23687\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__3300\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23674\
        );

    \I__3299\ : InMux
    port map (
            O => \N__23677\,
            I => \N__23671\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__23674\,
            I => \N__23667\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__23671\,
            I => \N__23664\
        );

    \I__3296\ : InMux
    port map (
            O => \N__23670\,
            I => \N__23661\
        );

    \I__3295\ : Span4Mux_v
    port map (
            O => \N__23667\,
            I => \N__23656\
        );

    \I__3294\ : Span4Mux_h
    port map (
            O => \N__23664\,
            I => \N__23656\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__23661\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__3292\ : Odrv4
    port map (
            O => \N__23656\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__3291\ : InMux
    port map (
            O => \N__23651\,
            I => \N__23647\
        );

    \I__3290\ : InMux
    port map (
            O => \N__23650\,
            I => \N__23644\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__23647\,
            I => \N__23640\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__23644\,
            I => \N__23637\
        );

    \I__3287\ : InMux
    port map (
            O => \N__23643\,
            I => \N__23633\
        );

    \I__3286\ : Span4Mux_h
    port map (
            O => \N__23640\,
            I => \N__23628\
        );

    \I__3285\ : Span4Mux_h
    port map (
            O => \N__23637\,
            I => \N__23628\
        );

    \I__3284\ : InMux
    port map (
            O => \N__23636\,
            I => \N__23625\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__23633\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__3282\ : Odrv4
    port map (
            O => \N__23628\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__23625\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__3280\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__3278\ : Span4Mux_h
    port map (
            O => \N__23612\,
            I => \N__23607\
        );

    \I__3277\ : InMux
    port map (
            O => \N__23611\,
            I => \N__23604\
        );

    \I__3276\ : InMux
    port map (
            O => \N__23610\,
            I => \N__23601\
        );

    \I__3275\ : Span4Mux_h
    port map (
            O => \N__23607\,
            I => \N__23598\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__23604\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__23601\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__3272\ : Odrv4
    port map (
            O => \N__23598\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__3271\ : InMux
    port map (
            O => \N__23591\,
            I => \N__23586\
        );

    \I__3270\ : InMux
    port map (
            O => \N__23590\,
            I => \N__23583\
        );

    \I__3269\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23580\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__23586\,
            I => \N__23576\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__23583\,
            I => \N__23571\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__23580\,
            I => \N__23571\
        );

    \I__3265\ : InMux
    port map (
            O => \N__23579\,
            I => \N__23568\
        );

    \I__3264\ : Span4Mux_v
    port map (
            O => \N__23576\,
            I => \N__23565\
        );

    \I__3263\ : Span4Mux_v
    port map (
            O => \N__23571\,
            I => \N__23562\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__23568\,
            I => \N__23559\
        );

    \I__3261\ : Span4Mux_v
    port map (
            O => \N__23565\,
            I => \N__23556\
        );

    \I__3260\ : Span4Mux_h
    port map (
            O => \N__23562\,
            I => \N__23551\
        );

    \I__3259\ : Span4Mux_v
    port map (
            O => \N__23559\,
            I => \N__23551\
        );

    \I__3258\ : Odrv4
    port map (
            O => \N__23556\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__3257\ : Odrv4
    port map (
            O => \N__23551\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__23546\,
            I => \N__23543\
        );

    \I__3255\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23537\
        );

    \I__3254\ : InMux
    port map (
            O => \N__23542\,
            I => \N__23537\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__23537\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\
        );

    \I__3252\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23529\
        );

    \I__3251\ : InMux
    port map (
            O => \N__23533\,
            I => \N__23526\
        );

    \I__3250\ : InMux
    port map (
            O => \N__23532\,
            I => \N__23523\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__23529\,
            I => \N__23520\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__23526\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__23523\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__3246\ : Odrv4
    port map (
            O => \N__23520\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__3245\ : InMux
    port map (
            O => \N__23513\,
            I => \N__23507\
        );

    \I__3244\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23504\
        );

    \I__3243\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23499\
        );

    \I__3242\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23499\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__23507\,
            I => \N__23496\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__23504\,
            I => \N__23493\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__23499\,
            I => \N__23490\
        );

    \I__3238\ : Span4Mux_v
    port map (
            O => \N__23496\,
            I => \N__23487\
        );

    \I__3237\ : Span4Mux_v
    port map (
            O => \N__23493\,
            I => \N__23484\
        );

    \I__3236\ : Span4Mux_h
    port map (
            O => \N__23490\,
            I => \N__23481\
        );

    \I__3235\ : Odrv4
    port map (
            O => \N__23487\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__3234\ : Odrv4
    port map (
            O => \N__23484\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__3233\ : Odrv4
    port map (
            O => \N__23481\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__3232\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23471\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__23471\,
            I => \N__23468\
        );

    \I__3230\ : Odrv4
    port map (
            O => \N__23468\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__3229\ : InMux
    port map (
            O => \N__23465\,
            I => \N__23460\
        );

    \I__3228\ : InMux
    port map (
            O => \N__23464\,
            I => \N__23457\
        );

    \I__3227\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23454\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__23460\,
            I => \N__23449\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__23457\,
            I => \N__23449\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__23454\,
            I => \N__23446\
        );

    \I__3223\ : Odrv4
    port map (
            O => \N__23449\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__3222\ : Odrv4
    port map (
            O => \N__23446\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__3221\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23436\
        );

    \I__3220\ : InMux
    port map (
            O => \N__23440\,
            I => \N__23433\
        );

    \I__3219\ : CascadeMux
    port map (
            O => \N__23439\,
            I => \N__23429\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__23436\,
            I => \N__23426\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__23433\,
            I => \N__23423\
        );

    \I__3216\ : InMux
    port map (
            O => \N__23432\,
            I => \N__23420\
        );

    \I__3215\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23417\
        );

    \I__3214\ : Span4Mux_h
    port map (
            O => \N__23426\,
            I => \N__23412\
        );

    \I__3213\ : Span4Mux_h
    port map (
            O => \N__23423\,
            I => \N__23412\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__23420\,
            I => \N__23409\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__23417\,
            I => \N__23406\
        );

    \I__3210\ : Span4Mux_v
    port map (
            O => \N__23412\,
            I => \N__23403\
        );

    \I__3209\ : Span4Mux_v
    port map (
            O => \N__23409\,
            I => \N__23400\
        );

    \I__3208\ : Span4Mux_h
    port map (
            O => \N__23406\,
            I => \N__23397\
        );

    \I__3207\ : Span4Mux_v
    port map (
            O => \N__23403\,
            I => \N__23392\
        );

    \I__3206\ : Span4Mux_v
    port map (
            O => \N__23400\,
            I => \N__23392\
        );

    \I__3205\ : Span4Mux_v
    port map (
            O => \N__23397\,
            I => \N__23389\
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__23392\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__23389\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__3202\ : InMux
    port map (
            O => \N__23384\,
            I => \N__23381\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__23381\,
            I => \N__23376\
        );

    \I__3200\ : InMux
    port map (
            O => \N__23380\,
            I => \N__23373\
        );

    \I__3199\ : InMux
    port map (
            O => \N__23379\,
            I => \N__23370\
        );

    \I__3198\ : Span4Mux_v
    port map (
            O => \N__23376\,
            I => \N__23365\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__23373\,
            I => \N__23365\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__23370\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__3195\ : Odrv4
    port map (
            O => \N__23365\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__3194\ : InMux
    port map (
            O => \N__23360\,
            I => \N__23354\
        );

    \I__3193\ : InMux
    port map (
            O => \N__23359\,
            I => \N__23354\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__23354\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__23351\,
            I => \N__23347\
        );

    \I__3190\ : InMux
    port map (
            O => \N__23350\,
            I => \N__23342\
        );

    \I__3189\ : InMux
    port map (
            O => \N__23347\,
            I => \N__23342\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__23342\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__3187\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23336\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__23336\,
            I => \N__23332\
        );

    \I__3185\ : InMux
    port map (
            O => \N__23335\,
            I => \N__23329\
        );

    \I__3184\ : Odrv4
    port map (
            O => \N__23332\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__23329\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\
        );

    \I__3182\ : InMux
    port map (
            O => \N__23324\,
            I => \N__23321\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__23321\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__23318\,
            I => \N__23315\
        );

    \I__3179\ : InMux
    port map (
            O => \N__23315\,
            I => \N__23312\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__23312\,
            I => \N__23309\
        );

    \I__3177\ : Span4Mux_h
    port map (
            O => \N__23309\,
            I => \N__23306\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__23306\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\
        );

    \I__3175\ : InMux
    port map (
            O => \N__23303\,
            I => \N__23300\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__23300\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__23297\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\
        );

    \I__3172\ : InMux
    port map (
            O => \N__23294\,
            I => \N__23289\
        );

    \I__3171\ : InMux
    port map (
            O => \N__23293\,
            I => \N__23286\
        );

    \I__3170\ : InMux
    port map (
            O => \N__23292\,
            I => \N__23283\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__23289\,
            I => \N__23277\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__23286\,
            I => \N__23277\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__23283\,
            I => \N__23274\
        );

    \I__3166\ : InMux
    port map (
            O => \N__23282\,
            I => \N__23271\
        );

    \I__3165\ : Span4Mux_s3_v
    port map (
            O => \N__23277\,
            I => \N__23268\
        );

    \I__3164\ : Span4Mux_s3_v
    port map (
            O => \N__23274\,
            I => \N__23265\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__23271\,
            I => \N__23262\
        );

    \I__3162\ : Span4Mux_v
    port map (
            O => \N__23268\,
            I => \N__23259\
        );

    \I__3161\ : Span4Mux_v
    port map (
            O => \N__23265\,
            I => \N__23254\
        );

    \I__3160\ : Span4Mux_h
    port map (
            O => \N__23262\,
            I => \N__23254\
        );

    \I__3159\ : Odrv4
    port map (
            O => \N__23259\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__3158\ : Odrv4
    port map (
            O => \N__23254\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__3157\ : InMux
    port map (
            O => \N__23249\,
            I => \N__23246\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__23246\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\
        );

    \I__3155\ : InMux
    port map (
            O => \N__23243\,
            I => \N__23240\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__23240\,
            I => \N__23236\
        );

    \I__3153\ : InMux
    port map (
            O => \N__23239\,
            I => \N__23231\
        );

    \I__3152\ : Span4Mux_h
    port map (
            O => \N__23236\,
            I => \N__23228\
        );

    \I__3151\ : InMux
    port map (
            O => \N__23235\,
            I => \N__23223\
        );

    \I__3150\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23223\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__23231\,
            I => \N__23220\
        );

    \I__3148\ : Odrv4
    port map (
            O => \N__23228\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__23223\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__3146\ : Odrv4
    port map (
            O => \N__23220\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__3145\ : InMux
    port map (
            O => \N__23213\,
            I => \N__23209\
        );

    \I__3144\ : InMux
    port map (
            O => \N__23212\,
            I => \N__23206\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__23209\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__23206\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__23201\,
            I => \N__23198\
        );

    \I__3140\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23194\
        );

    \I__3139\ : InMux
    port map (
            O => \N__23197\,
            I => \N__23191\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__23194\,
            I => \N__23188\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__23191\,
            I => \N__23185\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__23188\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\
        );

    \I__3135\ : Odrv12
    port map (
            O => \N__23185\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23175\
        );

    \I__3133\ : InMux
    port map (
            O => \N__23179\,
            I => \N__23172\
        );

    \I__3132\ : InMux
    port map (
            O => \N__23178\,
            I => \N__23169\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__23175\,
            I => \N__23166\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__23172\,
            I => \N__23163\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__23169\,
            I => \N__23159\
        );

    \I__3128\ : Span4Mux_v
    port map (
            O => \N__23166\,
            I => \N__23154\
        );

    \I__3127\ : Span4Mux_v
    port map (
            O => \N__23163\,
            I => \N__23154\
        );

    \I__3126\ : InMux
    port map (
            O => \N__23162\,
            I => \N__23151\
        );

    \I__3125\ : Span4Mux_v
    port map (
            O => \N__23159\,
            I => \N__23148\
        );

    \I__3124\ : Span4Mux_v
    port map (
            O => \N__23154\,
            I => \N__23145\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__23151\,
            I => \N__23142\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__23148\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__23145\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__3120\ : Odrv4
    port map (
            O => \N__23142\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__3119\ : InMux
    port map (
            O => \N__23135\,
            I => \N__23130\
        );

    \I__3118\ : InMux
    port map (
            O => \N__23134\,
            I => \N__23127\
        );

    \I__3117\ : InMux
    port map (
            O => \N__23133\,
            I => \N__23124\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__23130\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__23127\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__23124\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__3113\ : InMux
    port map (
            O => \N__23117\,
            I => \N__23112\
        );

    \I__3112\ : InMux
    port map (
            O => \N__23116\,
            I => \N__23109\
        );

    \I__3111\ : InMux
    port map (
            O => \N__23115\,
            I => \N__23106\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__23112\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__23109\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__23106\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__3107\ : InMux
    port map (
            O => \N__23099\,
            I => \N__23094\
        );

    \I__3106\ : CascadeMux
    port map (
            O => \N__23098\,
            I => \N__23090\
        );

    \I__3105\ : InMux
    port map (
            O => \N__23097\,
            I => \N__23087\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__23094\,
            I => \N__23084\
        );

    \I__3103\ : InMux
    port map (
            O => \N__23093\,
            I => \N__23081\
        );

    \I__3102\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23078\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__23087\,
            I => \N__23069\
        );

    \I__3100\ : Span4Mux_h
    port map (
            O => \N__23084\,
            I => \N__23069\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__23081\,
            I => \N__23069\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__23078\,
            I => \N__23069\
        );

    \I__3097\ : Odrv4
    port map (
            O => \N__23069\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__3096\ : InMux
    port map (
            O => \N__23066\,
            I => \N__23061\
        );

    \I__3095\ : InMux
    port map (
            O => \N__23065\,
            I => \N__23058\
        );

    \I__3094\ : InMux
    port map (
            O => \N__23064\,
            I => \N__23055\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__23061\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__23058\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__23055\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__3090\ : CascadeMux
    port map (
            O => \N__23048\,
            I => \N__23045\
        );

    \I__3089\ : InMux
    port map (
            O => \N__23045\,
            I => \N__23042\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__23042\,
            I => \N__23036\
        );

    \I__3087\ : InMux
    port map (
            O => \N__23041\,
            I => \N__23033\
        );

    \I__3086\ : InMux
    port map (
            O => \N__23040\,
            I => \N__23028\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23039\,
            I => \N__23028\
        );

    \I__3084\ : Odrv4
    port map (
            O => \N__23036\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__23033\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__23028\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__3081\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23016\
        );

    \I__3080\ : InMux
    port map (
            O => \N__23020\,
            I => \N__23013\
        );

    \I__3079\ : InMux
    port map (
            O => \N__23019\,
            I => \N__23010\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__23016\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__23013\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__23010\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__3075\ : InMux
    port map (
            O => \N__23003\,
            I => \N__23000\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__23000\,
            I => \N__22994\
        );

    \I__3073\ : InMux
    port map (
            O => \N__22999\,
            I => \N__22991\
        );

    \I__3072\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22986\
        );

    \I__3071\ : InMux
    port map (
            O => \N__22997\,
            I => \N__22986\
        );

    \I__3070\ : Span4Mux_h
    port map (
            O => \N__22994\,
            I => \N__22979\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__22991\,
            I => \N__22979\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__22986\,
            I => \N__22979\
        );

    \I__3067\ : Odrv4
    port map (
            O => \N__22979\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__3066\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22973\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__22973\,
            I => \N__22968\
        );

    \I__3064\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22965\
        );

    \I__3063\ : InMux
    port map (
            O => \N__22971\,
            I => \N__22962\
        );

    \I__3062\ : Span4Mux_h
    port map (
            O => \N__22968\,
            I => \N__22957\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__22965\,
            I => \N__22957\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__22962\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__22957\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__3058\ : InMux
    port map (
            O => \N__22952\,
            I => \N__22949\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__22949\,
            I => \N__22945\
        );

    \I__3056\ : InMux
    port map (
            O => \N__22948\,
            I => \N__22941\
        );

    \I__3055\ : Span4Mux_h
    port map (
            O => \N__22945\,
            I => \N__22938\
        );

    \I__3054\ : InMux
    port map (
            O => \N__22944\,
            I => \N__22935\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__22941\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__3052\ : Odrv4
    port map (
            O => \N__22938\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__22935\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__3050\ : InMux
    port map (
            O => \N__22928\,
            I => \N__22925\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__22925\,
            I => \N__22922\
        );

    \I__3048\ : Span4Mux_h
    port map (
            O => \N__22922\,
            I => \N__22918\
        );

    \I__3047\ : InMux
    port map (
            O => \N__22921\,
            I => \N__22915\
        );

    \I__3046\ : Sp12to4
    port map (
            O => \N__22918\,
            I => \N__22912\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__22915\,
            I => \N__22909\
        );

    \I__3044\ : Span12Mux_v
    port map (
            O => \N__22912\,
            I => \N__22904\
        );

    \I__3043\ : Span12Mux_v
    port map (
            O => \N__22909\,
            I => \N__22904\
        );

    \I__3042\ : Odrv12
    port map (
            O => \N__22904\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__3041\ : InMux
    port map (
            O => \N__22901\,
            I => \N__22897\
        );

    \I__3040\ : InMux
    port map (
            O => \N__22900\,
            I => \N__22894\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__22897\,
            I => \N__22891\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__22894\,
            I => \N__22888\
        );

    \I__3037\ : Span4Mux_h
    port map (
            O => \N__22891\,
            I => \N__22885\
        );

    \I__3036\ : Span4Mux_v
    port map (
            O => \N__22888\,
            I => \N__22882\
        );

    \I__3035\ : Sp12to4
    port map (
            O => \N__22885\,
            I => \N__22879\
        );

    \I__3034\ : Span4Mux_h
    port map (
            O => \N__22882\,
            I => \N__22876\
        );

    \I__3033\ : Odrv12
    port map (
            O => \N__22879\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__3032\ : Odrv4
    port map (
            O => \N__22876\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__3031\ : InMux
    port map (
            O => \N__22871\,
            I => \N__22868\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__22868\,
            I => \N__22864\
        );

    \I__3029\ : InMux
    port map (
            O => \N__22867\,
            I => \N__22861\
        );

    \I__3028\ : Span4Mux_h
    port map (
            O => \N__22864\,
            I => \N__22858\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__22861\,
            I => \N__22855\
        );

    \I__3026\ : Sp12to4
    port map (
            O => \N__22858\,
            I => \N__22850\
        );

    \I__3025\ : Span12Mux_s7_h
    port map (
            O => \N__22855\,
            I => \N__22850\
        );

    \I__3024\ : Odrv12
    port map (
            O => \N__22850\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__3023\ : InMux
    port map (
            O => \N__22847\,
            I => \N__22843\
        );

    \I__3022\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22840\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__22843\,
            I => \N__22837\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__22840\,
            I => \N__22834\
        );

    \I__3019\ : Sp12to4
    port map (
            O => \N__22837\,
            I => \N__22831\
        );

    \I__3018\ : Span4Mux_s3_h
    port map (
            O => \N__22834\,
            I => \N__22828\
        );

    \I__3017\ : Span12Mux_v
    port map (
            O => \N__22831\,
            I => \N__22825\
        );

    \I__3016\ : Span4Mux_h
    port map (
            O => \N__22828\,
            I => \N__22822\
        );

    \I__3015\ : Odrv12
    port map (
            O => \N__22825\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__3014\ : Odrv4
    port map (
            O => \N__22822\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__22817\,
            I => \N__22814\
        );

    \I__3012\ : InMux
    port map (
            O => \N__22814\,
            I => \N__22811\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__22811\,
            I => \N__22808\
        );

    \I__3010\ : Odrv12
    port map (
            O => \N__22808\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__3009\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22801\
        );

    \I__3008\ : InMux
    port map (
            O => \N__22804\,
            I => \N__22798\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__22801\,
            I => \N__22795\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__22798\,
            I => \N__22792\
        );

    \I__3005\ : Span4Mux_h
    port map (
            O => \N__22795\,
            I => \N__22789\
        );

    \I__3004\ : Span4Mux_s3_h
    port map (
            O => \N__22792\,
            I => \N__22786\
        );

    \I__3003\ : Sp12to4
    port map (
            O => \N__22789\,
            I => \N__22783\
        );

    \I__3002\ : Span4Mux_h
    port map (
            O => \N__22786\,
            I => \N__22780\
        );

    \I__3001\ : Odrv12
    port map (
            O => \N__22783\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__3000\ : Odrv4
    port map (
            O => \N__22780\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__22775\,
            I => \N__22772\
        );

    \I__2998\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22769\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__22769\,
            I => \N__22766\
        );

    \I__2996\ : Odrv4
    port map (
            O => \N__22766\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__22763\,
            I => \N__22760\
        );

    \I__2994\ : InMux
    port map (
            O => \N__22760\,
            I => \N__22757\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__22757\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__2992\ : InMux
    port map (
            O => \N__22754\,
            I => \N__22751\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__22751\,
            I => \N__22748\
        );

    \I__2990\ : Odrv4
    port map (
            O => \N__22748\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__2989\ : InMux
    port map (
            O => \N__22745\,
            I => \N__22742\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__22742\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__2987\ : InMux
    port map (
            O => \N__22739\,
            I => \N__22736\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__22736\,
            I => \N__22733\
        );

    \I__2985\ : Odrv12
    port map (
            O => \N__22733\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__2984\ : InMux
    port map (
            O => \N__22730\,
            I => \N__22727\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__22727\,
            I => \N__22724\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__22724\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__2981\ : CascadeMux
    port map (
            O => \N__22721\,
            I => \N__22718\
        );

    \I__2980\ : InMux
    port map (
            O => \N__22718\,
            I => \N__22715\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__22715\,
            I => \N__22712\
        );

    \I__2978\ : Odrv4
    port map (
            O => \N__22712\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__22709\,
            I => \N__22706\
        );

    \I__2976\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22703\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__22703\,
            I => \N__22700\
        );

    \I__2974\ : Odrv4
    port map (
            O => \N__22700\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__2973\ : InMux
    port map (
            O => \N__22697\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__2972\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22691\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__22691\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__22688\,
            I => \N__22685\
        );

    \I__2969\ : InMux
    port map (
            O => \N__22685\,
            I => \N__22682\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__22682\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__2967\ : InMux
    port map (
            O => \N__22679\,
            I => \N__22676\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__22676\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__2965\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22670\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__22670\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__2963\ : InMux
    port map (
            O => \N__22667\,
            I => \N__22664\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__22664\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__2961\ : CascadeMux
    port map (
            O => \N__22661\,
            I => \N__22658\
        );

    \I__2960\ : InMux
    port map (
            O => \N__22658\,
            I => \N__22655\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__22655\,
            I => \N__22652\
        );

    \I__2958\ : Odrv4
    port map (
            O => \N__22652\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__2957\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22646\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__22646\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__22643\,
            I => \N__22640\
        );

    \I__2954\ : InMux
    port map (
            O => \N__22640\,
            I => \N__22637\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__22637\,
            I => \N__22633\
        );

    \I__2952\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22630\
        );

    \I__2951\ : Span4Mux_h
    port map (
            O => \N__22633\,
            I => \N__22627\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__22630\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__22627\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__2948\ : InMux
    port map (
            O => \N__22622\,
            I => \N__22619\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__22619\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__2946\ : InMux
    port map (
            O => \N__22616\,
            I => \N__22613\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__22613\,
            I => \N__22610\
        );

    \I__2944\ : Span4Mux_h
    port map (
            O => \N__22610\,
            I => \N__22607\
        );

    \I__2943\ : Odrv4
    port map (
            O => \N__22607\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__2942\ : InMux
    port map (
            O => \N__22604\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__2941\ : InMux
    port map (
            O => \N__22601\,
            I => \N__22598\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__22598\,
            I => \N__22595\
        );

    \I__2939\ : Span4Mux_v
    port map (
            O => \N__22595\,
            I => \N__22592\
        );

    \I__2938\ : Odrv4
    port map (
            O => \N__22592\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__2937\ : InMux
    port map (
            O => \N__22589\,
            I => \bfn_9_15_0_\
        );

    \I__2936\ : InMux
    port map (
            O => \N__22586\,
            I => \N__22583\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__22583\,
            I => \N__22580\
        );

    \I__2934\ : Span4Mux_v
    port map (
            O => \N__22580\,
            I => \N__22577\
        );

    \I__2933\ : Odrv4
    port map (
            O => \N__22577\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__2932\ : InMux
    port map (
            O => \N__22574\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__2931\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22568\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__22568\,
            I => \N__22565\
        );

    \I__2929\ : Span4Mux_h
    port map (
            O => \N__22565\,
            I => \N__22562\
        );

    \I__2928\ : Odrv4
    port map (
            O => \N__22562\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__2927\ : InMux
    port map (
            O => \N__22559\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__2926\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22553\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__22553\,
            I => \N__22550\
        );

    \I__2924\ : Span4Mux_h
    port map (
            O => \N__22550\,
            I => \N__22547\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__22547\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__2922\ : InMux
    port map (
            O => \N__22544\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__2921\ : InMux
    port map (
            O => \N__22541\,
            I => \N__22538\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__22538\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__2919\ : InMux
    port map (
            O => \N__22535\,
            I => \N__22532\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__22532\,
            I => \N__22529\
        );

    \I__2917\ : Span4Mux_h
    port map (
            O => \N__22529\,
            I => \N__22526\
        );

    \I__2916\ : Odrv4
    port map (
            O => \N__22526\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__2915\ : InMux
    port map (
            O => \N__22523\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__2914\ : InMux
    port map (
            O => \N__22520\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__2913\ : InMux
    port map (
            O => \N__22517\,
            I => \N__22514\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__22514\,
            I => \N__22511\
        );

    \I__2911\ : Span4Mux_h
    port map (
            O => \N__22511\,
            I => \N__22507\
        );

    \I__2910\ : InMux
    port map (
            O => \N__22510\,
            I => \N__22504\
        );

    \I__2909\ : Odrv4
    port map (
            O => \N__22507\,
            I => \current_shift_inst.control_input_31\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__22504\,
            I => \current_shift_inst.control_input_31\
        );

    \I__2907\ : InMux
    port map (
            O => \N__22499\,
            I => \N__22496\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__22496\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__2905\ : InMux
    port map (
            O => \N__22493\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_28\
        );

    \I__2904\ : InMux
    port map (
            O => \N__22490\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30\
        );

    \I__2903\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22484\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__22484\,
            I => \N__22481\
        );

    \I__2901\ : Span4Mux_v
    port map (
            O => \N__22481\,
            I => \N__22478\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__22478\,
            I => \current_shift_inst.control_input_18\
        );

    \I__2899\ : InMux
    port map (
            O => \N__22475\,
            I => \N__22472\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__22472\,
            I => \N__22469\
        );

    \I__2897\ : Span4Mux_v
    port map (
            O => \N__22469\,
            I => \N__22466\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__22466\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__2895\ : InMux
    port map (
            O => \N__22463\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__2894\ : InMux
    port map (
            O => \N__22460\,
            I => \N__22457\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__22457\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__2892\ : InMux
    port map (
            O => \N__22454\,
            I => \N__22451\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__22451\,
            I => \N__22448\
        );

    \I__2890\ : Span4Mux_h
    port map (
            O => \N__22448\,
            I => \N__22445\
        );

    \I__2889\ : Odrv4
    port map (
            O => \N__22445\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__2888\ : InMux
    port map (
            O => \N__22442\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__2887\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22436\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__22436\,
            I => \N__22433\
        );

    \I__2885\ : Span4Mux_h
    port map (
            O => \N__22433\,
            I => \N__22430\
        );

    \I__2884\ : Odrv4
    port map (
            O => \N__22430\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__2883\ : InMux
    port map (
            O => \N__22427\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__2882\ : InMux
    port map (
            O => \N__22424\,
            I => \N__22421\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__22421\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__2880\ : InMux
    port map (
            O => \N__22418\,
            I => \N__22415\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__22415\,
            I => \N__22412\
        );

    \I__2878\ : Span4Mux_h
    port map (
            O => \N__22412\,
            I => \N__22409\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__22409\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__2876\ : InMux
    port map (
            O => \N__22406\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__2875\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22400\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__22400\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__2873\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22394\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__22394\,
            I => \N__22391\
        );

    \I__2871\ : Span4Mux_h
    port map (
            O => \N__22391\,
            I => \N__22388\
        );

    \I__2870\ : Odrv4
    port map (
            O => \N__22388\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__2869\ : InMux
    port map (
            O => \N__22385\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__2868\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22379\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__22379\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__2866\ : InMux
    port map (
            O => \N__22376\,
            I => \N__22373\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__22373\,
            I => \N__22370\
        );

    \I__2864\ : Span4Mux_h
    port map (
            O => \N__22370\,
            I => \N__22367\
        );

    \I__2863\ : Odrv4
    port map (
            O => \N__22367\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__2862\ : InMux
    port map (
            O => \N__22364\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__2861\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22358\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__2859\ : Span12Mux_v
    port map (
            O => \N__22355\,
            I => \N__22352\
        );

    \I__2858\ : Odrv12
    port map (
            O => \N__22352\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__2857\ : CascadeMux
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__2856\ : InMux
    port map (
            O => \N__22346\,
            I => \N__22343\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__22343\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__2854\ : InMux
    port map (
            O => \N__22340\,
            I => \N__22337\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__22337\,
            I => \N__22334\
        );

    \I__2852\ : Odrv12
    port map (
            O => \N__22334\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt18\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__22331\,
            I => \N__22328\
        );

    \I__2850\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__2848\ : Span4Mux_h
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__2847\ : Span4Mux_v
    port map (
            O => \N__22319\,
            I => \N__22316\
        );

    \I__2846\ : Odrv4
    port map (
            O => \N__22316\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\
        );

    \I__2845\ : InMux
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__2843\ : Odrv12
    port map (
            O => \N__22307\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\
        );

    \I__2842\ : CascadeMux
    port map (
            O => \N__22304\,
            I => \N__22301\
        );

    \I__2841\ : InMux
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__2839\ : Span4Mux_v
    port map (
            O => \N__22295\,
            I => \N__22292\
        );

    \I__2838\ : Odrv4
    port map (
            O => \N__22292\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt20\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22289\,
            I => \N__22286\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__22286\,
            I => \N__22283\
        );

    \I__2835\ : Span4Mux_h
    port map (
            O => \N__22283\,
            I => \N__22280\
        );

    \I__2834\ : Odrv4
    port map (
            O => \N__22280\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt22\
        );

    \I__2833\ : CascadeMux
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__2832\ : InMux
    port map (
            O => \N__22274\,
            I => \N__22271\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__22271\,
            I => \N__22268\
        );

    \I__2830\ : Span4Mux_h
    port map (
            O => \N__22268\,
            I => \N__22265\
        );

    \I__2829\ : Odrv4
    port map (
            O => \N__22265\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\
        );

    \I__2828\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22259\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__22259\,
            I => \N__22256\
        );

    \I__2826\ : Odrv12
    port map (
            O => \N__22256\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__2825\ : CascadeMux
    port map (
            O => \N__22253\,
            I => \N__22250\
        );

    \I__2824\ : InMux
    port map (
            O => \N__22250\,
            I => \N__22247\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__22247\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__2822\ : InMux
    port map (
            O => \N__22244\,
            I => \N__22241\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__22241\,
            I => \N__22238\
        );

    \I__2820\ : Odrv4
    port map (
            O => \N__22238\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__22235\,
            I => \N__22232\
        );

    \I__2818\ : InMux
    port map (
            O => \N__22232\,
            I => \N__22229\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__22229\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__22226\,
            I => \N__22223\
        );

    \I__2815\ : InMux
    port map (
            O => \N__22223\,
            I => \N__22220\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__22220\,
            I => \N__22217\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__22217\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__2812\ : InMux
    port map (
            O => \N__22214\,
            I => \N__22211\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__22211\,
            I => \N__22208\
        );

    \I__2810\ : Span4Mux_h
    port map (
            O => \N__22208\,
            I => \N__22205\
        );

    \I__2809\ : Odrv4
    port map (
            O => \N__22205\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__2808\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22199\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__22199\,
            I => \N__22196\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__22196\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__22193\,
            I => \N__22190\
        );

    \I__2804\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__22187\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__2802\ : InMux
    port map (
            O => \N__22184\,
            I => \N__22181\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__2800\ : Odrv12
    port map (
            O => \N__22178\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__2799\ : CascadeMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__2798\ : InMux
    port map (
            O => \N__22172\,
            I => \N__22169\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__2796\ : Odrv4
    port map (
            O => \N__22166\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__2795\ : InMux
    port map (
            O => \N__22163\,
            I => \N__22160\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__22160\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__22157\,
            I => \N__22154\
        );

    \I__2792\ : InMux
    port map (
            O => \N__22154\,
            I => \N__22151\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__22151\,
            I => \N__22148\
        );

    \I__2790\ : Odrv4
    port map (
            O => \N__22148\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__2789\ : InMux
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__2787\ : Span4Mux_v
    port map (
            O => \N__22139\,
            I => \N__22136\
        );

    \I__2786\ : Odrv4
    port map (
            O => \N__22136\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__22133\,
            I => \N__22130\
        );

    \I__2784\ : InMux
    port map (
            O => \N__22130\,
            I => \N__22127\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__22127\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__22124\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__22121\,
            I => \N__22118\
        );

    \I__2780\ : InMux
    port map (
            O => \N__22118\,
            I => \N__22115\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__22115\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__2778\ : InMux
    port map (
            O => \N__22112\,
            I => \N__22109\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__22109\,
            I => \N__22106\
        );

    \I__2776\ : Odrv4
    port map (
            O => \N__22106\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__2775\ : CascadeMux
    port map (
            O => \N__22103\,
            I => \N__22100\
        );

    \I__2774\ : InMux
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__22097\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__2772\ : CascadeMux
    port map (
            O => \N__22094\,
            I => \N__22091\
        );

    \I__2771\ : InMux
    port map (
            O => \N__22091\,
            I => \N__22088\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__22088\,
            I => \N__22085\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__22085\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__2768\ : InMux
    port map (
            O => \N__22082\,
            I => \N__22079\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__22079\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__2766\ : InMux
    port map (
            O => \N__22076\,
            I => \N__22073\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__22073\,
            I => \N__22070\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__22070\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__22067\,
            I => \N__22064\
        );

    \I__2762\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22061\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__22061\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__2760\ : InMux
    port map (
            O => \N__22058\,
            I => \N__22055\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__22055\,
            I => \N__22052\
        );

    \I__2758\ : Span4Mux_v
    port map (
            O => \N__22052\,
            I => \N__22049\
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__22049\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__22046\,
            I => \N__22043\
        );

    \I__2755\ : InMux
    port map (
            O => \N__22043\,
            I => \N__22040\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__22040\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__2753\ : InMux
    port map (
            O => \N__22037\,
            I => \N__22034\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__22034\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\
        );

    \I__2751\ : CascadeMux
    port map (
            O => \N__22031\,
            I => \N__22028\
        );

    \I__2750\ : InMux
    port map (
            O => \N__22028\,
            I => \N__22025\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__22025\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__2748\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22018\
        );

    \I__2747\ : InMux
    port map (
            O => \N__22021\,
            I => \N__22015\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__22018\,
            I => \N__22012\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__22015\,
            I => \N__22009\
        );

    \I__2744\ : Odrv4
    port map (
            O => \N__22012\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__2743\ : Odrv4
    port map (
            O => \N__22009\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__2742\ : InMux
    port map (
            O => \N__22004\,
            I => \N__22001\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__22001\,
            I => \N__21997\
        );

    \I__2740\ : InMux
    port map (
            O => \N__22000\,
            I => \N__21994\
        );

    \I__2739\ : Span4Mux_h
    port map (
            O => \N__21997\,
            I => \N__21991\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__21994\,
            I => \N__21988\
        );

    \I__2737\ : Odrv4
    port map (
            O => \N__21991\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__2736\ : Odrv4
    port map (
            O => \N__21988\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__2735\ : InMux
    port map (
            O => \N__21983\,
            I => \N__21977\
        );

    \I__2734\ : InMux
    port map (
            O => \N__21982\,
            I => \N__21977\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__21977\,
            I => \N__21974\
        );

    \I__2732\ : Span4Mux_v
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__2731\ : Odrv4
    port map (
            O => \N__21971\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\
        );

    \I__2730\ : InMux
    port map (
            O => \N__21968\,
            I => \N__21965\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__21965\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__21962\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21_cascade_\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__21959\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\
        );

    \I__2726\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21952\
        );

    \I__2725\ : InMux
    port map (
            O => \N__21955\,
            I => \N__21948\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__21952\,
            I => \N__21945\
        );

    \I__2723\ : InMux
    port map (
            O => \N__21951\,
            I => \N__21942\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__21948\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__2721\ : Odrv12
    port map (
            O => \N__21945\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__21942\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__21935\,
            I => \N__21932\
        );

    \I__2718\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__21929\,
            I => \N__21924\
        );

    \I__2716\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21921\
        );

    \I__2715\ : InMux
    port map (
            O => \N__21927\,
            I => \N__21918\
        );

    \I__2714\ : Span4Mux_v
    port map (
            O => \N__21924\,
            I => \N__21915\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__21921\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__21918\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__2711\ : Odrv4
    port map (
            O => \N__21915\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__2710\ : InMux
    port map (
            O => \N__21908\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__2709\ : InMux
    port map (
            O => \N__21905\,
            I => \N__21901\
        );

    \I__2708\ : InMux
    port map (
            O => \N__21904\,
            I => \N__21898\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__21901\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__21898\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__2705\ : IoInMux
    port map (
            O => \N__21893\,
            I => \N__21890\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__21890\,
            I => \N__21887\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__21887\,
            I => s4_phy_c
        );

    \I__2702\ : IoInMux
    port map (
            O => \N__21884\,
            I => \N__21881\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__21881\,
            I => \GB_BUFFER_clock_output_0_THRU_CO\
        );

    \I__2700\ : InMux
    port map (
            O => \N__21878\,
            I => \N__21875\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__21875\,
            I => \N__21872\
        );

    \I__2698\ : Odrv4
    port map (
            O => \N__21872\,
            I => il_min_comp1_c
        );

    \I__2697\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21864\
        );

    \I__2696\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21861\
        );

    \I__2695\ : InMux
    port map (
            O => \N__21867\,
            I => \N__21858\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__21864\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__21861\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__21858\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__2691\ : InMux
    port map (
            O => \N__21851\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__21848\,
            I => \N__21844\
        );

    \I__2689\ : InMux
    port map (
            O => \N__21847\,
            I => \N__21840\
        );

    \I__2688\ : InMux
    port map (
            O => \N__21844\,
            I => \N__21837\
        );

    \I__2687\ : InMux
    port map (
            O => \N__21843\,
            I => \N__21834\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__21840\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__21837\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__21834\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__2683\ : InMux
    port map (
            O => \N__21827\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__21824\,
            I => \N__21820\
        );

    \I__2681\ : InMux
    port map (
            O => \N__21823\,
            I => \N__21816\
        );

    \I__2680\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21813\
        );

    \I__2679\ : InMux
    port map (
            O => \N__21819\,
            I => \N__21810\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__21816\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__21813\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__21810\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__2675\ : InMux
    port map (
            O => \N__21803\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__21800\,
            I => \N__21796\
        );

    \I__2673\ : InMux
    port map (
            O => \N__21799\,
            I => \N__21792\
        );

    \I__2672\ : InMux
    port map (
            O => \N__21796\,
            I => \N__21789\
        );

    \I__2671\ : InMux
    port map (
            O => \N__21795\,
            I => \N__21786\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__21792\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__21789\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__21786\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__2667\ : InMux
    port map (
            O => \N__21779\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__21776\,
            I => \N__21772\
        );

    \I__2665\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21768\
        );

    \I__2664\ : InMux
    port map (
            O => \N__21772\,
            I => \N__21765\
        );

    \I__2663\ : InMux
    port map (
            O => \N__21771\,
            I => \N__21762\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__21768\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__21765\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__21762\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__2659\ : InMux
    port map (
            O => \N__21755\,
            I => \bfn_8_22_0_\
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__21752\,
            I => \N__21748\
        );

    \I__2657\ : InMux
    port map (
            O => \N__21751\,
            I => \N__21744\
        );

    \I__2656\ : InMux
    port map (
            O => \N__21748\,
            I => \N__21741\
        );

    \I__2655\ : InMux
    port map (
            O => \N__21747\,
            I => \N__21738\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__21744\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__21741\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__21738\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__2651\ : InMux
    port map (
            O => \N__21731\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__21728\,
            I => \N__21724\
        );

    \I__2649\ : InMux
    port map (
            O => \N__21727\,
            I => \N__21720\
        );

    \I__2648\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21717\
        );

    \I__2647\ : InMux
    port map (
            O => \N__21723\,
            I => \N__21714\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__21720\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__21717\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__21714\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__2643\ : InMux
    port map (
            O => \N__21707\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__21704\,
            I => \N__21700\
        );

    \I__2641\ : InMux
    port map (
            O => \N__21703\,
            I => \N__21696\
        );

    \I__2640\ : InMux
    port map (
            O => \N__21700\,
            I => \N__21693\
        );

    \I__2639\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21690\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__21696\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__21693\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__21690\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__2635\ : InMux
    port map (
            O => \N__21683\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__2634\ : InMux
    port map (
            O => \N__21680\,
            I => \N__21676\
        );

    \I__2633\ : InMux
    port map (
            O => \N__21679\,
            I => \N__21673\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__21676\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__21673\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__2630\ : InMux
    port map (
            O => \N__21668\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__21665\,
            I => \N__21661\
        );

    \I__2628\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21657\
        );

    \I__2627\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21654\
        );

    \I__2626\ : InMux
    port map (
            O => \N__21660\,
            I => \N__21651\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__21657\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__21654\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__21651\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__2622\ : InMux
    port map (
            O => \N__21644\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__21641\,
            I => \N__21637\
        );

    \I__2620\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21633\
        );

    \I__2619\ : InMux
    port map (
            O => \N__21637\,
            I => \N__21630\
        );

    \I__2618\ : InMux
    port map (
            O => \N__21636\,
            I => \N__21627\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__21633\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__21630\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__21627\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__2614\ : InMux
    port map (
            O => \N__21620\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__21617\,
            I => \N__21613\
        );

    \I__2612\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21609\
        );

    \I__2611\ : InMux
    port map (
            O => \N__21613\,
            I => \N__21606\
        );

    \I__2610\ : InMux
    port map (
            O => \N__21612\,
            I => \N__21603\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__21609\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__21606\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__21603\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__2606\ : InMux
    port map (
            O => \N__21596\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__21593\,
            I => \N__21589\
        );

    \I__2604\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21585\
        );

    \I__2603\ : InMux
    port map (
            O => \N__21589\,
            I => \N__21582\
        );

    \I__2602\ : InMux
    port map (
            O => \N__21588\,
            I => \N__21579\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__21585\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__21582\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__21579\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__2598\ : InMux
    port map (
            O => \N__21572\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__21569\,
            I => \N__21565\
        );

    \I__2596\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21561\
        );

    \I__2595\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21558\
        );

    \I__2594\ : InMux
    port map (
            O => \N__21564\,
            I => \N__21555\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__21561\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__21558\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__21555\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__2590\ : InMux
    port map (
            O => \N__21548\,
            I => \bfn_8_21_0_\
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__21545\,
            I => \N__21541\
        );

    \I__2588\ : InMux
    port map (
            O => \N__21544\,
            I => \N__21537\
        );

    \I__2587\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21534\
        );

    \I__2586\ : InMux
    port map (
            O => \N__21540\,
            I => \N__21531\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__21537\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__21534\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__21531\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__2582\ : InMux
    port map (
            O => \N__21524\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__2581\ : CascadeMux
    port map (
            O => \N__21521\,
            I => \N__21517\
        );

    \I__2580\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21513\
        );

    \I__2579\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21510\
        );

    \I__2578\ : InMux
    port map (
            O => \N__21516\,
            I => \N__21507\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__21513\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__21510\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__21507\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__2574\ : InMux
    port map (
            O => \N__21500\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__21497\,
            I => \N__21493\
        );

    \I__2572\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21489\
        );

    \I__2571\ : InMux
    port map (
            O => \N__21493\,
            I => \N__21486\
        );

    \I__2570\ : InMux
    port map (
            O => \N__21492\,
            I => \N__21483\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__21489\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__21486\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__21483\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__2566\ : InMux
    port map (
            O => \N__21476\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__21473\,
            I => \N__21469\
        );

    \I__2564\ : InMux
    port map (
            O => \N__21472\,
            I => \N__21465\
        );

    \I__2563\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21462\
        );

    \I__2562\ : InMux
    port map (
            O => \N__21468\,
            I => \N__21459\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__21465\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__21462\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__21459\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__21452\,
            I => \N__21448\
        );

    \I__2557\ : InMux
    port map (
            O => \N__21451\,
            I => \N__21444\
        );

    \I__2556\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21441\
        );

    \I__2555\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21438\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__21444\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__21441\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__21438\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__2551\ : InMux
    port map (
            O => \N__21431\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__21428\,
            I => \N__21424\
        );

    \I__2549\ : InMux
    port map (
            O => \N__21427\,
            I => \N__21420\
        );

    \I__2548\ : InMux
    port map (
            O => \N__21424\,
            I => \N__21417\
        );

    \I__2547\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21414\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__21420\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__21417\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__21414\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__2543\ : InMux
    port map (
            O => \N__21407\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__21404\,
            I => \N__21400\
        );

    \I__2541\ : InMux
    port map (
            O => \N__21403\,
            I => \N__21396\
        );

    \I__2540\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21393\
        );

    \I__2539\ : InMux
    port map (
            O => \N__21399\,
            I => \N__21390\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__21396\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__21393\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__21390\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__2535\ : InMux
    port map (
            O => \N__21383\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__21380\,
            I => \N__21376\
        );

    \I__2533\ : InMux
    port map (
            O => \N__21379\,
            I => \N__21372\
        );

    \I__2532\ : InMux
    port map (
            O => \N__21376\,
            I => \N__21369\
        );

    \I__2531\ : InMux
    port map (
            O => \N__21375\,
            I => \N__21366\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__21372\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__21369\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__21366\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__2527\ : InMux
    port map (
            O => \N__21359\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__21356\,
            I => \N__21352\
        );

    \I__2525\ : InMux
    port map (
            O => \N__21355\,
            I => \N__21348\
        );

    \I__2524\ : InMux
    port map (
            O => \N__21352\,
            I => \N__21345\
        );

    \I__2523\ : InMux
    port map (
            O => \N__21351\,
            I => \N__21342\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__21348\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__21345\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__21342\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__2519\ : InMux
    port map (
            O => \N__21335\,
            I => \bfn_8_20_0_\
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__21332\,
            I => \N__21328\
        );

    \I__2517\ : InMux
    port map (
            O => \N__21331\,
            I => \N__21324\
        );

    \I__2516\ : InMux
    port map (
            O => \N__21328\,
            I => \N__21321\
        );

    \I__2515\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21318\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__21324\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__21321\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__21318\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__2511\ : InMux
    port map (
            O => \N__21311\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__21308\,
            I => \N__21304\
        );

    \I__2509\ : InMux
    port map (
            O => \N__21307\,
            I => \N__21300\
        );

    \I__2508\ : InMux
    port map (
            O => \N__21304\,
            I => \N__21297\
        );

    \I__2507\ : InMux
    port map (
            O => \N__21303\,
            I => \N__21294\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__21300\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__21297\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__21294\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__2503\ : InMux
    port map (
            O => \N__21287\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__2502\ : CascadeMux
    port map (
            O => \N__21284\,
            I => \N__21280\
        );

    \I__2501\ : InMux
    port map (
            O => \N__21283\,
            I => \N__21276\
        );

    \I__2500\ : InMux
    port map (
            O => \N__21280\,
            I => \N__21273\
        );

    \I__2499\ : InMux
    port map (
            O => \N__21279\,
            I => \N__21270\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__21276\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__21273\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__21270\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__2495\ : InMux
    port map (
            O => \N__21263\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__2494\ : InMux
    port map (
            O => \N__21260\,
            I => \N__21257\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__21257\,
            I => \N__21252\
        );

    \I__2492\ : InMux
    port map (
            O => \N__21256\,
            I => \N__21249\
        );

    \I__2491\ : InMux
    port map (
            O => \N__21255\,
            I => \N__21246\
        );

    \I__2490\ : Odrv4
    port map (
            O => \N__21252\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__21249\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__21246\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__2487\ : InMux
    port map (
            O => \N__21239\,
            I => \bfn_8_19_0_\
        );

    \I__2486\ : InMux
    port map (
            O => \N__21236\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__21233\,
            I => \N__21228\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__21232\,
            I => \N__21225\
        );

    \I__2483\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21222\
        );

    \I__2482\ : InMux
    port map (
            O => \N__21228\,
            I => \N__21217\
        );

    \I__2481\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21217\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__21222\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__21217\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__2478\ : InMux
    port map (
            O => \N__21212\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__21209\,
            I => \N__21204\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__21208\,
            I => \N__21201\
        );

    \I__2475\ : InMux
    port map (
            O => \N__21207\,
            I => \N__21198\
        );

    \I__2474\ : InMux
    port map (
            O => \N__21204\,
            I => \N__21193\
        );

    \I__2473\ : InMux
    port map (
            O => \N__21201\,
            I => \N__21193\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__21198\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__21193\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__2470\ : InMux
    port map (
            O => \N__21188\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__2469\ : InMux
    port map (
            O => \N__21185\,
            I => \N__21182\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__21182\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__21179\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\
        );

    \I__2466\ : CascadeMux
    port map (
            O => \N__21176\,
            I => \N__21173\
        );

    \I__2465\ : InMux
    port map (
            O => \N__21173\,
            I => \N__21169\
        );

    \I__2464\ : InMux
    port map (
            O => \N__21172\,
            I => \N__21166\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__21169\,
            I => \N__21160\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__21166\,
            I => \N__21160\
        );

    \I__2461\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21157\
        );

    \I__2460\ : Span4Mux_v
    port map (
            O => \N__21160\,
            I => \N__21154\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__21157\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__2458\ : Odrv4
    port map (
            O => \N__21154\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__2457\ : InMux
    port map (
            O => \N__21149\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__2456\ : InMux
    port map (
            O => \N__21146\,
            I => \N__21142\
        );

    \I__2455\ : InMux
    port map (
            O => \N__21145\,
            I => \N__21139\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__21142\,
            I => \N__21136\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__21139\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__2452\ : Odrv12
    port map (
            O => \N__21136\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__21131\,
            I => \N__21128\
        );

    \I__2450\ : InMux
    port map (
            O => \N__21128\,
            I => \N__21123\
        );

    \I__2449\ : InMux
    port map (
            O => \N__21127\,
            I => \N__21120\
        );

    \I__2448\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21117\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__21123\,
            I => \N__21112\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__21120\,
            I => \N__21112\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__21117\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__2444\ : Odrv12
    port map (
            O => \N__21112\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__2443\ : InMux
    port map (
            O => \N__21107\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__2442\ : InMux
    port map (
            O => \N__21104\,
            I => \N__21100\
        );

    \I__2441\ : InMux
    port map (
            O => \N__21103\,
            I => \N__21097\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__21100\,
            I => \N__21094\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__21097\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__2438\ : Odrv12
    port map (
            O => \N__21094\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__2437\ : CascadeMux
    port map (
            O => \N__21089\,
            I => \N__21086\
        );

    \I__2436\ : InMux
    port map (
            O => \N__21086\,
            I => \N__21081\
        );

    \I__2435\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21078\
        );

    \I__2434\ : InMux
    port map (
            O => \N__21084\,
            I => \N__21075\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__21081\,
            I => \N__21070\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__21078\,
            I => \N__21070\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__21075\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__2430\ : Odrv12
    port map (
            O => \N__21070\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__2429\ : InMux
    port map (
            O => \N__21065\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__2428\ : InMux
    port map (
            O => \N__21062\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__2427\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21056\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__21056\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__21053\,
            I => \N__21050\
        );

    \I__2424\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21046\
        );

    \I__2423\ : InMux
    port map (
            O => \N__21049\,
            I => \N__21043\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__21046\,
            I => \N__21037\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__21043\,
            I => \N__21037\
        );

    \I__2420\ : InMux
    port map (
            O => \N__21042\,
            I => \N__21034\
        );

    \I__2419\ : Span4Mux_v
    port map (
            O => \N__21037\,
            I => \N__21031\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__21034\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__2417\ : Odrv4
    port map (
            O => \N__21031\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__2416\ : InMux
    port map (
            O => \N__21026\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__21023\,
            I => \N__21020\
        );

    \I__2414\ : InMux
    port map (
            O => \N__21020\,
            I => \N__21015\
        );

    \I__2413\ : InMux
    port map (
            O => \N__21019\,
            I => \N__21012\
        );

    \I__2412\ : InMux
    port map (
            O => \N__21018\,
            I => \N__21009\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__21015\,
            I => \N__21004\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__21012\,
            I => \N__21004\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__21009\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__2408\ : Odrv12
    port map (
            O => \N__21004\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__2407\ : InMux
    port map (
            O => \N__20999\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__2406\ : InMux
    port map (
            O => \N__20996\,
            I => \N__20989\
        );

    \I__2405\ : InMux
    port map (
            O => \N__20995\,
            I => \N__20989\
        );

    \I__2404\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20986\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__20989\,
            I => \N__20983\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__20986\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__2401\ : Odrv12
    port map (
            O => \N__20983\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__2400\ : InMux
    port map (
            O => \N__20978\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__2399\ : InMux
    port map (
            O => \N__20975\,
            I => \N__20968\
        );

    \I__2398\ : InMux
    port map (
            O => \N__20974\,
            I => \N__20968\
        );

    \I__2397\ : InMux
    port map (
            O => \N__20973\,
            I => \N__20965\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__20968\,
            I => \N__20962\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__20965\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__2394\ : Odrv12
    port map (
            O => \N__20962\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__2393\ : InMux
    port map (
            O => \N__20957\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__20954\,
            I => \N__20950\
        );

    \I__2391\ : InMux
    port map (
            O => \N__20953\,
            I => \N__20946\
        );

    \I__2390\ : InMux
    port map (
            O => \N__20950\,
            I => \N__20943\
        );

    \I__2389\ : InMux
    port map (
            O => \N__20949\,
            I => \N__20940\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__20946\,
            I => \N__20935\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__20943\,
            I => \N__20935\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__20940\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__2385\ : Odrv12
    port map (
            O => \N__20935\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__2384\ : InMux
    port map (
            O => \N__20930\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__2383\ : CascadeMux
    port map (
            O => \N__20927\,
            I => \N__20923\
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__20926\,
            I => \N__20920\
        );

    \I__2381\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20915\
        );

    \I__2380\ : InMux
    port map (
            O => \N__20920\,
            I => \N__20915\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__20915\,
            I => \N__20911\
        );

    \I__2378\ : InMux
    port map (
            O => \N__20914\,
            I => \N__20908\
        );

    \I__2377\ : Span4Mux_v
    port map (
            O => \N__20911\,
            I => \N__20905\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__20908\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__20905\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__2374\ : InMux
    port map (
            O => \N__20900\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__20897\,
            I => \N__20893\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__20896\,
            I => \N__20890\
        );

    \I__2371\ : InMux
    port map (
            O => \N__20893\,
            I => \N__20884\
        );

    \I__2370\ : InMux
    port map (
            O => \N__20890\,
            I => \N__20884\
        );

    \I__2369\ : InMux
    port map (
            O => \N__20889\,
            I => \N__20881\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__20884\,
            I => \N__20878\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__20881\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__2366\ : Odrv12
    port map (
            O => \N__20878\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__2365\ : InMux
    port map (
            O => \N__20873\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__20870\,
            I => \N__20867\
        );

    \I__2363\ : InMux
    port map (
            O => \N__20867\,
            I => \N__20863\
        );

    \I__2362\ : InMux
    port map (
            O => \N__20866\,
            I => \N__20860\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__20863\,
            I => \N__20854\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__20860\,
            I => \N__20854\
        );

    \I__2359\ : InMux
    port map (
            O => \N__20859\,
            I => \N__20851\
        );

    \I__2358\ : Span4Mux_v
    port map (
            O => \N__20854\,
            I => \N__20848\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__20851\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__20848\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__2355\ : InMux
    port map (
            O => \N__20843\,
            I => \bfn_8_14_0_\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__20840\,
            I => \N__20837\
        );

    \I__2353\ : InMux
    port map (
            O => \N__20837\,
            I => \N__20833\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__20836\,
            I => \N__20830\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__20833\,
            I => \N__20826\
        );

    \I__2350\ : InMux
    port map (
            O => \N__20830\,
            I => \N__20823\
        );

    \I__2349\ : InMux
    port map (
            O => \N__20829\,
            I => \N__20820\
        );

    \I__2348\ : Sp12to4
    port map (
            O => \N__20826\,
            I => \N__20815\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__20823\,
            I => \N__20815\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__20820\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__2345\ : Odrv12
    port map (
            O => \N__20815\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__2344\ : InMux
    port map (
            O => \N__20810\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__2343\ : InMux
    port map (
            O => \N__20807\,
            I => \N__20801\
        );

    \I__2342\ : InMux
    port map (
            O => \N__20806\,
            I => \N__20801\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__20801\,
            I => \N__20797\
        );

    \I__2340\ : InMux
    port map (
            O => \N__20800\,
            I => \N__20794\
        );

    \I__2339\ : Span4Mux_v
    port map (
            O => \N__20797\,
            I => \N__20791\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__20794\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__2337\ : Odrv4
    port map (
            O => \N__20791\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__2336\ : InMux
    port map (
            O => \N__20786\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__2335\ : InMux
    port map (
            O => \N__20783\,
            I => \N__20776\
        );

    \I__2334\ : InMux
    port map (
            O => \N__20782\,
            I => \N__20776\
        );

    \I__2333\ : InMux
    port map (
            O => \N__20781\,
            I => \N__20773\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__20776\,
            I => \N__20770\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__20773\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__2330\ : Odrv12
    port map (
            O => \N__20770\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__2329\ : InMux
    port map (
            O => \N__20765\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__2328\ : CascadeMux
    port map (
            O => \N__20762\,
            I => \N__20758\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__20761\,
            I => \N__20755\
        );

    \I__2326\ : InMux
    port map (
            O => \N__20758\,
            I => \N__20749\
        );

    \I__2325\ : InMux
    port map (
            O => \N__20755\,
            I => \N__20749\
        );

    \I__2324\ : InMux
    port map (
            O => \N__20754\,
            I => \N__20746\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__20749\,
            I => \N__20743\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__20746\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__2321\ : Odrv12
    port map (
            O => \N__20743\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__2320\ : InMux
    port map (
            O => \N__20738\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__20735\,
            I => \N__20731\
        );

    \I__2318\ : CascadeMux
    port map (
            O => \N__20734\,
            I => \N__20728\
        );

    \I__2317\ : InMux
    port map (
            O => \N__20731\,
            I => \N__20722\
        );

    \I__2316\ : InMux
    port map (
            O => \N__20728\,
            I => \N__20722\
        );

    \I__2315\ : InMux
    port map (
            O => \N__20727\,
            I => \N__20719\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__20722\,
            I => \N__20716\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__20719\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__2312\ : Odrv12
    port map (
            O => \N__20716\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__2311\ : InMux
    port map (
            O => \N__20711\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__20708\,
            I => \N__20705\
        );

    \I__2309\ : InMux
    port map (
            O => \N__20705\,
            I => \N__20701\
        );

    \I__2308\ : InMux
    port map (
            O => \N__20704\,
            I => \N__20698\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__20701\,
            I => \N__20692\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__20698\,
            I => \N__20692\
        );

    \I__2305\ : InMux
    port map (
            O => \N__20697\,
            I => \N__20689\
        );

    \I__2304\ : Span4Mux_v
    port map (
            O => \N__20692\,
            I => \N__20686\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__20689\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__20686\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__2301\ : InMux
    port map (
            O => \N__20681\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__20678\,
            I => \N__20675\
        );

    \I__2299\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20671\
        );

    \I__2298\ : InMux
    port map (
            O => \N__20674\,
            I => \N__20668\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__20671\,
            I => \N__20662\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__20668\,
            I => \N__20662\
        );

    \I__2295\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20659\
        );

    \I__2294\ : Span4Mux_v
    port map (
            O => \N__20662\,
            I => \N__20656\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__20659\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__2292\ : Odrv4
    port map (
            O => \N__20656\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__2291\ : InMux
    port map (
            O => \N__20651\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__2290\ : CascadeMux
    port map (
            O => \N__20648\,
            I => \N__20645\
        );

    \I__2289\ : InMux
    port map (
            O => \N__20645\,
            I => \N__20640\
        );

    \I__2288\ : InMux
    port map (
            O => \N__20644\,
            I => \N__20637\
        );

    \I__2287\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20634\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__20640\,
            I => \N__20629\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__20637\,
            I => \N__20629\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__20634\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__2283\ : Odrv12
    port map (
            O => \N__20629\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__2282\ : InMux
    port map (
            O => \N__20624\,
            I => \bfn_8_13_0_\
        );

    \I__2281\ : InMux
    port map (
            O => \N__20621\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__20618\,
            I => \N__20614\
        );

    \I__2279\ : InMux
    port map (
            O => \N__20617\,
            I => \N__20611\
        );

    \I__2278\ : InMux
    port map (
            O => \N__20614\,
            I => \N__20608\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__20611\,
            I => \N__20602\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__20608\,
            I => \N__20602\
        );

    \I__2275\ : InMux
    port map (
            O => \N__20607\,
            I => \N__20599\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__20602\,
            I => \N__20596\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__20599\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__20596\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__2271\ : InMux
    port map (
            O => \N__20591\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__2270\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20582\
        );

    \I__2269\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20582\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__20582\,
            I => \N__20578\
        );

    \I__2267\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20575\
        );

    \I__2266\ : Span4Mux_v
    port map (
            O => \N__20578\,
            I => \N__20572\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__20575\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__20572\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__2263\ : InMux
    port map (
            O => \N__20567\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__20564\,
            I => \N__20560\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__20563\,
            I => \N__20557\
        );

    \I__2260\ : InMux
    port map (
            O => \N__20560\,
            I => \N__20551\
        );

    \I__2259\ : InMux
    port map (
            O => \N__20557\,
            I => \N__20551\
        );

    \I__2258\ : InMux
    port map (
            O => \N__20556\,
            I => \N__20548\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__20551\,
            I => \N__20545\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__20548\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__2255\ : Odrv12
    port map (
            O => \N__20545\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__2254\ : InMux
    port map (
            O => \N__20540\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__20537\,
            I => \N__20533\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__20536\,
            I => \N__20530\
        );

    \I__2251\ : InMux
    port map (
            O => \N__20533\,
            I => \N__20524\
        );

    \I__2250\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20524\
        );

    \I__2249\ : InMux
    port map (
            O => \N__20529\,
            I => \N__20521\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__20524\,
            I => \N__20518\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__20521\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__2246\ : Odrv12
    port map (
            O => \N__20518\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__2245\ : InMux
    port map (
            O => \N__20513\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__2244\ : InMux
    port map (
            O => \N__20510\,
            I => \N__20504\
        );

    \I__2243\ : InMux
    port map (
            O => \N__20509\,
            I => \N__20504\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__20504\,
            I => \N__20500\
        );

    \I__2241\ : InMux
    port map (
            O => \N__20503\,
            I => \N__20497\
        );

    \I__2240\ : Span4Mux_v
    port map (
            O => \N__20500\,
            I => \N__20494\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__20497\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__20494\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__2237\ : InMux
    port map (
            O => \N__20489\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__2236\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20480\
        );

    \I__2235\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20480\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__20480\,
            I => \N__20476\
        );

    \I__2233\ : InMux
    port map (
            O => \N__20479\,
            I => \N__20473\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__20476\,
            I => \N__20470\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__20473\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__20470\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__2229\ : InMux
    port map (
            O => \N__20465\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__20462\,
            I => \N__20458\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__20461\,
            I => \N__20455\
        );

    \I__2226\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20452\
        );

    \I__2225\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20449\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__20452\,
            I => \N__20443\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__20449\,
            I => \N__20443\
        );

    \I__2222\ : InMux
    port map (
            O => \N__20448\,
            I => \N__20440\
        );

    \I__2221\ : Span4Mux_v
    port map (
            O => \N__20443\,
            I => \N__20437\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__20440\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__20437\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__2218\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20427\
        );

    \I__2217\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20424\
        );

    \I__2216\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20421\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__20427\,
            I => \N__20418\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__20424\,
            I => \N__20415\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__20421\,
            I => \N__20411\
        );

    \I__2212\ : Span4Mux_v
    port map (
            O => \N__20418\,
            I => \N__20406\
        );

    \I__2211\ : Span4Mux_h
    port map (
            O => \N__20415\,
            I => \N__20406\
        );

    \I__2210\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20403\
        );

    \I__2209\ : Odrv12
    port map (
            O => \N__20411\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__2208\ : Odrv4
    port map (
            O => \N__20406\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__20403\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__2206\ : InMux
    port map (
            O => \N__20396\,
            I => \bfn_8_12_0_\
        );

    \I__2205\ : InMux
    port map (
            O => \N__20393\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__2204\ : InMux
    port map (
            O => \N__20390\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__2203\ : InMux
    port map (
            O => \N__20387\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__2202\ : InMux
    port map (
            O => \N__20384\,
            I => \bfn_8_10_0_\
        );

    \I__2201\ : InMux
    port map (
            O => \N__20381\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__2200\ : InMux
    port map (
            O => \N__20378\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__2199\ : InMux
    port map (
            O => \N__20375\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__2198\ : InMux
    port map (
            O => \N__20372\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__2197\ : InMux
    port map (
            O => \N__20369\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__2196\ : InMux
    port map (
            O => \N__20366\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__2195\ : InMux
    port map (
            O => \N__20363\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__2194\ : InMux
    port map (
            O => \N__20360\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__2193\ : InMux
    port map (
            O => \N__20357\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__2192\ : InMux
    port map (
            O => \N__20354\,
            I => \bfn_8_9_0_\
        );

    \I__2191\ : InMux
    port map (
            O => \N__20351\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__2190\ : InMux
    port map (
            O => \N__20348\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__2189\ : InMux
    port map (
            O => \N__20345\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__2188\ : InMux
    port map (
            O => \N__20342\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__2187\ : InMux
    port map (
            O => \N__20339\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__2186\ : InMux
    port map (
            O => \N__20336\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__2185\ : InMux
    port map (
            O => \N__20333\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__2184\ : InMux
    port map (
            O => \N__20330\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__2183\ : InMux
    port map (
            O => \N__20327\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__2182\ : InMux
    port map (
            O => \N__20324\,
            I => \bfn_8_8_0_\
        );

    \I__2181\ : InMux
    port map (
            O => \N__20321\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__2180\ : InMux
    port map (
            O => \N__20318\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__2179\ : InMux
    port map (
            O => \N__20315\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__2178\ : InMux
    port map (
            O => \N__20312\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__2177\ : InMux
    port map (
            O => \N__20309\,
            I => \N__20305\
        );

    \I__2176\ : InMux
    port map (
            O => \N__20308\,
            I => \N__20302\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__20305\,
            I => \N__20299\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__20302\,
            I => \N__20296\
        );

    \I__2173\ : Span4Mux_v
    port map (
            O => \N__20299\,
            I => \N__20293\
        );

    \I__2172\ : Span12Mux_v
    port map (
            O => \N__20296\,
            I => \N__20290\
        );

    \I__2171\ : Span4Mux_h
    port map (
            O => \N__20293\,
            I => \N__20287\
        );

    \I__2170\ : Odrv12
    port map (
            O => \N__20290\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__20287\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__2168\ : InMux
    port map (
            O => \N__20282\,
            I => \N__20279\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__20279\,
            I => \N__20276\
        );

    \I__2166\ : Odrv12
    port map (
            O => \N__20276\,
            I => il_max_comp1_c
        );

    \I__2165\ : InMux
    port map (
            O => \N__20273\,
            I => \bfn_8_7_0_\
        );

    \I__2164\ : InMux
    port map (
            O => \N__20270\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__2163\ : InMux
    port map (
            O => \N__20267\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__2162\ : InMux
    port map (
            O => \N__20264\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__2161\ : InMux
    port map (
            O => \N__20261\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__2160\ : InMux
    port map (
            O => \N__20258\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__2159\ : InMux
    port map (
            O => \N__20255\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__2158\ : InMux
    port map (
            O => \N__20252\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__2157\ : InMux
    port map (
            O => \N__20249\,
            I => \bfn_7_23_0_\
        );

    \I__2156\ : InMux
    port map (
            O => \N__20246\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__2155\ : InMux
    port map (
            O => \N__20243\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__2154\ : InMux
    port map (
            O => \N__20240\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__2153\ : InMux
    port map (
            O => \N__20237\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__2152\ : InMux
    port map (
            O => \N__20234\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__2151\ : InMux
    port map (
            O => \N__20231\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__2150\ : InMux
    port map (
            O => \N__20228\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__2149\ : InMux
    port map (
            O => \N__20225\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__2148\ : InMux
    port map (
            O => \N__20222\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__2147\ : InMux
    port map (
            O => \N__20219\,
            I => \bfn_7_22_0_\
        );

    \I__2146\ : InMux
    port map (
            O => \N__20216\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__2145\ : InMux
    port map (
            O => \N__20213\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__2144\ : InMux
    port map (
            O => \N__20210\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__2143\ : InMux
    port map (
            O => \N__20207\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__2142\ : InMux
    port map (
            O => \N__20204\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20201\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__2140\ : InMux
    port map (
            O => \N__20198\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__2139\ : InMux
    port map (
            O => \N__20195\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__2138\ : InMux
    port map (
            O => \N__20192\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__2137\ : InMux
    port map (
            O => \N__20189\,
            I => \bfn_7_21_0_\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20186\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__2135\ : InMux
    port map (
            O => \N__20183\,
            I => \bfn_7_14_0_\
        );

    \I__2134\ : InMux
    port map (
            O => \N__20180\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__2133\ : InMux
    port map (
            O => \N__20177\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__2132\ : InMux
    port map (
            O => \N__20174\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__2131\ : InMux
    port map (
            O => \N__20171\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__2130\ : InMux
    port map (
            O => \N__20168\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__2129\ : InMux
    port map (
            O => \N__20165\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__2128\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20159\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__20159\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__2126\ : InMux
    port map (
            O => \N__20156\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__2125\ : InMux
    port map (
            O => \N__20153\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__2124\ : InMux
    port map (
            O => \N__20150\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__2123\ : InMux
    port map (
            O => \N__20147\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__2122\ : InMux
    port map (
            O => \N__20144\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__2121\ : InMux
    port map (
            O => \N__20141\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__2120\ : InMux
    port map (
            O => \N__20138\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__2119\ : CascadeMux
    port map (
            O => \N__20135\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_\
        );

    \I__2118\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20129\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__20129\,
            I => \N__20126\
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__20126\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__20123\,
            I => \N__20119\
        );

    \I__2114\ : InMux
    port map (
            O => \N__20122\,
            I => \N__20114\
        );

    \I__2113\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20114\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__20114\,
            I => \N__20111\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__20111\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\
        );

    \I__2110\ : InMux
    port map (
            O => \N__20108\,
            I => \N__20102\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20107\,
            I => \N__20102\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__20102\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\
        );

    \I__2107\ : InMux
    port map (
            O => \N__20099\,
            I => \N__20096\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__20096\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\
        );

    \I__2105\ : InMux
    port map (
            O => \N__20093\,
            I => \N__20090\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__20090\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__2103\ : InMux
    port map (
            O => \N__20087\,
            I => \N__20084\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__20084\,
            I => \N__20081\
        );

    \I__2101\ : Glb2LocalMux
    port map (
            O => \N__20081\,
            I => \N__20078\
        );

    \I__2100\ : GlobalMux
    port map (
            O => \N__20078\,
            I => clk_12mhz
        );

    \I__2099\ : IoInMux
    port map (
            O => \N__20075\,
            I => \N__20072\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__20072\,
            I => \N__20069\
        );

    \I__2097\ : IoSpan4Mux
    port map (
            O => \N__20069\,
            I => \N__20066\
        );

    \I__2096\ : Span4Mux_s0_v
    port map (
            O => \N__20066\,
            I => \N__20063\
        );

    \I__2095\ : Odrv4
    port map (
            O => \N__20063\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__2094\ : InMux
    port map (
            O => \N__20060\,
            I => \N__20057\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__20057\,
            I => \N__20052\
        );

    \I__2092\ : InMux
    port map (
            O => \N__20056\,
            I => \N__20049\
        );

    \I__2091\ : InMux
    port map (
            O => \N__20055\,
            I => \N__20046\
        );

    \I__2090\ : Span4Mux_h
    port map (
            O => \N__20052\,
            I => \N__20043\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__20049\,
            I => \N__20040\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__20046\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__20043\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__20040\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__20033\,
            I => \N__20030\
        );

    \I__2084\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20027\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__20027\,
            I => \N__20024\
        );

    \I__2082\ : Odrv4
    port map (
            O => \N__20024\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__2081\ : CascadeMux
    port map (
            O => \N__20021\,
            I => \N__20018\
        );

    \I__2080\ : InMux
    port map (
            O => \N__20018\,
            I => \N__20015\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__20015\,
            I => \N__20012\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__20012\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__2077\ : InMux
    port map (
            O => \N__20009\,
            I => \N__20005\
        );

    \I__2076\ : InMux
    port map (
            O => \N__20008\,
            I => \N__20002\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__20005\,
            I => \N__19992\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__20002\,
            I => \N__19992\
        );

    \I__2073\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19987\
        );

    \I__2072\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19987\
        );

    \I__2071\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19984\
        );

    \I__2070\ : InMux
    port map (
            O => \N__19998\,
            I => \N__19973\
        );

    \I__2069\ : InMux
    port map (
            O => \N__19997\,
            I => \N__19970\
        );

    \I__2068\ : Span4Mux_v
    port map (
            O => \N__19992\,
            I => \N__19953\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__19987\,
            I => \N__19953\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__19984\,
            I => \N__19950\
        );

    \I__2065\ : InMux
    port map (
            O => \N__19983\,
            I => \N__19947\
        );

    \I__2064\ : InMux
    port map (
            O => \N__19982\,
            I => \N__19940\
        );

    \I__2063\ : InMux
    port map (
            O => \N__19981\,
            I => \N__19940\
        );

    \I__2062\ : InMux
    port map (
            O => \N__19980\,
            I => \N__19940\
        );

    \I__2061\ : InMux
    port map (
            O => \N__19979\,
            I => \N__19931\
        );

    \I__2060\ : InMux
    port map (
            O => \N__19978\,
            I => \N__19931\
        );

    \I__2059\ : InMux
    port map (
            O => \N__19977\,
            I => \N__19931\
        );

    \I__2058\ : InMux
    port map (
            O => \N__19976\,
            I => \N__19931\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__19973\,
            I => \N__19928\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__19970\,
            I => \N__19922\
        );

    \I__2055\ : InMux
    port map (
            O => \N__19969\,
            I => \N__19907\
        );

    \I__2054\ : InMux
    port map (
            O => \N__19968\,
            I => \N__19907\
        );

    \I__2053\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19907\
        );

    \I__2052\ : InMux
    port map (
            O => \N__19966\,
            I => \N__19907\
        );

    \I__2051\ : InMux
    port map (
            O => \N__19965\,
            I => \N__19907\
        );

    \I__2050\ : InMux
    port map (
            O => \N__19964\,
            I => \N__19907\
        );

    \I__2049\ : InMux
    port map (
            O => \N__19963\,
            I => \N__19907\
        );

    \I__2048\ : InMux
    port map (
            O => \N__19962\,
            I => \N__19896\
        );

    \I__2047\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19896\
        );

    \I__2046\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19896\
        );

    \I__2045\ : InMux
    port map (
            O => \N__19959\,
            I => \N__19896\
        );

    \I__2044\ : InMux
    port map (
            O => \N__19958\,
            I => \N__19896\
        );

    \I__2043\ : Span4Mux_v
    port map (
            O => \N__19953\,
            I => \N__19892\
        );

    \I__2042\ : Span4Mux_v
    port map (
            O => \N__19950\,
            I => \N__19887\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__19947\,
            I => \N__19887\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__19940\,
            I => \N__19882\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__19931\,
            I => \N__19882\
        );

    \I__2038\ : Span4Mux_h
    port map (
            O => \N__19928\,
            I => \N__19879\
        );

    \I__2037\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19872\
        );

    \I__2036\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19872\
        );

    \I__2035\ : InMux
    port map (
            O => \N__19925\,
            I => \N__19872\
        );

    \I__2034\ : Span4Mux_h
    port map (
            O => \N__19922\,
            I => \N__19865\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__19907\,
            I => \N__19865\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__19896\,
            I => \N__19865\
        );

    \I__2031\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19862\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__19892\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__19887\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2028\ : Odrv12
    port map (
            O => \N__19882\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2027\ : Odrv4
    port map (
            O => \N__19879\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__19872\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2025\ : Odrv4
    port map (
            O => \N__19865\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__19862\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2023\ : CascadeMux
    port map (
            O => \N__19847\,
            I => \N__19844\
        );

    \I__2022\ : InMux
    port map (
            O => \N__19844\,
            I => \N__19841\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__19841\,
            I => \N__19838\
        );

    \I__2020\ : Span4Mux_h
    port map (
            O => \N__19838\,
            I => \N__19835\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__19835\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__19832\,
            I => \N__19825\
        );

    \I__2017\ : InMux
    port map (
            O => \N__19831\,
            I => \N__19811\
        );

    \I__2016\ : InMux
    port map (
            O => \N__19830\,
            I => \N__19808\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__19829\,
            I => \N__19799\
        );

    \I__2014\ : InMux
    port map (
            O => \N__19828\,
            I => \N__19796\
        );

    \I__2013\ : InMux
    port map (
            O => \N__19825\,
            I => \N__19789\
        );

    \I__2012\ : InMux
    port map (
            O => \N__19824\,
            I => \N__19789\
        );

    \I__2011\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19789\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__19822\,
            I => \N__19785\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__19821\,
            I => \N__19782\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__19820\,
            I => \N__19779\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__19819\,
            I => \N__19773\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__19818\,
            I => \N__19770\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__19817\,
            I => \N__19767\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__19816\,
            I => \N__19764\
        );

    \I__2003\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19761\
        );

    \I__2002\ : InMux
    port map (
            O => \N__19814\,
            I => \N__19758\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__19811\,
            I => \N__19755\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__19808\,
            I => \N__19752\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__19807\,
            I => \N__19749\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__19806\,
            I => \N__19744\
        );

    \I__1997\ : InMux
    port map (
            O => \N__19805\,
            I => \N__19741\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__19804\,
            I => \N__19735\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__19803\,
            I => \N__19732\
        );

    \I__1994\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19729\
        );

    \I__1993\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19726\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__19796\,
            I => \N__19721\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__19789\,
            I => \N__19721\
        );

    \I__1990\ : InMux
    port map (
            O => \N__19788\,
            I => \N__19712\
        );

    \I__1989\ : InMux
    port map (
            O => \N__19785\,
            I => \N__19712\
        );

    \I__1988\ : InMux
    port map (
            O => \N__19782\,
            I => \N__19712\
        );

    \I__1987\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19712\
        );

    \I__1986\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19697\
        );

    \I__1985\ : InMux
    port map (
            O => \N__19777\,
            I => \N__19697\
        );

    \I__1984\ : InMux
    port map (
            O => \N__19776\,
            I => \N__19697\
        );

    \I__1983\ : InMux
    port map (
            O => \N__19773\,
            I => \N__19697\
        );

    \I__1982\ : InMux
    port map (
            O => \N__19770\,
            I => \N__19697\
        );

    \I__1981\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19697\
        );

    \I__1980\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19697\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__19761\,
            I => \N__19694\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__19758\,
            I => \N__19687\
        );

    \I__1977\ : Span4Mux_h
    port map (
            O => \N__19755\,
            I => \N__19687\
        );

    \I__1976\ : Span4Mux_s3_h
    port map (
            O => \N__19752\,
            I => \N__19687\
        );

    \I__1975\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19684\
        );

    \I__1974\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19677\
        );

    \I__1973\ : InMux
    port map (
            O => \N__19747\,
            I => \N__19677\
        );

    \I__1972\ : InMux
    port map (
            O => \N__19744\,
            I => \N__19677\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__19741\,
            I => \N__19674\
        );

    \I__1970\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19663\
        );

    \I__1969\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19663\
        );

    \I__1968\ : InMux
    port map (
            O => \N__19738\,
            I => \N__19663\
        );

    \I__1967\ : InMux
    port map (
            O => \N__19735\,
            I => \N__19663\
        );

    \I__1966\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19663\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__19729\,
            I => \N__19658\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__19726\,
            I => \N__19658\
        );

    \I__1963\ : Span4Mux_h
    port map (
            O => \N__19721\,
            I => \N__19649\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__19712\,
            I => \N__19649\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__19697\,
            I => \N__19649\
        );

    \I__1960\ : Span4Mux_h
    port map (
            O => \N__19694\,
            I => \N__19649\
        );

    \I__1959\ : Span4Mux_v
    port map (
            O => \N__19687\,
            I => \N__19646\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__19684\,
            I => \N__19635\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__19677\,
            I => \N__19635\
        );

    \I__1956\ : Span4Mux_h
    port map (
            O => \N__19674\,
            I => \N__19635\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__19663\,
            I => \N__19635\
        );

    \I__1954\ : Span4Mux_h
    port map (
            O => \N__19658\,
            I => \N__19635\
        );

    \I__1953\ : Span4Mux_v
    port map (
            O => \N__19649\,
            I => \N__19632\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__19646\,
            I => \N__19629\
        );

    \I__1951\ : Span4Mux_v
    port map (
            O => \N__19635\,
            I => \N__19626\
        );

    \I__1950\ : Span4Mux_v
    port map (
            O => \N__19632\,
            I => \N__19623\
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__19629\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__19626\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__1947\ : Odrv4
    port map (
            O => \N__19623\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__19616\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\
        );

    \I__1945\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__19610\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__19607\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\
        );

    \I__1942\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19601\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__19601\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\
        );

    \I__1940\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__19595\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__19592\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\
        );

    \I__1937\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19586\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__19586\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\
        );

    \I__1935\ : CascadeMux
    port map (
            O => \N__19583\,
            I => \current_shift_inst.PI_CTRL.N_77_cascade_\
        );

    \I__1934\ : InMux
    port map (
            O => \N__19580\,
            I => \N__19577\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__19577\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__1932\ : InMux
    port map (
            O => \N__19574\,
            I => \N__19571\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__19571\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__19568\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\
        );

    \I__1929\ : InMux
    port map (
            O => \N__19565\,
            I => \N__19562\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__19562\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__19559\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_\
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__19556\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__19553\,
            I => \current_shift_inst.PI_CTRL.N_44_cascade_\
        );

    \I__1924\ : InMux
    port map (
            O => \N__19550\,
            I => \N__19547\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__19547\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\
        );

    \I__1922\ : InMux
    port map (
            O => \N__19544\,
            I => \N__19541\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__19541\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__19538\,
            I => \N__19535\
        );

    \I__1919\ : InMux
    port map (
            O => \N__19535\,
            I => \N__19532\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__19532\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__1917\ : InMux
    port map (
            O => \N__19529\,
            I => \N__19526\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__19526\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__19523\,
            I => \N__19520\
        );

    \I__1914\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19517\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__19517\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__1912\ : CascadeMux
    port map (
            O => \N__19514\,
            I => \N__19511\
        );

    \I__1911\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__19508\,
            I => \N__19505\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__19505\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__19502\,
            I => \N__19499\
        );

    \I__1907\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__19496\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__1905\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__19490\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__1903\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19484\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__19484\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__19481\,
            I => \N__19478\
        );

    \I__1900\ : InMux
    port map (
            O => \N__19478\,
            I => \N__19475\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__19475\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__1898\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19469\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__19469\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__1896\ : InMux
    port map (
            O => \N__19466\,
            I => \N__19463\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__19463\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__1894\ : InMux
    port map (
            O => \N__19460\,
            I => \N__19457\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__19457\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__1892\ : InMux
    port map (
            O => \N__19454\,
            I => \N__19451\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__19451\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__1890\ : InMux
    port map (
            O => \N__19448\,
            I => \N__19445\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__19445\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__1888\ : CascadeMux
    port map (
            O => \N__19442\,
            I => \N__19439\
        );

    \I__1887\ : InMux
    port map (
            O => \N__19439\,
            I => \N__19436\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__19436\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__1885\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19430\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__19430\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__19427\,
            I => \N__19424\
        );

    \I__1882\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19421\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__19421\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__1880\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19415\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__19415\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__1878\ : InMux
    port map (
            O => \N__19412\,
            I => \N__19409\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__19409\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__1876\ : InMux
    port map (
            O => \N__19406\,
            I => \N__19403\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__19403\,
            I => \N__19400\
        );

    \I__1874\ : Span4Mux_v
    port map (
            O => \N__19400\,
            I => \N__19397\
        );

    \I__1873\ : Span4Mux_v
    port map (
            O => \N__19397\,
            I => \N__19394\
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__19394\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__19391\,
            I => \N__19388\
        );

    \I__1870\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__19385\,
            I => \N__19382\
        );

    \I__1868\ : Span4Mux_v
    port map (
            O => \N__19382\,
            I => \N__19379\
        );

    \I__1867\ : Odrv4
    port map (
            O => \N__19379\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\
        );

    \I__1866\ : InMux
    port map (
            O => \N__19376\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__1865\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__19370\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__1862\ : InMux
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__19361\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__1859\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19352\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__19349\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__1856\ : InMux
    port map (
            O => \N__19346\,
            I => \N__19343\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__19343\,
            I => \N__19340\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__19340\,
            I => \N_38_i_i\
        );

    \I__1853\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19334\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__19334\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__1851\ : InMux
    port map (
            O => \N__19331\,
            I => \N__19328\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__19328\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__19325\,
            I => \N__19322\
        );

    \I__1848\ : InMux
    port map (
            O => \N__19322\,
            I => \N__19319\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__19316\,
            I => \N__19313\
        );

    \I__1845\ : Odrv4
    port map (
            O => \N__19313\,
            I => \current_shift_inst.PI_CTRL.integrator_1_23\
        );

    \I__1844\ : InMux
    port map (
            O => \N__19310\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__1843\ : InMux
    port map (
            O => \N__19307\,
            I => \N__19304\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__19304\,
            I => \N__19301\
        );

    \I__1841\ : Span4Mux_v
    port map (
            O => \N__19301\,
            I => \N__19298\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__19298\,
            I => \current_shift_inst.PI_CTRL.integrator_1_24\
        );

    \I__1839\ : InMux
    port map (
            O => \N__19295\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__1837\ : InMux
    port map (
            O => \N__19289\,
            I => \N__19286\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__19286\,
            I => \N__19283\
        );

    \I__1835\ : Span4Mux_h
    port map (
            O => \N__19283\,
            I => \N__19280\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__19280\,
            I => \N__19277\
        );

    \I__1833\ : Odrv4
    port map (
            O => \N__19277\,
            I => \current_shift_inst.PI_CTRL.integrator_1_25\
        );

    \I__1832\ : InMux
    port map (
            O => \N__19274\,
            I => \bfn_3_16_0_\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__19271\,
            I => \N__19268\
        );

    \I__1830\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__19265\,
            I => \N__19262\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__19262\,
            I => \N__19259\
        );

    \I__1827\ : Odrv4
    port map (
            O => \N__19259\,
            I => \current_shift_inst.PI_CTRL.integrator_1_26\
        );

    \I__1826\ : InMux
    port map (
            O => \N__19256\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__19253\,
            I => \N__19250\
        );

    \I__1824\ : InMux
    port map (
            O => \N__19250\,
            I => \N__19247\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__19247\,
            I => \N__19244\
        );

    \I__1822\ : Span4Mux_h
    port map (
            O => \N__19244\,
            I => \N__19241\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__19241\,
            I => \N__19238\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__19238\,
            I => \current_shift_inst.PI_CTRL.integrator_1_27\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__1818\ : InMux
    port map (
            O => \N__19232\,
            I => \N__19229\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__19229\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__1816\ : InMux
    port map (
            O => \N__19226\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__1814\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19217\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__19217\,
            I => \N__19214\
        );

    \I__1812\ : Span4Mux_h
    port map (
            O => \N__19214\,
            I => \N__19211\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__19211\,
            I => \N__19208\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__19208\,
            I => \current_shift_inst.PI_CTRL.integrator_1_28\
        );

    \I__1809\ : InMux
    port map (
            O => \N__19205\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__19202\,
            I => \N__19199\
        );

    \I__1807\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19196\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__19193\,
            I => \N__19190\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__19190\,
            I => \current_shift_inst.PI_CTRL.integrator_1_29\
        );

    \I__1803\ : InMux
    port map (
            O => \N__19187\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__1802\ : InMux
    port map (
            O => \N__19184\,
            I => \N__19181\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__19181\,
            I => \N__19178\
        );

    \I__1800\ : Span4Mux_v
    port map (
            O => \N__19178\,
            I => \N__19175\
        );

    \I__1799\ : Odrv4
    port map (
            O => \N__19175\,
            I => \current_shift_inst.PI_CTRL.integrator_1_30\
        );

    \I__1798\ : InMux
    port map (
            O => \N__19172\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__19169\,
            I => \N__19166\
        );

    \I__1796\ : InMux
    port map (
            O => \N__19166\,
            I => \N__19163\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__19163\,
            I => \N__19160\
        );

    \I__1794\ : Span4Mux_h
    port map (
            O => \N__19160\,
            I => \N__19157\
        );

    \I__1793\ : Odrv4
    port map (
            O => \N__19157\,
            I => \current_shift_inst.PI_CTRL.integrator_1_14\
        );

    \I__1792\ : InMux
    port map (
            O => \N__19154\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__1791\ : CascadeMux
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__1790\ : InMux
    port map (
            O => \N__19148\,
            I => \N__19145\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__19145\,
            I => \N__19142\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__19142\,
            I => \N__19139\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__19139\,
            I => \current_shift_inst.PI_CTRL.integrator_1_15\
        );

    \I__1786\ : InMux
    port map (
            O => \N__19136\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__19133\,
            I => \N__19130\
        );

    \I__1784\ : InMux
    port map (
            O => \N__19130\,
            I => \N__19127\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__19127\,
            I => \N__19124\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__19124\,
            I => \N__19121\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__19121\,
            I => \current_shift_inst.PI_CTRL.integrator_1_16\
        );

    \I__1780\ : InMux
    port map (
            O => \N__19118\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__19115\,
            I => \N__19112\
        );

    \I__1778\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__19109\,
            I => \N__19106\
        );

    \I__1776\ : Span4Mux_h
    port map (
            O => \N__19106\,
            I => \N__19103\
        );

    \I__1775\ : Span4Mux_v
    port map (
            O => \N__19103\,
            I => \N__19100\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__19100\,
            I => \current_shift_inst.PI_CTRL.integrator_1_17\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19097\,
            I => \bfn_3_15_0_\
        );

    \I__1772\ : CascadeMux
    port map (
            O => \N__19094\,
            I => \N__19091\
        );

    \I__1771\ : InMux
    port map (
            O => \N__19091\,
            I => \N__19088\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__19088\,
            I => \N__19085\
        );

    \I__1769\ : Span4Mux_v
    port map (
            O => \N__19085\,
            I => \N__19082\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__19082\,
            I => \current_shift_inst.PI_CTRL.integrator_1_18\
        );

    \I__1767\ : InMux
    port map (
            O => \N__19079\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__19076\,
            I => \N__19073\
        );

    \I__1765\ : InMux
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__1763\ : Span4Mux_h
    port map (
            O => \N__19067\,
            I => \N__19064\
        );

    \I__1762\ : Span4Mux_v
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__19061\,
            I => \current_shift_inst.PI_CTRL.integrator_1_19\
        );

    \I__1760\ : InMux
    port map (
            O => \N__19058\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__19055\,
            I => \N__19052\
        );

    \I__1758\ : InMux
    port map (
            O => \N__19052\,
            I => \N__19049\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__19049\,
            I => \N__19046\
        );

    \I__1756\ : Span12Mux_h
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__1755\ : Odrv12
    port map (
            O => \N__19043\,
            I => \current_shift_inst.PI_CTRL.integrator_1_20\
        );

    \I__1754\ : InMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__19037\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__1752\ : InMux
    port map (
            O => \N__19034\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__19031\,
            I => \N__19028\
        );

    \I__1750\ : InMux
    port map (
            O => \N__19028\,
            I => \N__19025\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__19025\,
            I => \N__19022\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__19022\,
            I => \N__19019\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__19019\,
            I => \current_shift_inst.PI_CTRL.integrator_1_21\
        );

    \I__1746\ : InMux
    port map (
            O => \N__19016\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__19013\,
            I => \N__19010\
        );

    \I__1744\ : InMux
    port map (
            O => \N__19010\,
            I => \N__19007\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__19007\,
            I => \N__19004\
        );

    \I__1742\ : Span4Mux_v
    port map (
            O => \N__19004\,
            I => \N__19001\
        );

    \I__1741\ : Odrv4
    port map (
            O => \N__19001\,
            I => \current_shift_inst.PI_CTRL.integrator_1_22\
        );

    \I__1740\ : InMux
    port map (
            O => \N__18998\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__18995\,
            I => \N__18992\
        );

    \I__1738\ : InMux
    port map (
            O => \N__18992\,
            I => \N__18989\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__18989\,
            I => \N__18986\
        );

    \I__1736\ : Span4Mux_h
    port map (
            O => \N__18986\,
            I => \N__18983\
        );

    \I__1735\ : Odrv4
    port map (
            O => \N__18983\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__1734\ : InMux
    port map (
            O => \N__18980\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__18977\,
            I => \N__18974\
        );

    \I__1732\ : InMux
    port map (
            O => \N__18974\,
            I => \N__18971\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__18971\,
            I => \N__18968\
        );

    \I__1730\ : Span4Mux_h
    port map (
            O => \N__18968\,
            I => \N__18965\
        );

    \I__1729\ : Odrv4
    port map (
            O => \N__18965\,
            I => \current_shift_inst.PI_CTRL.integrator_1_7\
        );

    \I__1728\ : InMux
    port map (
            O => \N__18962\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__18959\,
            I => \N__18956\
        );

    \I__1726\ : InMux
    port map (
            O => \N__18956\,
            I => \N__18953\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__18953\,
            I => \N__18950\
        );

    \I__1724\ : Span4Mux_h
    port map (
            O => \N__18950\,
            I => \N__18947\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__18947\,
            I => \current_shift_inst.PI_CTRL.integrator_1_8\
        );

    \I__1722\ : InMux
    port map (
            O => \N__18944\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__18941\,
            I => \N__18938\
        );

    \I__1720\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18935\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__18935\,
            I => \N__18932\
        );

    \I__1718\ : Span4Mux_v
    port map (
            O => \N__18932\,
            I => \N__18929\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__18929\,
            I => \current_shift_inst.PI_CTRL.integrator_1_9\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__18926\,
            I => \N__18923\
        );

    \I__1715\ : InMux
    port map (
            O => \N__18923\,
            I => \N__18920\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__18920\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__1713\ : InMux
    port map (
            O => \N__18917\,
            I => \bfn_3_14_0_\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__18914\,
            I => \N__18911\
        );

    \I__1711\ : InMux
    port map (
            O => \N__18911\,
            I => \N__18908\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__18908\,
            I => \N__18905\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__18905\,
            I => \N__18902\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__18902\,
            I => \current_shift_inst.PI_CTRL.integrator_1_10\
        );

    \I__1707\ : InMux
    port map (
            O => \N__18899\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__1705\ : InMux
    port map (
            O => \N__18893\,
            I => \N__18890\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__1703\ : Span4Mux_v
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__18884\,
            I => \current_shift_inst.PI_CTRL.integrator_1_11\
        );

    \I__1701\ : InMux
    port map (
            O => \N__18881\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__1700\ : InMux
    port map (
            O => \N__18878\,
            I => \N__18875\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__18875\,
            I => \N__18872\
        );

    \I__1698\ : Span4Mux_h
    port map (
            O => \N__18872\,
            I => \N__18869\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__18869\,
            I => \current_shift_inst.PI_CTRL.integrator_1_12\
        );

    \I__1696\ : InMux
    port map (
            O => \N__18866\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__1695\ : CascadeMux
    port map (
            O => \N__18863\,
            I => \N__18860\
        );

    \I__1694\ : InMux
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__18857\,
            I => \N__18854\
        );

    \I__1692\ : Span4Mux_h
    port map (
            O => \N__18854\,
            I => \N__18851\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__18851\,
            I => \current_shift_inst.PI_CTRL.integrator_1_13\
        );

    \I__1690\ : InMux
    port map (
            O => \N__18848\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__1689\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__18842\,
            I => \N__18839\
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__18839\,
            I => \rgb_drv_RNOZ0\
        );

    \I__1686\ : ClkMux
    port map (
            O => \N__18836\,
            I => \N__18830\
        );

    \I__1685\ : ClkMux
    port map (
            O => \N__18835\,
            I => \N__18830\
        );

    \I__1684\ : GlobalMux
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__1683\ : gio2CtrlBuf
    port map (
            O => \N__18827\,
            I => delay_hc_input_c_g
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__1681\ : InMux
    port map (
            O => \N__18821\,
            I => \N__18817\
        );

    \I__1680\ : InMux
    port map (
            O => \N__18820\,
            I => \N__18814\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__18817\,
            I => \N__18809\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__18814\,
            I => \N__18809\
        );

    \I__1677\ : Span4Mux_v
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__18806\,
            I => \current_shift_inst.PI_CTRL.un1_integrator\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__18803\,
            I => \N__18800\
        );

    \I__1674\ : InMux
    port map (
            O => \N__18800\,
            I => \N__18797\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__18791\,
            I => \current_shift_inst.PI_CTRL.integrator_1_2\
        );

    \I__1670\ : InMux
    port map (
            O => \N__18788\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__1668\ : InMux
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__18779\,
            I => \N__18776\
        );

    \I__1666\ : Span4Mux_v
    port map (
            O => \N__18776\,
            I => \N__18773\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__18773\,
            I => \current_shift_inst.PI_CTRL.integrator_1_3\
        );

    \I__1664\ : InMux
    port map (
            O => \N__18770\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__18767\,
            I => \N__18764\
        );

    \I__1662\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18761\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__18761\,
            I => \N__18758\
        );

    \I__1660\ : Span4Mux_v
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__18755\,
            I => \current_shift_inst.PI_CTRL.integrator_1_4\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__18752\,
            I => \N__18749\
        );

    \I__1657\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18746\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__18746\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__1655\ : InMux
    port map (
            O => \N__18743\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__18740\,
            I => \N__18737\
        );

    \I__1653\ : InMux
    port map (
            O => \N__18737\,
            I => \N__18734\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__18734\,
            I => \N__18731\
        );

    \I__1651\ : Span4Mux_h
    port map (
            O => \N__18731\,
            I => \N__18728\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__18728\,
            I => \current_shift_inst.PI_CTRL.integrator_1_5\
        );

    \I__1649\ : InMux
    port map (
            O => \N__18725\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__1648\ : InMux
    port map (
            O => \N__18722\,
            I => \N__18719\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__18719\,
            I => \N__18716\
        );

    \I__1646\ : Span4Mux_v
    port map (
            O => \N__18716\,
            I => \N__18713\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__18713\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_11\
        );

    \I__1644\ : InMux
    port map (
            O => \N__18710\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\
        );

    \I__1643\ : InMux
    port map (
            O => \N__18707\,
            I => \N__18704\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__18704\,
            I => \N__18701\
        );

    \I__1641\ : Span4Mux_v
    port map (
            O => \N__18701\,
            I => \N__18698\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__18698\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_12\
        );

    \I__1639\ : InMux
    port map (
            O => \N__18695\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\
        );

    \I__1638\ : InMux
    port map (
            O => \N__18692\,
            I => \N__18689\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__18689\,
            I => \N__18686\
        );

    \I__1636\ : Span4Mux_v
    port map (
            O => \N__18686\,
            I => \N__18683\
        );

    \I__1635\ : Odrv4
    port map (
            O => \N__18683\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_13\
        );

    \I__1634\ : InMux
    port map (
            O => \N__18680\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\
        );

    \I__1633\ : InMux
    port map (
            O => \N__18677\,
            I => \N__18674\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__1631\ : Span4Mux_v
    port map (
            O => \N__18671\,
            I => \N__18668\
        );

    \I__1630\ : Odrv4
    port map (
            O => \N__18668\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_14\
        );

    \I__1629\ : InMux
    port map (
            O => \N__18665\,
            I => \N__18651\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__18664\,
            I => \N__18648\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__18663\,
            I => \N__18645\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__18662\,
            I => \N__18642\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__18661\,
            I => \N__18639\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__18660\,
            I => \N__18636\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__18659\,
            I => \N__18633\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__18658\,
            I => \N__18630\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__18657\,
            I => \N__18627\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__18656\,
            I => \N__18624\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__18655\,
            I => \N__18621\
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__18654\,
            I => \N__18618\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__18651\,
            I => \N__18615\
        );

    \I__1616\ : InMux
    port map (
            O => \N__18648\,
            I => \N__18608\
        );

    \I__1615\ : InMux
    port map (
            O => \N__18645\,
            I => \N__18608\
        );

    \I__1614\ : InMux
    port map (
            O => \N__18642\,
            I => \N__18608\
        );

    \I__1613\ : InMux
    port map (
            O => \N__18639\,
            I => \N__18599\
        );

    \I__1612\ : InMux
    port map (
            O => \N__18636\,
            I => \N__18599\
        );

    \I__1611\ : InMux
    port map (
            O => \N__18633\,
            I => \N__18599\
        );

    \I__1610\ : InMux
    port map (
            O => \N__18630\,
            I => \N__18599\
        );

    \I__1609\ : InMux
    port map (
            O => \N__18627\,
            I => \N__18594\
        );

    \I__1608\ : InMux
    port map (
            O => \N__18624\,
            I => \N__18594\
        );

    \I__1607\ : InMux
    port map (
            O => \N__18621\,
            I => \N__18589\
        );

    \I__1606\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18589\
        );

    \I__1605\ : Odrv4
    port map (
            O => \N__18615\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__18608\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__18599\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__18594\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__18589\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1600\ : InMux
    port map (
            O => \N__18578\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\
        );

    \I__1599\ : InMux
    port map (
            O => \N__18575\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\
        );

    \I__1598\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18569\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__18569\,
            I => \N__18566\
        );

    \I__1596\ : Span4Mux_v
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__18563\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_3\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__18560\,
            I => \N__18557\
        );

    \I__1593\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__18554\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_18\
        );

    \I__1591\ : InMux
    port map (
            O => \N__18551\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\
        );

    \I__1590\ : InMux
    port map (
            O => \N__18548\,
            I => \N__18545\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__18545\,
            I => \N__18542\
        );

    \I__1588\ : Span4Mux_v
    port map (
            O => \N__18542\,
            I => \N__18539\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__18539\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_4\
        );

    \I__1586\ : InMux
    port map (
            O => \N__18536\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\
        );

    \I__1585\ : InMux
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__1583\ : Span4Mux_v
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__18524\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_5\
        );

    \I__1581\ : InMux
    port map (
            O => \N__18521\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\
        );

    \I__1580\ : InMux
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__1578\ : Span4Mux_v
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__18509\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_6\
        );

    \I__1576\ : InMux
    port map (
            O => \N__18506\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\
        );

    \I__1575\ : InMux
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__1573\ : Span4Mux_v
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__1572\ : Odrv4
    port map (
            O => \N__18494\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_7\
        );

    \I__1571\ : InMux
    port map (
            O => \N__18491\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\
        );

    \I__1570\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18485\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__18485\,
            I => \N__18482\
        );

    \I__1568\ : Span4Mux_v
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__18479\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_8\
        );

    \I__1566\ : InMux
    port map (
            O => \N__18476\,
            I => \bfn_1_12_0_\
        );

    \I__1565\ : InMux
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__18470\,
            I => \N__18467\
        );

    \I__1563\ : Span4Mux_v
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__1562\ : Odrv4
    port map (
            O => \N__18464\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_9\
        );

    \I__1561\ : InMux
    port map (
            O => \N__18461\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\
        );

    \I__1560\ : InMux
    port map (
            O => \N__18458\,
            I => \N__18455\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__18455\,
            I => \N__18452\
        );

    \I__1558\ : Span4Mux_v
    port map (
            O => \N__18452\,
            I => \N__18449\
        );

    \I__1557\ : Odrv4
    port map (
            O => \N__18449\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_10\
        );

    \I__1556\ : InMux
    port map (
            O => \N__18446\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\
        );

    \I__1555\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__18440\,
            I => \N__18437\
        );

    \I__1553\ : Span4Mux_v
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__18434\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_15\
        );

    \I__1551\ : InMux
    port map (
            O => \N__18431\,
            I => \N__18428\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__18428\,
            I => \N__18425\
        );

    \I__1549\ : Span4Mux_v
    port map (
            O => \N__18425\,
            I => \N__18422\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__18422\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_0\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__1546\ : InMux
    port map (
            O => \N__18416\,
            I => \N__18413\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__18413\,
            I => \N__18410\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__18410\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_15\
        );

    \I__1543\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18404\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__1541\ : Span4Mux_v
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__18398\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_1\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__1538\ : InMux
    port map (
            O => \N__18392\,
            I => \N__18389\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__18389\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_16\
        );

    \I__1536\ : InMux
    port map (
            O => \N__18386\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\
        );

    \I__1535\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18380\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__18380\,
            I => \N__18377\
        );

    \I__1533\ : Span4Mux_v
    port map (
            O => \N__18377\,
            I => \N__18374\
        );

    \I__1532\ : Odrv4
    port map (
            O => \N__18374\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_2\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__18371\,
            I => \N__18368\
        );

    \I__1530\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18365\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__18365\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_17\
        );

    \I__1528\ : InMux
    port map (
            O => \N__18362\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\
        );

    \I__1527\ : IoInMux
    port map (
            O => \N__18359\,
            I => \N__18356\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__18356\,
            I => \N__18353\
        );

    \I__1525\ : Span4Mux_s1_v
    port map (
            O => \N__18353\,
            I => \N__18350\
        );

    \I__1524\ : Span4Mux_h
    port map (
            O => \N__18350\,
            I => \N__18347\
        );

    \I__1523\ : Sp12to4
    port map (
            O => \N__18347\,
            I => \N__18344\
        );

    \I__1522\ : Span12Mux_s9_v
    port map (
            O => \N__18344\,
            I => \N__18341\
        );

    \I__1521\ : Span12Mux_v
    port map (
            O => \N__18341\,
            I => \N__18338\
        );

    \I__1520\ : Odrv12
    port map (
            O => \N__18338\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1519\ : IoInMux
    port map (
            O => \N__18335\,
            I => \N__18332\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__18332\,
            I => \N__18329\
        );

    \I__1517\ : IoSpan4Mux
    port map (
            O => \N__18329\,
            I => \N__18326\
        );

    \I__1516\ : IoSpan4Mux
    port map (
            O => \N__18326\,
            I => \N__18323\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__18323\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_14_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_28_0_\
        );

    \IN_MUX_bfv_14_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_7\,
            carryinitout => \bfn_14_29_0_\
        );

    \IN_MUX_bfv_14_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_15\,
            carryinitout => \bfn_14_30_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_12_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_12_7_0_\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_12_8_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_3_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_13_0_\
        );

    \IN_MUX_bfv_3_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryinitout => \bfn_3_14_0_\
        );

    \IN_MUX_bfv_3_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryinitout => \bfn_3_15_0_\
        );

    \IN_MUX_bfv_3_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryinitout => \bfn_3_16_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_15_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryinitout => \bfn_15_24_0_\
        );

    \IN_MUX_bfv_15_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryinitout => \bfn_15_25_0_\
        );

    \IN_MUX_bfv_15_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryinitout => \bfn_15_26_0_\
        );

    \IN_MUX_bfv_13_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_28_0_\
        );

    \IN_MUX_bfv_13_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            carryinitout => \bfn_13_29_0_\
        );

    \IN_MUX_bfv_13_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            carryinitout => \bfn_13_30_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_13_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_cry_7\,
            carryinitout => \bfn_13_25_0_\
        );

    \IN_MUX_bfv_14_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_25_0_\
        );

    \IN_MUX_bfv_14_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_7\,
            carryinitout => \bfn_14_26_0_\
        );

    \IN_MUX_bfv_14_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_15\,
            carryinitout => \bfn_14_27_0_\
        );

    \IN_MUX_bfv_11_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_23_0_\
        );

    \IN_MUX_bfv_11_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_11_24_0_\
        );

    \IN_MUX_bfv_12_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_21_0_\
        );

    \IN_MUX_bfv_12_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_12_22_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_18_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_10_0_\
        );

    \IN_MUX_bfv_18_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_18_11_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_7_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_7_21_0_\
        );

    \IN_MUX_bfv_7_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_7_22_0_\
        );

    \IN_MUX_bfv_7_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_7_23_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_10_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_10_20_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_8_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_8_21_0_\
        );

    \IN_MUX_bfv_8_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_8_22_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_7_14_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18359\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18335\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__32600\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_162_i_g\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__36125\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__26204\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__37792\,
            CLKHFEN => \N__37794\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__37793\,
            RGB2PWM => \N__19346\,
            RGB1 => rgb_g_wire,
            CURREN => \N__37913\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__18845\,
            RGB0PWM => \N__48311\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18443\,
            in2 => \_gnd_net_\,
            in3 => \N__18665\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18431\,
            in2 => \N__18419\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_16\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18407\,
            in2 => \N__18395\,
            in3 => \N__18386\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18383\,
            in2 => \N__18371\,
            in3 => \N__18362\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18572\,
            in2 => \N__18560\,
            in3 => \N__18551\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18548\,
            in2 => \N__18654\,
            in3 => \N__18536\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18533\,
            in2 => \N__18656\,
            in3 => \N__18521\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18518\,
            in2 => \N__18655\,
            in3 => \N__18506\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18503\,
            in2 => \N__18657\,
            in3 => \N__18491\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18488\,
            in2 => \N__18658\,
            in3 => \N__18476\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_24\,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18473\,
            in2 => \N__18662\,
            in3 => \N__18461\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18458\,
            in2 => \N__18659\,
            in3 => \N__18446\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18722\,
            in2 => \N__18663\,
            in3 => \N__18710\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18707\,
            in2 => \N__18660\,
            in3 => \N__18695\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18692\,
            in2 => \N__18664\,
            in3 => \N__18680\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18677\,
            in2 => \N__18661\,
            in3 => \N__18578\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18575\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29142\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18836\,
            ce => 'H',
            sr => \N__48255\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__41042\,
            in1 => \N__20008\,
            in2 => \N__18752\,
            in3 => \N__19815\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48794\,
            ce => 'H',
            sr => \N__48261\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101001001000"
        )
    port map (
            in0 => \N__39835\,
            in1 => \N__20009\,
            in2 => \N__18824\,
            in3 => \N__19830\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48785\,
            ce => 'H',
            sr => \N__48264\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000010110001"
        )
    port map (
            in0 => \N__20001\,
            in1 => \N__41041\,
            in2 => \N__18926\,
            in3 => \N__19802\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48773\,
            ce => 'H',
            sr => \N__48268\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__20000\,
            in1 => \N__41040\,
            in2 => \N__19829\,
            in3 => \N__19040\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48773\,
            ce => 'H',
            sr => \N__48268\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__19998\,
            in1 => \N__41046\,
            in2 => \N__19235\,
            in3 => \N__19814\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48755\,
            ce => 'H',
            sr => \N__48277\
        );

    \rgb_drv_RNO_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__43025\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48310\,
            lcout => \rgb_drv_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29143\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18835\,
            ce => 'H',
            sr => \N__48247\
        );

    \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18820\,
            in2 => \N__39857\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39786\,
            in2 => \N__18803\,
            in3 => \N__18788\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39729\,
            in2 => \N__18785\,
            in3 => \N__18770\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39666\,
            in2 => \N__18767\,
            in3 => \N__18743\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39638\,
            in2 => \N__18740\,
            in3 => \N__18725\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39557\,
            in2 => \N__18995\,
            in3 => \N__18980\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39512\,
            in2 => \N__18977\,
            in3 => \N__18962\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39458\,
            in2 => \N__18959\,
            in3 => \N__18944\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40302\,
            in2 => \N__18941\,
            in3 => \N__18917\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_3_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40254\,
            in2 => \N__18914\,
            in3 => \N__18899\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40181\,
            in2 => \N__18896\,
            in3 => \N__18881\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18878\,
            in2 => \N__40118\,
            in3 => \N__18866\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40067\,
            in2 => \N__18863\,
            in3 => \N__18848\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40021\,
            in2 => \N__19169\,
            in3 => \N__19154\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39965\,
            in2 => \N__19151\,
            in3 => \N__19136\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39920\,
            in2 => \N__19133\,
            in3 => \N__19118\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40709\,
            in2 => \N__19115\,
            in3 => \N__19097\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_3_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40665\,
            in2 => \N__19094\,
            in3 => \N__19079\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40604\,
            in2 => \N__19076\,
            in3 => \N__19058\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40550\,
            in2 => \N__19055\,
            in3 => \N__19034\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40514\,
            in2 => \N__19031\,
            in3 => \N__19016\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40469\,
            in2 => \N__19013\,
            in3 => \N__18998\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40412\,
            in2 => \N__19325\,
            in3 => \N__19310\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19307\,
            in2 => \N__40379\,
            in3 => \N__19295\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41297\,
            in2 => \N__19292\,
            in3 => \N__19274\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_3_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41258\,
            in2 => \N__19271\,
            in3 => \N__19256\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41211\,
            in2 => \N__19253\,
            in3 => \N__19226\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41169\,
            in2 => \N__19223\,
            in3 => \N__19205\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41120\,
            in2 => \N__19202\,
            in3 => \N__19187\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19184\,
            in2 => \N__41088\,
            in3 => \N__19172\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__40971\,
            in1 => \N__19406\,
            in2 => \N__19391\,
            in3 => \N__19376\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000100010"
        )
    port map (
            in0 => \N__41008\,
            in1 => \N__19927\,
            in2 => \N__19806\,
            in3 => \N__19373\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48742\,
            ce => 'H',
            sr => \N__48273\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__19926\,
            in1 => \N__41010\,
            in2 => \N__19367\,
            in3 => \N__19748\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48742\,
            ce => 'H',
            sr => \N__48273\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__19925\,
            in1 => \N__41009\,
            in2 => \N__19358\,
            in3 => \N__19747\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48742\,
            ce => 'H',
            sr => \N__48273\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41304\,
            in1 => \N__41207\,
            in2 => \N__41270\,
            in3 => \N__41168\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40614\,
            in1 => \N__40661\,
            in2 => \N__40725\,
            in3 => \N__40477\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_0_LC_3_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__48309\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43024\,
            lcout => \N_38_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__19981\,
            in1 => \N__19823\,
            in2 => \_gnd_net_\,
            in3 => \N__19337\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48774\,
            ce => 'H',
            sr => \N__48248\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101000"
        )
    port map (
            in0 => \N__19331\,
            in1 => \N__19980\,
            in2 => \N__19832\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48774\,
            ce => 'H',
            sr => \N__48248\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111100000001"
        )
    port map (
            in0 => \N__19982\,
            in1 => \N__19824\,
            in2 => \N__41050\,
            in3 => \N__19466\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48774\,
            ce => 'H',
            sr => \N__48248\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100000001"
        )
    port map (
            in0 => \N__19978\,
            in1 => \N__41033\,
            in2 => \N__19821\,
            in3 => \N__19460\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48765\,
            ce => 'H',
            sr => \N__48256\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__19977\,
            in1 => \N__41032\,
            in2 => \N__19820\,
            in3 => \N__19454\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48765\,
            ce => 'H',
            sr => \N__48256\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100000001"
        )
    port map (
            in0 => \N__19979\,
            in1 => \N__41034\,
            in2 => \N__19822\,
            in3 => \N__19448\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48765\,
            ce => 'H',
            sr => \N__48256\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__41031\,
            in1 => \N__19976\,
            in2 => \N__19442\,
            in3 => \N__19788\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48765\,
            ce => 'H',
            sr => \N__48256\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__19965\,
            in1 => \N__41004\,
            in2 => \N__19817\,
            in3 => \N__19433\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48756\,
            ce => 'H',
            sr => \N__48262\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__41002\,
            in1 => \N__19968\,
            in2 => \N__19427\,
            in3 => \N__19778\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48756\,
            ce => 'H',
            sr => \N__48262\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__19967\,
            in1 => \N__41005\,
            in2 => \N__19818\,
            in3 => \N__19418\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48756\,
            ce => 'H',
            sr => \N__48262\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__19969\,
            in1 => \N__41006\,
            in2 => \N__19819\,
            in3 => \N__19412\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48756\,
            ce => 'H',
            sr => \N__48262\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__41000\,
            in1 => \N__19776\,
            in2 => \N__19538\,
            in3 => \N__19963\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48756\,
            ce => 'H',
            sr => \N__48262\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__19964\,
            in1 => \N__41003\,
            in2 => \N__19816\,
            in3 => \N__19529\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48756\,
            ce => 'H',
            sr => \N__48262\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__41001\,
            in1 => \N__19966\,
            in2 => \N__19523\,
            in3 => \N__19777\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48756\,
            ce => 'H',
            sr => \N__48262\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__40995\,
            in1 => \N__19958\,
            in2 => \N__19514\,
            in3 => \N__19739\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48743\,
            ce => 'H',
            sr => \N__48265\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__40997\,
            in1 => \N__19740\,
            in2 => \N__19502\,
            in3 => \N__19961\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48743\,
            ce => 'H',
            sr => \N__48265\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__19962\,
            in1 => \N__40998\,
            in2 => \N__19804\,
            in3 => \N__19493\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48743\,
            ce => 'H',
            sr => \N__48265\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111001000"
        )
    port map (
            in0 => \N__19960\,
            in1 => \N__19487\,
            in2 => \N__19803\,
            in3 => \N__40999\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48743\,
            ce => 'H',
            sr => \N__48265\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__40996\,
            in1 => \N__19959\,
            in2 => \N__19481\,
            in3 => \N__19738\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48743\,
            ce => 'H',
            sr => \N__48265\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__19895\,
            in1 => \N__41011\,
            in2 => \N__19807\,
            in3 => \N__19472\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48732\,
            ce => 'H',
            sr => \N__48269\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39966\,
            in1 => \N__40250\,
            in2 => \N__40081\,
            in3 => \N__39925\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__40194\,
            in1 => \N__40020\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40129\,
            in1 => \N__19574\,
            in2 => \N__19568\,
            in3 => \N__41078\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20099\,
            in1 => \N__19565\,
            in2 => \N__19559\,
            in3 => \N__19544\,
            lcout => \current_shift_inst.PI_CTRL.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39519\,
            in1 => \N__39472\,
            in2 => \N__39581\,
            in3 => \N__40323\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__39645\,
            in1 => \N__39690\,
            in2 => \N__19556\,
            in3 => \N__39748\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__41136\,
            in1 => \N__40413\,
            in2 => \N__19553\,
            in3 => \N__19550\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39921\,
            in1 => \N__40016\,
            in2 => \N__40198\,
            in3 => \N__40128\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41259\,
            in2 => \_gnd_net_\,
            in3 => \N__40515\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41179\,
            in1 => \N__41224\,
            in2 => \N__41314\,
            in3 => \N__41092\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40560\,
            in1 => \N__40383\,
            in2 => \N__19616\,
            in3 => \N__19613\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__40615\,
            in1 => \N__40669\,
            in2 => \N__40735\,
            in3 => \N__40473\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__41013\,
            in1 => \N__40420\,
            in2 => \N__19607\,
            in3 => \N__19604\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20093\,
            in1 => \N__19598\,
            in2 => \N__19592\,
            in3 => \N__19580\,
            lcout => \current_shift_inst.PI_CTRL.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__39523\,
            in1 => \N__39647\,
            in2 => \_gnd_net_\,
            in3 => \N__39471\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110111"
        )
    port map (
            in0 => \N__39796\,
            in1 => \N__39747\,
            in2 => \N__39877\,
            in3 => \N__39694\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__19589\,
            in1 => \N__40327\,
            in2 => \N__19583\,
            in3 => \N__39573\,
            lcout => \current_shift_inst.PI_CTRL.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23611\,
            in1 => \N__23589\,
            in2 => \_gnd_net_\,
            in3 => \N__41887\,
            lcout => \elapsed_time_ns_1_RNI7ADN9_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_29_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23610\,
            in1 => \N__23590\,
            in2 => \_gnd_net_\,
            in3 => \N__41816\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48804\,
            ce => \N__28504\,
            sr => \N__48215\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41884\,
            in1 => \N__23670\,
            in2 => \_gnd_net_\,
            in3 => \N__23650\,
            lcout => \elapsed_time_ns_1_RNIL73T9_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__28283\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28209\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23883\,
            in1 => \N__23864\,
            in2 => \_gnd_net_\,
            in3 => \N__41881\,
            lcout => \elapsed_time_ns_1_RNIDV2T9_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20055\,
            in1 => \N__20431\,
            in2 => \_gnd_net_\,
            in3 => \N__41883\,
            lcout => \elapsed_time_ns_1_RNIUVBN9_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31533\,
            in1 => \N__31503\,
            in2 => \_gnd_net_\,
            in3 => \N__41882\,
            lcout => \elapsed_time_ns_1_RNI03DN9_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_22_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41886\,
            in1 => \N__31534\,
            in2 => \_gnd_net_\,
            in3 => \N__31510\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48775\,
            ce => \N__28502\,
            sr => \N__48237\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41885\,
            in1 => \N__20056\,
            in2 => \_gnd_net_\,
            in3 => \N__20430\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48775\,
            ce => \N__28502\,
            sr => \N__48237\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011010001"
        )
    port map (
            in0 => \N__41036\,
            in1 => \N__19999\,
            in2 => \N__20033\,
            in3 => \N__19828\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48766\,
            ce => 'H',
            sr => \N__48242\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__41035\,
            in1 => \N__19997\,
            in2 => \N__20021\,
            in3 => \N__19831\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48757\,
            ce => 'H',
            sr => \N__48249\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__41007\,
            in1 => \N__19983\,
            in2 => \N__19847\,
            in3 => \N__19805\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48744\,
            ce => 'H',
            sr => \N__48257\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40384\,
            in1 => \N__40573\,
            in2 => \N__40529\,
            in3 => \N__41012\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39979\,
            in1 => \N__40080\,
            in2 => \N__40261\,
            in3 => \N__41140\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20087\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22971\,
            in1 => \N__24058\,
            in2 => \_gnd_net_\,
            in3 => \N__41878\,
            lcout => \elapsed_time_ns_1_RNI68CN9_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23938\,
            in1 => \N__23379\,
            in2 => \_gnd_net_\,
            in3 => \N__41898\,
            lcout => \elapsed_time_ns_1_RNI04EN9_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22972\,
            in1 => \N__24062\,
            in2 => \_gnd_net_\,
            in3 => \N__41899\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48799\,
            ce => \N__28508\,
            sr => \N__48191\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23736\,
            in1 => \N__23713\,
            in2 => \_gnd_net_\,
            in3 => \N__41814\,
            lcout => \elapsed_time_ns_1_RNITUBN9_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41815\,
            in1 => \N__20060\,
            in2 => \_gnd_net_\,
            in3 => \N__20432\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48795\,
            ce => \N__36595\,
            sr => \N__48201\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31612\,
            in1 => \N__31585\,
            in2 => \_gnd_net_\,
            in3 => \N__41861\,
            lcout => \elapsed_time_ns_1_RNI14DN9_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__22021\,
            in1 => \N__25963\,
            in2 => \N__25996\,
            in3 => \N__22000\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23239\,
            in2 => \_gnd_net_\,
            in3 => \N__25080\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24916\,
            in1 => \N__23162\,
            in2 => \N__20135\,
            in3 => \N__20132\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28706\,
            in1 => \N__28744\,
            in2 => \_gnd_net_\,
            in3 => \N__41903\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48776\,
            ce => \N__36444\,
            sr => \N__48216\
        );

    \phase_controller_inst2.state_RNIG7JF_2_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31768\,
            in2 => \_gnd_net_\,
            in3 => \N__31801\,
            lcout => \phase_controller_inst2.state_RNIG7JFZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20414\,
            in1 => \N__23699\,
            in2 => \N__28739\,
            in3 => \N__23636\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__20108\,
            in1 => \N__20122\,
            in2 => \N__25886\,
            in3 => \N__25859\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101010001"
        )
    port map (
            in0 => \N__25858\,
            in1 => \N__25885\,
            in2 => \N__20123\,
            in3 => \N__20107\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_23_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41901\,
            in1 => \N__31608\,
            in2 => \_gnd_net_\,
            in3 => \N__31574\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48758\,
            ce => \N__28503\,
            sr => \N__48227\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23643\,
            in1 => \N__23678\,
            in2 => \_gnd_net_\,
            in3 => \N__41902\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48758\,
            ce => \N__28503\,
            sr => \N__48227\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41900\,
            in1 => \N__23737\,
            in2 => \_gnd_net_\,
            in3 => \N__23703\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48758\,
            ce => \N__28503\,
            sr => \N__48227\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20162\,
            in2 => \_gnd_net_\,
            in3 => \N__22487\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22475\,
            in2 => \_gnd_net_\,
            in3 => \N__20156\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__48745\,
            ce => 'H',
            sr => \N__48232\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22454\,
            in2 => \_gnd_net_\,
            in3 => \N__20153\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__48745\,
            ce => 'H',
            sr => \N__48232\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22439\,
            in2 => \_gnd_net_\,
            in3 => \N__20150\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__48745\,
            ce => 'H',
            sr => \N__48232\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22418\,
            in2 => \_gnd_net_\,
            in3 => \N__20147\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__48745\,
            ce => 'H',
            sr => \N__48232\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22397\,
            in2 => \_gnd_net_\,
            in3 => \N__20144\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__48745\,
            ce => 'H',
            sr => \N__48232\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22376\,
            in2 => \_gnd_net_\,
            in3 => \N__20141\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__48745\,
            ce => 'H',
            sr => \N__48232\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22616\,
            in2 => \_gnd_net_\,
            in3 => \N__20138\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__48745\,
            ce => 'H',
            sr => \N__48232\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22601\,
            in2 => \_gnd_net_\,
            in3 => \N__20183\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__48733\,
            ce => 'H',
            sr => \N__48238\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22586\,
            in2 => \_gnd_net_\,
            in3 => \N__20180\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__48733\,
            ce => 'H',
            sr => \N__48238\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22571\,
            in2 => \_gnd_net_\,
            in3 => \N__20177\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__48733\,
            ce => 'H',
            sr => \N__48238\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22556\,
            in2 => \_gnd_net_\,
            in3 => \N__20174\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__48733\,
            ce => 'H',
            sr => \N__48238\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22535\,
            in2 => \_gnd_net_\,
            in3 => \N__20171\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__48733\,
            ce => 'H',
            sr => \N__48238\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21059\,
            in2 => \_gnd_net_\,
            in3 => \N__20168\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__48733\,
            ce => 'H',
            sr => \N__48238\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22517\,
            in2 => \_gnd_net_\,
            in3 => \N__20165\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48733\,
            ce => 'H',
            sr => \N__48238\
        );

    \phase_controller_inst2.state_1_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__27793\,
            in1 => \N__31830\,
            in2 => \_gnd_net_\,
            in3 => \N__31715\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48733\,
            ce => 'H',
            sr => \N__48238\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__26911\,
            in1 => \N__32143\,
            in2 => \_gnd_net_\,
            in3 => \N__32112\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__26910\,
            in1 => \N__33695\,
            in2 => \_gnd_net_\,
            in3 => \N__33649\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32400\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24231\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29784\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32652\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29600\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24421\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29519\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32318\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21255\,
            in2 => \N__21232\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_7_20_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__48684\,
            ce => \N__33740\,
            sr => \N__48270\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23955\,
            in2 => \N__21208\,
            in3 => \N__20210\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__48684\,
            ce => \N__33740\,
            sr => \N__48270\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21447\,
            in2 => \N__21233\,
            in3 => \N__20207\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__48684\,
            ce => \N__33740\,
            sr => \N__48270\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21423\,
            in2 => \N__21209\,
            in3 => \N__20204\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__48684\,
            ce => \N__33740\,
            sr => \N__48270\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21399\,
            in2 => \N__21452\,
            in3 => \N__20201\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__48684\,
            ce => \N__33740\,
            sr => \N__48270\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21375\,
            in2 => \N__21428\,
            in3 => \N__20198\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__48684\,
            ce => \N__33740\,
            sr => \N__48270\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21351\,
            in2 => \N__21404\,
            in3 => \N__20195\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__48684\,
            ce => \N__33740\,
            sr => \N__48270\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21327\,
            in2 => \N__21380\,
            in3 => \N__20192\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__48684\,
            ce => \N__33740\,
            sr => \N__48270\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21303\,
            in2 => \N__21356\,
            in3 => \N__20189\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_7_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__48679\,
            ce => \N__33739\,
            sr => \N__48274\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21279\,
            in2 => \N__21332\,
            in3 => \N__20186\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__48679\,
            ce => \N__33739\,
            sr => \N__48274\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21660\,
            in2 => \N__21308\,
            in3 => \N__20237\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__48679\,
            ce => \N__33739\,
            sr => \N__48274\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21636\,
            in2 => \N__21284\,
            in3 => \N__20234\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__48679\,
            ce => \N__33739\,
            sr => \N__48274\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21612\,
            in2 => \N__21665\,
            in3 => \N__20231\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__48679\,
            ce => \N__33739\,
            sr => \N__48274\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21588\,
            in2 => \N__21641\,
            in3 => \N__20228\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__48679\,
            ce => \N__33739\,
            sr => \N__48274\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21564\,
            in2 => \N__21617\,
            in3 => \N__20225\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__48679\,
            ce => \N__33739\,
            sr => \N__48274\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21540\,
            in2 => \N__21593\,
            in3 => \N__20222\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__48679\,
            ce => \N__33739\,
            sr => \N__48274\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21516\,
            in2 => \N__21569\,
            in3 => \N__20219\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_7_22_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__48675\,
            ce => \N__33738\,
            sr => \N__48278\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21492\,
            in2 => \N__21545\,
            in3 => \N__20216\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__48675\,
            ce => \N__33738\,
            sr => \N__48278\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21468\,
            in2 => \N__21521\,
            in3 => \N__20213\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__48675\,
            ce => \N__33738\,
            sr => \N__48278\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21843\,
            in2 => \N__21497\,
            in3 => \N__20264\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__48675\,
            ce => \N__33738\,
            sr => \N__48278\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21819\,
            in2 => \N__21473\,
            in3 => \N__20261\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__48675\,
            ce => \N__33738\,
            sr => \N__48278\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21795\,
            in2 => \N__21848\,
            in3 => \N__20258\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__48675\,
            ce => \N__33738\,
            sr => \N__48278\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21771\,
            in2 => \N__21824\,
            in3 => \N__20255\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__48675\,
            ce => \N__33738\,
            sr => \N__48278\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21747\,
            in2 => \N__21800\,
            in3 => \N__20252\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__48675\,
            ce => \N__33738\,
            sr => \N__48278\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21723\,
            in2 => \N__21776\,
            in3 => \N__20249\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_7_23_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__48669\,
            ce => \N__33737\,
            sr => \N__48281\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21699\,
            in2 => \N__21752\,
            in3 => \N__20246\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__48669\,
            ce => \N__33737\,
            sr => \N__48281\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21679\,
            in2 => \N__21728\,
            in3 => \N__20243\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__48669\,
            ce => \N__33737\,
            sr => \N__48281\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21904\,
            in2 => \N__21704\,
            in3 => \N__20240\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__48669\,
            ce => \N__33737\,
            sr => \N__48281\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20312\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20308\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48665\,
            ce => 'H',
            sr => \N__48282\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21869\,
            in1 => \N__23292\,
            in2 => \_gnd_net_\,
            in3 => \N__41890\,
            lcout => \elapsed_time_ns_1_RNI24CN9_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20282\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22948\,
            in1 => \N__24023\,
            in2 => \_gnd_net_\,
            in3 => \N__41825\,
            lcout => \elapsed_time_ns_1_RNI57CN9_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30725\,
            in1 => \N__30767\,
            in2 => \_gnd_net_\,
            in3 => \N__41833\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48800\,
            ce => \N__28511\,
            sr => \N__48173\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41832\,
            in1 => \N__22944\,
            in2 => \_gnd_net_\,
            in3 => \N__24021\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48800\,
            ce => \N__28511\,
            sr => \N__48173\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29116\,
            in1 => \N__21951\,
            in2 => \_gnd_net_\,
            in3 => \N__20273\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__48796\,
            ce => \N__29219\,
            sr => \N__48182\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29112\,
            in1 => \N__21927\,
            in2 => \_gnd_net_\,
            in3 => \N__20270\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__48796\,
            ce => \N__29219\,
            sr => \N__48182\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29117\,
            in1 => \N__20607\,
            in2 => \_gnd_net_\,
            in3 => \N__20267\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__48796\,
            ce => \N__29219\,
            sr => \N__48182\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29113\,
            in1 => \N__20581\,
            in2 => \_gnd_net_\,
            in3 => \N__20339\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__48796\,
            ce => \N__29219\,
            sr => \N__48182\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29118\,
            in1 => \N__20556\,
            in2 => \_gnd_net_\,
            in3 => \N__20336\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__48796\,
            ce => \N__29219\,
            sr => \N__48182\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29114\,
            in1 => \N__20529\,
            in2 => \_gnd_net_\,
            in3 => \N__20333\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__48796\,
            ce => \N__29219\,
            sr => \N__48182\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29119\,
            in1 => \N__20503\,
            in2 => \_gnd_net_\,
            in3 => \N__20330\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__48796\,
            ce => \N__29219\,
            sr => \N__48182\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29115\,
            in1 => \N__20479\,
            in2 => \_gnd_net_\,
            in3 => \N__20327\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__48796\,
            ce => \N__29219\,
            sr => \N__48182\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29111\,
            in1 => \N__20448\,
            in2 => \_gnd_net_\,
            in3 => \N__20324\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__48786\,
            ce => \N__29218\,
            sr => \N__48192\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29123\,
            in1 => \N__20829\,
            in2 => \_gnd_net_\,
            in3 => \N__20321\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__48786\,
            ce => \N__29218\,
            sr => \N__48192\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29108\,
            in1 => \N__20800\,
            in2 => \_gnd_net_\,
            in3 => \N__20318\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__48786\,
            ce => \N__29218\,
            sr => \N__48192\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29120\,
            in1 => \N__20781\,
            in2 => \_gnd_net_\,
            in3 => \N__20315\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__48786\,
            ce => \N__29218\,
            sr => \N__48192\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29109\,
            in1 => \N__20754\,
            in2 => \_gnd_net_\,
            in3 => \N__20366\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__48786\,
            ce => \N__29218\,
            sr => \N__48192\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29121\,
            in1 => \N__20727\,
            in2 => \_gnd_net_\,
            in3 => \N__20363\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__48786\,
            ce => \N__29218\,
            sr => \N__48192\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29110\,
            in1 => \N__20697\,
            in2 => \_gnd_net_\,
            in3 => \N__20360\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__48786\,
            ce => \N__29218\,
            sr => \N__48192\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29122\,
            in1 => \N__20667\,
            in2 => \_gnd_net_\,
            in3 => \N__20357\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__48786\,
            ce => \N__29218\,
            sr => \N__48192\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29100\,
            in1 => \N__20643\,
            in2 => \_gnd_net_\,
            in3 => \N__20354\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__48777\,
            ce => \N__29217\,
            sr => \N__48202\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29104\,
            in1 => \N__21042\,
            in2 => \_gnd_net_\,
            in3 => \N__20351\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__48777\,
            ce => \N__29217\,
            sr => \N__48202\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29101\,
            in1 => \N__21018\,
            in2 => \_gnd_net_\,
            in3 => \N__20348\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__48777\,
            ce => \N__29217\,
            sr => \N__48202\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29105\,
            in1 => \N__20994\,
            in2 => \_gnd_net_\,
            in3 => \N__20345\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__48777\,
            ce => \N__29217\,
            sr => \N__48202\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29102\,
            in1 => \N__20973\,
            in2 => \_gnd_net_\,
            in3 => \N__20342\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__48777\,
            ce => \N__29217\,
            sr => \N__48202\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29106\,
            in1 => \N__20949\,
            in2 => \_gnd_net_\,
            in3 => \N__20393\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__48777\,
            ce => \N__29217\,
            sr => \N__48202\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29103\,
            in1 => \N__20914\,
            in2 => \_gnd_net_\,
            in3 => \N__20390\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__48777\,
            ce => \N__29217\,
            sr => \N__48202\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29107\,
            in1 => \N__20889\,
            in2 => \_gnd_net_\,
            in3 => \N__20387\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__48777\,
            ce => \N__29217\,
            sr => \N__48202\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29058\,
            in1 => \N__20859\,
            in2 => \_gnd_net_\,
            in3 => \N__20384\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__48767\,
            ce => \N__29210\,
            sr => \N__48209\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29062\,
            in1 => \N__21165\,
            in2 => \_gnd_net_\,
            in3 => \N__20381\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__48767\,
            ce => \N__29210\,
            sr => \N__48209\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29059\,
            in1 => \N__21126\,
            in2 => \_gnd_net_\,
            in3 => \N__20378\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__48767\,
            ce => \N__29210\,
            sr => \N__48209\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29063\,
            in1 => \N__21084\,
            in2 => \_gnd_net_\,
            in3 => \N__20375\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__48767\,
            ce => \N__29210\,
            sr => \N__48209\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__29060\,
            in1 => \N__21145\,
            in2 => \_gnd_net_\,
            in3 => \N__20372\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__48767\,
            ce => \N__29210\,
            sr => \N__48209\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21103\,
            in1 => \N__29061\,
            in2 => \_gnd_net_\,
            in3 => \N__20369\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48767\,
            ce => \N__29210\,
            sr => \N__48209\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21956\,
            in2 => \N__20618\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__48759\,
            ce => \N__29882\,
            sr => \N__48217\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20587\,
            in2 => \N__21935\,
            in3 => \N__20621\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__48759\,
            ce => \N__29882\,
            sr => \N__48217\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20617\,
            in2 => \N__20563\,
            in3 => \N__20591\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__48759\,
            ce => \N__29882\,
            sr => \N__48217\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20588\,
            in2 => \N__20536\,
            in3 => \N__20567\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__48759\,
            ce => \N__29882\,
            sr => \N__48217\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20509\,
            in2 => \N__20564\,
            in3 => \N__20540\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__48759\,
            ce => \N__29882\,
            sr => \N__48217\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20485\,
            in2 => \N__20537\,
            in3 => \N__20513\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__48759\,
            ce => \N__29882\,
            sr => \N__48217\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20510\,
            in2 => \N__20461\,
            in3 => \N__20489\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__48759\,
            ce => \N__29882\,
            sr => \N__48217\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20486\,
            in2 => \N__20836\,
            in3 => \N__20465\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__48759\,
            ce => \N__29882\,
            sr => \N__48217\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20806\,
            in2 => \N__20462\,
            in3 => \N__20396\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__48746\,
            ce => \N__29887\,
            sr => \N__48221\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20782\,
            in2 => \N__20840\,
            in3 => \N__20810\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__48746\,
            ce => \N__29887\,
            sr => \N__48221\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20807\,
            in2 => \N__20761\,
            in3 => \N__20786\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__48746\,
            ce => \N__29887\,
            sr => \N__48221\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20783\,
            in2 => \N__20734\,
            in3 => \N__20765\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__48746\,
            ce => \N__29887\,
            sr => \N__48221\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20704\,
            in2 => \N__20762\,
            in3 => \N__20738\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__48746\,
            ce => \N__29887\,
            sr => \N__48221\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20674\,
            in2 => \N__20735\,
            in3 => \N__20711\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__48746\,
            ce => \N__29887\,
            sr => \N__48221\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20644\,
            in2 => \N__20708\,
            in3 => \N__20681\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__48746\,
            ce => \N__29887\,
            sr => \N__48221\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21049\,
            in2 => \N__20678\,
            in3 => \N__20651\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__48746\,
            ce => \N__29887\,
            sr => \N__48221\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21019\,
            in2 => \N__20648\,
            in3 => \N__20624\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__48734\,
            ce => \N__29886\,
            sr => \N__48228\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20995\,
            in2 => \N__21053\,
            in3 => \N__21026\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__48734\,
            ce => \N__29886\,
            sr => \N__48228\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20974\,
            in2 => \N__21023\,
            in3 => \N__20999\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__48734\,
            ce => \N__29886\,
            sr => \N__48228\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20996\,
            in2 => \N__20954\,
            in3 => \N__20978\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__48734\,
            ce => \N__29886\,
            sr => \N__48228\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20975\,
            in2 => \N__20926\,
            in3 => \N__20957\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__48734\,
            ce => \N__29886\,
            sr => \N__48228\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20953\,
            in2 => \N__20896\,
            in3 => \N__20930\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__48734\,
            ce => \N__29886\,
            sr => \N__48228\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20866\,
            in2 => \N__20927\,
            in3 => \N__20900\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__48734\,
            ce => \N__29886\,
            sr => \N__48228\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21172\,
            in2 => \N__20897\,
            in3 => \N__20873\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__48734\,
            ce => \N__29886\,
            sr => \N__48228\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21127\,
            in2 => \N__20870\,
            in3 => \N__20843\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__48724\,
            ce => \N__29875\,
            sr => \N__48233\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21085\,
            in2 => \N__21176\,
            in3 => \N__21149\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__48724\,
            ce => \N__29875\,
            sr => \N__48233\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21146\,
            in2 => \N__21131\,
            in3 => \N__21107\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__48724\,
            ce => \N__29875\,
            sr => \N__48233\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21104\,
            in2 => \N__21089\,
            in3 => \N__21065\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__48724\,
            ce => \N__29875\,
            sr => \N__48233\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21062\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48724\,
            ce => \N__29875\,
            sr => \N__48233\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__26375\,
            in1 => \N__28865\,
            in2 => \_gnd_net_\,
            in3 => \N__29309\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__26435\,
            in1 => \N__28967\,
            in2 => \_gnd_net_\,
            in3 => \N__29306\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__29310\,
            in1 => \N__26360\,
            in2 => \_gnd_net_\,
            in3 => \N__28838\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22510\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__29308\,
            in1 => \N__28898\,
            in2 => \_gnd_net_\,
            in3 => \N__26390\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29311\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__29307\,
            in1 => \N__28928\,
            in2 => \_gnd_net_\,
            in3 => \N__26405\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33648\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21260\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48704\,
            ce => \N__33742\,
            sr => \N__48243\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33772\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48704\,
            ce => \N__33742\,
            sr => \N__48243\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__37879\,
            in1 => \N__21185\,
            in2 => \_gnd_net_\,
            in3 => \N__22636\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37880\,
            in2 => \N__21179\,
            in3 => \N__29446\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__27126\,
            in1 => \N__33611\,
            in2 => \_gnd_net_\,
            in3 => \N__27086\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__33615\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33272\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111000101"
        )
    port map (
            in0 => \N__24148\,
            in1 => \N__24787\,
            in2 => \N__33617\,
            in3 => \N__33273\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__26922\,
            in1 => \N__24147\,
            in2 => \_gnd_net_\,
            in3 => \N__24786\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33771\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48696\,
            ce => \N__33741\,
            sr => \N__48250\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26549\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24378\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__26550\,
            in1 => \N__26921\,
            in2 => \_gnd_net_\,
            in3 => \N__26528\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29675\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34219\,
            in1 => \N__21256\,
            in2 => \_gnd_net_\,
            in3 => \N__21239\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__48685\,
            ce => \N__32582\,
            sr => \N__48263\
        );

    \current_shift_inst.timer_s1.counter_1_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34223\,
            in1 => \N__23956\,
            in2 => \_gnd_net_\,
            in3 => \N__21236\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__48685\,
            ce => \N__32582\,
            sr => \N__48263\
        );

    \current_shift_inst.timer_s1.counter_2_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34220\,
            in1 => \N__21231\,
            in2 => \_gnd_net_\,
            in3 => \N__21212\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__48685\,
            ce => \N__32582\,
            sr => \N__48263\
        );

    \current_shift_inst.timer_s1.counter_3_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34224\,
            in1 => \N__21207\,
            in2 => \_gnd_net_\,
            in3 => \N__21188\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__48685\,
            ce => \N__32582\,
            sr => \N__48263\
        );

    \current_shift_inst.timer_s1.counter_4_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34221\,
            in1 => \N__21451\,
            in2 => \_gnd_net_\,
            in3 => \N__21431\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__48685\,
            ce => \N__32582\,
            sr => \N__48263\
        );

    \current_shift_inst.timer_s1.counter_5_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34225\,
            in1 => \N__21427\,
            in2 => \_gnd_net_\,
            in3 => \N__21407\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__48685\,
            ce => \N__32582\,
            sr => \N__48263\
        );

    \current_shift_inst.timer_s1.counter_6_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34222\,
            in1 => \N__21403\,
            in2 => \_gnd_net_\,
            in3 => \N__21383\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__48685\,
            ce => \N__32582\,
            sr => \N__48263\
        );

    \current_shift_inst.timer_s1.counter_7_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34226\,
            in1 => \N__21379\,
            in2 => \_gnd_net_\,
            in3 => \N__21359\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__48685\,
            ce => \N__32582\,
            sr => \N__48263\
        );

    \current_shift_inst.timer_s1.counter_8_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34157\,
            in1 => \N__21355\,
            in2 => \_gnd_net_\,
            in3 => \N__21335\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__48680\,
            ce => \N__32584\,
            sr => \N__48266\
        );

    \current_shift_inst.timer_s1.counter_9_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34161\,
            in1 => \N__21331\,
            in2 => \_gnd_net_\,
            in3 => \N__21311\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__48680\,
            ce => \N__32584\,
            sr => \N__48266\
        );

    \current_shift_inst.timer_s1.counter_10_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34154\,
            in1 => \N__21307\,
            in2 => \_gnd_net_\,
            in3 => \N__21287\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__48680\,
            ce => \N__32584\,
            sr => \N__48266\
        );

    \current_shift_inst.timer_s1.counter_11_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34158\,
            in1 => \N__21283\,
            in2 => \_gnd_net_\,
            in3 => \N__21263\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__48680\,
            ce => \N__32584\,
            sr => \N__48266\
        );

    \current_shift_inst.timer_s1.counter_12_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34155\,
            in1 => \N__21664\,
            in2 => \_gnd_net_\,
            in3 => \N__21644\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__48680\,
            ce => \N__32584\,
            sr => \N__48266\
        );

    \current_shift_inst.timer_s1.counter_13_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34159\,
            in1 => \N__21640\,
            in2 => \_gnd_net_\,
            in3 => \N__21620\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__48680\,
            ce => \N__32584\,
            sr => \N__48266\
        );

    \current_shift_inst.timer_s1.counter_14_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34156\,
            in1 => \N__21616\,
            in2 => \_gnd_net_\,
            in3 => \N__21596\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__48680\,
            ce => \N__32584\,
            sr => \N__48266\
        );

    \current_shift_inst.timer_s1.counter_15_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34160\,
            in1 => \N__21592\,
            in2 => \_gnd_net_\,
            in3 => \N__21572\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__48680\,
            ce => \N__32584\,
            sr => \N__48266\
        );

    \current_shift_inst.timer_s1.counter_16_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34191\,
            in1 => \N__21568\,
            in2 => \_gnd_net_\,
            in3 => \N__21548\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_21_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__48676\,
            ce => \N__32583\,
            sr => \N__48271\
        );

    \current_shift_inst.timer_s1.counter_17_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34121\,
            in1 => \N__21544\,
            in2 => \_gnd_net_\,
            in3 => \N__21524\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__48676\,
            ce => \N__32583\,
            sr => \N__48271\
        );

    \current_shift_inst.timer_s1.counter_18_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34192\,
            in1 => \N__21520\,
            in2 => \_gnd_net_\,
            in3 => \N__21500\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__48676\,
            ce => \N__32583\,
            sr => \N__48271\
        );

    \current_shift_inst.timer_s1.counter_19_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34122\,
            in1 => \N__21496\,
            in2 => \_gnd_net_\,
            in3 => \N__21476\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__48676\,
            ce => \N__32583\,
            sr => \N__48271\
        );

    \current_shift_inst.timer_s1.counter_20_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34193\,
            in1 => \N__21472\,
            in2 => \_gnd_net_\,
            in3 => \N__21851\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__48676\,
            ce => \N__32583\,
            sr => \N__48271\
        );

    \current_shift_inst.timer_s1.counter_21_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34123\,
            in1 => \N__21847\,
            in2 => \_gnd_net_\,
            in3 => \N__21827\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__48676\,
            ce => \N__32583\,
            sr => \N__48271\
        );

    \current_shift_inst.timer_s1.counter_22_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34194\,
            in1 => \N__21823\,
            in2 => \_gnd_net_\,
            in3 => \N__21803\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__48676\,
            ce => \N__32583\,
            sr => \N__48271\
        );

    \current_shift_inst.timer_s1.counter_23_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34124\,
            in1 => \N__21799\,
            in2 => \_gnd_net_\,
            in3 => \N__21779\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__48676\,
            ce => \N__32583\,
            sr => \N__48271\
        );

    \current_shift_inst.timer_s1.counter_24_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34204\,
            in1 => \N__21775\,
            in2 => \_gnd_net_\,
            in3 => \N__21755\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_22_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__48670\,
            ce => \N__32588\,
            sr => \N__48275\
        );

    \current_shift_inst.timer_s1.counter_25_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34208\,
            in1 => \N__21751\,
            in2 => \_gnd_net_\,
            in3 => \N__21731\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__48670\,
            ce => \N__32588\,
            sr => \N__48275\
        );

    \current_shift_inst.timer_s1.counter_26_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34205\,
            in1 => \N__21727\,
            in2 => \_gnd_net_\,
            in3 => \N__21707\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__48670\,
            ce => \N__32588\,
            sr => \N__48275\
        );

    \current_shift_inst.timer_s1.counter_27_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34209\,
            in1 => \N__21703\,
            in2 => \_gnd_net_\,
            in3 => \N__21683\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__48670\,
            ce => \N__32588\,
            sr => \N__48275\
        );

    \current_shift_inst.timer_s1.counter_28_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34206\,
            in1 => \N__21680\,
            in2 => \_gnd_net_\,
            in3 => \N__21668\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__48670\,
            ce => \N__32588\,
            sr => \N__48275\
        );

    \current_shift_inst.timer_s1.counter_29_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21905\,
            in1 => \N__34207\,
            in2 => \_gnd_net_\,
            in3 => \N__21908\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48670\,
            ce => \N__32588\,
            sr => \N__48275\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30286\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30555\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S2_LC_8_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31732\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48648\,
            ce => 'H',
            sr => \N__48286\
        );

    \GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48812\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clock_output_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21878\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21867\,
            in1 => \N__23293\,
            in2 => \_gnd_net_\,
            in3 => \N__41891\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48807\,
            ce => \N__28514\,
            sr => \N__48141\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21868\,
            in1 => \N__23294\,
            in2 => \_gnd_net_\,
            in3 => \N__41895\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48806\,
            ce => \N__36608\,
            sr => \N__48149\
        );

    \phase_controller_inst2.stoper_hc.target_time_20_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31374\,
            in1 => \N__31357\,
            in2 => \_gnd_net_\,
            in3 => \N__41879\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48801\,
            ce => \N__28513\,
            sr => \N__48157\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41850\,
            in1 => \N__25058\,
            in2 => \_gnd_net_\,
            in3 => \N__25102\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48797\,
            ce => \N__28512\,
            sr => \N__48166\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41849\,
            in1 => \N__23178\,
            in2 => \_gnd_net_\,
            in3 => \N__23134\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48797\,
            ce => \N__28512\,
            sr => \N__48166\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31584\,
            in1 => \N__31502\,
            in2 => \N__41943\,
            in3 => \N__38249\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23579\,
            in1 => \N__28577\,
            in2 => \N__23439\,
            in3 => \N__28640\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21968\,
            in1 => \N__23981\,
            in2 => \N__21962\,
            in3 => \N__23249\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23532\,
            in1 => \N__41668\,
            in2 => \_gnd_net_\,
            in3 => \N__23513\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48787\,
            ce => \N__36601\,
            sr => \N__48174\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22997\,
            in1 => \N__23039\,
            in2 => \N__23098\,
            in3 => \N__23852\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31878\,
            in2 => \N__21959\,
            in3 => \N__28166\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21955\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48778\,
            ce => \N__29888\,
            sr => \N__48183\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21928\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48778\,
            ce => \N__29888\,
            sr => \N__48183\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23040\,
            in1 => \N__23066\,
            in2 => \_gnd_net_\,
            in3 => \N__41743\,
            lcout => \elapsed_time_ns_1_RNIE03T9_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22998\,
            in1 => \N__41653\,
            in2 => \_gnd_net_\,
            in3 => \N__23021\,
            lcout => \elapsed_time_ns_1_RNIF13T9_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23093\,
            in1 => \N__23117\,
            in2 => \_gnd_net_\,
            in3 => \N__41742\,
            lcout => \elapsed_time_ns_1_RNIG23T9_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__22022\,
            in1 => \N__25964\,
            in2 => \N__25997\,
            in3 => \N__22004\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23041\,
            in1 => \N__23064\,
            in2 => \_gnd_net_\,
            in3 => \N__41666\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48768\,
            ce => \N__28509\,
            sr => \N__48193\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41665\,
            in1 => \N__23019\,
            in2 => \_gnd_net_\,
            in3 => \N__22999\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48768\,
            ce => \N__28509\,
            sr => \N__48193\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23115\,
            in1 => \N__23097\,
            in2 => \_gnd_net_\,
            in3 => \N__41667\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48768\,
            ce => \N__28509\,
            sr => \N__48193\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__25936\,
            in1 => \N__23542\,
            in2 => \N__25913\,
            in3 => \N__21983\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011111011"
        )
    port map (
            in0 => \N__21982\,
            in1 => \N__25937\,
            in2 => \N__23546\,
            in3 => \N__25912\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41787\,
            in1 => \N__24909\,
            in2 => \_gnd_net_\,
            in3 => \N__24944\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48760\,
            ce => \N__28505\,
            sr => \N__48203\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23234\,
            in1 => \N__41786\,
            in2 => \_gnd_net_\,
            in3 => \N__23212\,
            lcout => \elapsed_time_ns_1_RNIK63T9_0_8\,
            ltout => \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__41788\,
            in1 => \_gnd_net_\,
            in2 => \N__22124\,
            in3 => \N__23235\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48760\,
            ce => \N__28505\,
            sr => \N__48203\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23831\,
            in2 => \N__22121\,
            in3 => \N__25416\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22112\,
            in2 => \N__22103\,
            in3 => \N__25682\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22082\,
            in2 => \N__22094\,
            in3 => \N__25655\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22076\,
            in2 => \N__22067\,
            in3 => \N__25637\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22058\,
            in2 => \N__22046\,
            in3 => \N__25616\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25598\,
            in1 => \N__22037\,
            in2 => \N__22031\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22262\,
            in2 => \N__22253\,
            in3 => \N__25580\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22244\,
            in2 => \N__22235\,
            in3 => \N__25559\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22214\,
            in2 => \N__22226\,
            in3 => \N__25541\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22202\,
            in2 => \N__22193\,
            in3 => \N__25826\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25808\,
            in1 => \N__22184\,
            in2 => \N__22175\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22163\,
            in2 => \N__28679\,
            in3 => \N__25790\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23474\,
            in2 => \N__22157\,
            in3 => \N__25772\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25754\,
            in1 => \N__22145\,
            in2 => \N__22133\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25736\,
            in1 => \N__22361\,
            in2 => \N__22349\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24068\,
            in2 => \N__24164\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22340\,
            in2 => \N__22331\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22313\,
            in2 => \N__22304\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22289\,
            in2 => \N__22277\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27953\,
            in2 => \N__28004\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24197\,
            in2 => \N__28382\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28103\,
            in2 => \N__28019\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23765\,
            in2 => \N__23810\,
            in3 => \N__22493\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22490\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24293\,
            in2 => \N__24284\,
            in3 => \N__24282\,
            lcout => \current_shift_inst.control_input_18\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22499\,
            in2 => \_gnd_net_\,
            in3 => \N__22463\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22460\,
            in2 => \_gnd_net_\,
            in3 => \N__22442\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22649\,
            in2 => \_gnd_net_\,
            in3 => \N__22427\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22424\,
            in2 => \_gnd_net_\,
            in3 => \N__22406\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22403\,
            in2 => \_gnd_net_\,
            in3 => \N__22385\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22382\,
            in2 => \_gnd_net_\,
            in3 => \N__22364\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22622\,
            in2 => \_gnd_net_\,
            in3 => \N__22604\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29366\,
            in2 => \_gnd_net_\,
            in3 => \N__22589\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29342\,
            in2 => \_gnd_net_\,
            in3 => \N__22574\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29231\,
            in2 => \_gnd_net_\,
            in3 => \N__22559\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29390\,
            in2 => \_gnd_net_\,
            in3 => \N__22544\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22541\,
            in2 => \_gnd_net_\,
            in3 => \N__22523\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29305\,
            in2 => \_gnd_net_\,
            in3 => \N__22520\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__29303\,
            in1 => \N__26450\,
            in2 => \_gnd_net_\,
            in3 => \N__28979\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__26420\,
            in1 => \N__28955\,
            in2 => \_gnd_net_\,
            in3 => \N__29304\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31958\,
            in2 => \N__22643\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37866\,
            in2 => \N__24215\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24320\,
            in2 => \N__37906\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37870\,
            in2 => \N__24587\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24326\,
            in2 => \N__37907\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37874\,
            in2 => \N__24356\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24170\,
            in2 => \N__37908\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37878\,
            in2 => \N__24347\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22667\,
            in2 => \N__37905\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37865\,
            in2 => \N__24308\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22754\,
            in2 => \N__37902\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37853\,
            in2 => \N__24335\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22739\,
            in2 => \N__37903\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37857\,
            in2 => \N__22661\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24314\,
            in2 => \N__37904\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37861\,
            in2 => \N__24404\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37834\,
            in2 => \N__22775\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26855\,
            in2 => \N__37898\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37838\,
            in2 => \N__22817\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26660\,
            in2 => \N__37899\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37842\,
            in2 => \N__26687\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22673\,
            in2 => \N__37900\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37846\,
            in2 => \N__26702\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22730\,
            in2 => \N__37901\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37717\,
            in2 => \N__22688\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22694\,
            in2 => \N__37831\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37721\,
            in2 => \N__22721\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22679\,
            in2 => \N__37832\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37725\,
            in2 => \N__22709\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22745\,
            in2 => \N__37833\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37729\,
            in2 => \N__22763\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33589\,
            in2 => \_gnd_net_\,
            in3 => \N__22697\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33607\,
            in1 => \N__27189\,
            in2 => \_gnd_net_\,
            in3 => \N__27148\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__26984\,
            in1 => \N__27051\,
            in2 => \_gnd_net_\,
            in3 => \N__27009\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__33608\,
            in1 => \N__33849\,
            in2 => \N__33811\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__29532\,
            in1 => \N__26983\,
            in2 => \_gnd_net_\,
            in3 => \N__29478\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__33610\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31999\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__30405\,
            in1 => \N__26981\,
            in2 => \_gnd_net_\,
            in3 => \N__30369\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33609\,
            in1 => \N__30573\,
            in2 => \_gnd_net_\,
            in3 => \N__30525\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32328\,
            in1 => \N__26982\,
            in2 => \_gnd_net_\,
            in3 => \N__32283\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__26977\,
            in1 => \N__30069\,
            in2 => \_gnd_net_\,
            in3 => \N__30090\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32139\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33547\,
            in1 => \N__26643\,
            in2 => \_gnd_net_\,
            in3 => \N__26604\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27044\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30396\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30159\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__26976\,
            in1 => \N__29964\,
            in2 => \_gnd_net_\,
            in3 => \N__30007\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32459\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24135\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27180\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30056\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27119\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30236\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22805\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48661\,
            ce => 'H',
            sr => \N__48276\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22928\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48661\,
            ce => 'H',
            sr => \N__48276\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22901\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48661\,
            ce => 'H',
            sr => \N__48276\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22871\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48658\,
            ce => 'H',
            sr => \N__48279\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22847\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48658\,
            ce => 'H',
            sr => \N__48279\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31378\,
            in1 => \N__31356\,
            in2 => \_gnd_net_\,
            in3 => \N__41779\,
            lcout => \elapsed_time_ns_1_RNIU0DN9_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__23335\,
            in1 => \N__27709\,
            in2 => \N__27743\,
            in3 => \N__23197\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41783\,
            in1 => \N__23179\,
            in2 => \_gnd_net_\,
            in3 => \N__23135\,
            lcout => \elapsed_time_ns_1_RNIH33T9_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_30_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41771\,
            in1 => \N__23463\,
            in2 => \_gnd_net_\,
            in3 => \N__23440\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48780\,
            ce => \N__36597\,
            sr => \N__48150\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25101\,
            in1 => \N__25053\,
            in2 => \_gnd_net_\,
            in3 => \N__41775\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48780\,
            ce => \N__36597\,
            sr => \N__48150\
        );

    \phase_controller_inst1.stoper_hc.target_time_31_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41772\,
            in1 => \N__23939\,
            in2 => \_gnd_net_\,
            in3 => \N__23380\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48780\,
            ce => \N__36597\,
            sr => \N__48150\
        );

    \phase_controller_inst1.stoper_hc.target_time_24_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38200\,
            in1 => \N__38260\,
            in2 => \_gnd_net_\,
            in3 => \N__41774\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48780\,
            ce => \N__36597\,
            sr => \N__48150\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41773\,
            in1 => \N__23180\,
            in2 => \_gnd_net_\,
            in3 => \N__23133\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48780\,
            ce => \N__36597\,
            sr => \N__48150\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23116\,
            in1 => \N__23099\,
            in2 => \_gnd_net_\,
            in3 => \N__41659\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48769\,
            ce => \N__36605\,
            sr => \N__48158\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__41655\,
            in1 => \N__23065\,
            in2 => \N__23048\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48769\,
            ce => \N__36605\,
            sr => \N__48158\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41656\,
            in1 => \N__23020\,
            in2 => \_gnd_net_\,
            in3 => \N__23003\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48769\,
            ce => \N__36605\,
            sr => \N__48158\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22976\,
            in1 => \N__24057\,
            in2 => \_gnd_net_\,
            in3 => \N__41658\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48769\,
            ce => \N__36605\,
            sr => \N__48158\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41654\,
            in1 => \N__23891\,
            in2 => \_gnd_net_\,
            in3 => \N__23856\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48769\,
            ce => \N__36605\,
            sr => \N__48158\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22952\,
            in1 => \N__24022\,
            in2 => \_gnd_net_\,
            in3 => \N__41657\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48769\,
            ce => \N__36605\,
            sr => \N__48158\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__27776\,
            in1 => \N__23350\,
            in2 => \N__27554\,
            in3 => \N__23360\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__23359\,
            in1 => \N__27775\,
            in2 => \N__23351\,
            in3 => \N__27553\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__27739\,
            in1 => \N__23339\,
            in2 => \N__23201\,
            in3 => \N__27710\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__23937\,
            in1 => \N__23324\,
            in2 => \N__23318\,
            in3 => \N__23303\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27297\,
            in1 => \_gnd_net_\,
            in2 => \N__23297\,
            in3 => \N__27327\,
            lcout => \elapsed_time_ns_1_RNI35CN9_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41652\,
            in1 => \N__23465\,
            in2 => \_gnd_net_\,
            in3 => \N__23432\,
            lcout => \elapsed_time_ns_1_RNIV2EN9_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23511\,
            in1 => \N__23533\,
            in2 => \_gnd_net_\,
            in3 => \N__41651\,
            lcout => \elapsed_time_ns_1_RNI02CN9_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23282\,
            in1 => \N__23510\,
            in2 => \N__30769\,
            in3 => \N__27296\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23243\,
            in1 => \N__41663\,
            in2 => \_gnd_net_\,
            in3 => \N__23213\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48748\,
            ce => \N__36606\,
            sr => \N__48175\
        );

    \phase_controller_inst1.stoper_hc.target_time_25_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41660\,
            in1 => \N__28662\,
            in2 => \_gnd_net_\,
            in3 => \N__28645\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48748\,
            ce => \N__36606\,
            sr => \N__48175\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23741\,
            in1 => \N__23714\,
            in2 => \_gnd_net_\,
            in3 => \N__41664\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48748\,
            ce => \N__36606\,
            sr => \N__48175\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41662\,
            in1 => \N__23677\,
            in2 => \_gnd_net_\,
            in3 => \N__23651\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48748\,
            ce => \N__36606\,
            sr => \N__48175\
        );

    \phase_controller_inst1.stoper_hc.target_time_29_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41661\,
            in1 => \N__23618\,
            in2 => \_gnd_net_\,
            in3 => \N__23591\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48748\,
            ce => \N__36606\,
            sr => \N__48175\
        );

    \phase_controller_inst2.stoper_hc.target_time_21_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41419\,
            in1 => \N__41942\,
            in2 => \_gnd_net_\,
            in3 => \N__41794\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48736\,
            ce => \N__28506\,
            sr => \N__48184\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27328\,
            in1 => \N__27301\,
            in2 => \_gnd_net_\,
            in3 => \N__41793\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48736\,
            ce => \N__28506\,
            sr => \N__48184\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41789\,
            in1 => \N__25127\,
            in2 => \_gnd_net_\,
            in3 => \N__25165\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48736\,
            ce => \N__28506\,
            sr => \N__48184\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23534\,
            in1 => \N__41792\,
            in2 => \_gnd_net_\,
            in3 => \N__23512\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48736\,
            ce => \N__28506\,
            sr => \N__48184\
        );

    \phase_controller_inst2.stoper_hc.target_time_30_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41791\,
            in1 => \N__23464\,
            in2 => \_gnd_net_\,
            in3 => \N__23441\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48736\,
            ce => \N__28506\,
            sr => \N__48184\
        );

    \phase_controller_inst2.stoper_hc.target_time_31_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41795\,
            in1 => \N__23384\,
            in2 => \_gnd_net_\,
            in3 => \N__23933\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48736\,
            ce => \N__28506\,
            sr => \N__48184\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41790\,
            in1 => \N__23884\,
            in2 => \_gnd_net_\,
            in3 => \N__23863\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48736\,
            ce => \N__28506\,
            sr => \N__48184\
        );

    \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__23776\,
            in1 => \N__26232\,
            in2 => \N__26045\,
            in3 => \N__23788\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.stoper_hc.un4_running_df30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101011101"
        )
    port map (
            in0 => \N__28210\,
            in1 => \N__23800\,
            in2 => \N__23825\,
            in3 => \N__23822\,
            lcout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23813\,
            in3 => \N__28256\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001110"
        )
    port map (
            in0 => \N__23787\,
            in1 => \N__26040\,
            in2 => \N__26236\,
            in3 => \N__23775\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28257\,
            in2 => \_gnd_net_\,
            in3 => \N__23752\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110011101111"
        )
    port map (
            in0 => \N__23789\,
            in1 => \N__26044\,
            in2 => \N__26237\,
            in3 => \N__23777\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__26203\,
            in1 => \N__25420\,
            in2 => \N__23756\,
            in3 => \N__28261\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48726\,
            ce => 'H',
            sr => \N__48194\
        );

    \phase_controller_inst2.stoper_hc.running_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101111101010000"
        )
    port map (
            in0 => \N__28211\,
            in1 => \N__28237\,
            in2 => \N__28262\,
            in3 => \N__28297\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48726\,
            ce => 'H',
            sr => \N__48194\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33606\,
            in1 => \N__30259\,
            in2 => \N__33278\,
            in3 => \N__30212\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010110010"
        )
    port map (
            in0 => \N__24098\,
            in1 => \N__25699\,
            in2 => \N__24085\,
            in3 => \N__25717\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33605\,
            in1 => \N__24152\,
            in2 => \N__33277\,
            in3 => \N__24788\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24113\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48716\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010111011"
        )
    port map (
            in0 => \N__24097\,
            in1 => \N__25698\,
            in2 => \N__24086\,
            in3 => \N__25716\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24042\,
            in1 => \N__25154\,
            in2 => \N__31346\,
            in3 => \N__24005\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__33603\,
            in1 => \N__24568\,
            in2 => \N__28331\,
            in3 => \N__24187\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23966\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48706\,
            ce => \N__33743\,
            sr => \N__48210\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001011"
        )
    port map (
            in0 => \N__24569\,
            in1 => \N__33604\,
            in2 => \N__24191\,
            in3 => \N__28330\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__26985\,
            in1 => \N__24567\,
            in2 => \_gnd_net_\,
            in3 => \N__24186\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33551\,
            in1 => \N__24262\,
            in2 => \N__33280\,
            in3 => \N__24697\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__32426\,
            in1 => \N__33550\,
            in2 => \N__32384\,
            in3 => \N__33228\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33553\,
            in1 => \N__24440\,
            in2 => \N__33279\,
            in3 => \N__24620\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__24394\,
            in1 => \N__33229\,
            in2 => \N__24500\,
            in3 => \N__33549\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__28469\,
            in1 => \N__28449\,
            in2 => \N__28426\,
            in3 => \N__28400\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24185\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__29582\,
            in1 => \N__33230\,
            in2 => \N__29636\,
            in3 => \N__33552\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__26964\,
            in1 => \N__29628\,
            in2 => \_gnd_net_\,
            in3 => \N__29574\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__26965\,
            in1 => \N__24249\,
            in2 => \_gnd_net_\,
            in3 => \N__24696\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__26312\,
            in1 => \N__28796\,
            in2 => \_gnd_net_\,
            in3 => \N__29301\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => \current_shift_inst.control_input_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24287\,
            in3 => \N__24283\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48689\,
            ce => 'H',
            sr => \N__48222\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29302\,
            lcout => \current_shift_inst.N_1288_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__33555\,
            in1 => \N__24395\,
            in2 => \N__24499\,
            in3 => \N__33209\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__24619\,
            in1 => \N__33560\,
            in2 => \N__33276\,
            in3 => \N__24436\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__33556\,
            in1 => \N__33210\,
            in2 => \N__29693\,
            in3 => \N__29719\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__30500\,
            in1 => \N__33558\,
            in2 => \N__33274\,
            in3 => \N__30452\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__33554\,
            in1 => \N__33208\,
            in2 => \N__29816\,
            in3 => \N__29768\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__33211\,
            in1 => \N__24698\,
            in2 => \N__24263\,
            in3 => \N__33557\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__24435\,
            in1 => \N__26993\,
            in2 => \_gnd_net_\,
            in3 => \N__24618\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32338\,
            in1 => \N__33559\,
            in2 => \N__33275\,
            in3 => \N__32290\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__24387\,
            in1 => \N__26939\,
            in2 => \_gnd_net_\,
            in3 => \N__24483\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33234\,
            in1 => \N__33561\,
            in2 => \N__26566\,
            in3 => \N__26526\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__29691\,
            in1 => \N__26940\,
            in2 => \_gnd_net_\,
            in3 => \N__29709\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__26941\,
            in1 => \N__30495\,
            in2 => \_gnd_net_\,
            in3 => \N__30450\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32418\,
            in1 => \N__26938\,
            in2 => \_gnd_net_\,
            in3 => \N__32362\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__26936\,
            in1 => \N__32667\,
            in2 => \_gnd_net_\,
            in3 => \N__32625\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__32238\,
            in1 => \N__26942\,
            in2 => \_gnd_net_\,
            in3 => \N__32187\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__26937\,
            in1 => \N__29802\,
            in2 => \_gnd_net_\,
            in3 => \N__29760\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24578\,
            in2 => \N__33712\,
            in3 => \N__33708\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24554\,
            in2 => \_gnd_net_\,
            in3 => \N__24542\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24539\,
            in2 => \_gnd_net_\,
            in3 => \N__24527\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24524\,
            in2 => \_gnd_net_\,
            in3 => \N__24512\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24509\,
            in2 => \_gnd_net_\,
            in3 => \N__24470\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24467\,
            in2 => \_gnd_net_\,
            in3 => \N__24455\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24452\,
            in2 => \_gnd_net_\,
            in3 => \N__24443\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24719\,
            in2 => \_gnd_net_\,
            in3 => \N__24710\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24707\,
            in2 => \_gnd_net_\,
            in3 => \N__24674\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_10_19_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24671\,
            in2 => \_gnd_net_\,
            in3 => \N__24662\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26495\,
            in2 => \_gnd_net_\,
            in3 => \N__24659\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24656\,
            in2 => \_gnd_net_\,
            in3 => \N__24647\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24644\,
            in2 => \_gnd_net_\,
            in3 => \N__24635\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26489\,
            in2 => \_gnd_net_\,
            in3 => \N__24632\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24629\,
            in2 => \_gnd_net_\,
            in3 => \N__24602\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24599\,
            in2 => \_gnd_net_\,
            in3 => \N__24590\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24833\,
            in2 => \_gnd_net_\,
            in3 => \N__24827\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_10_20_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24845\,
            in2 => \_gnd_net_\,
            in3 => \N__24824\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24821\,
            in3 => \N__24809\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24806\,
            in2 => \_gnd_net_\,
            in3 => \N__24800\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24797\,
            in2 => \_gnd_net_\,
            in3 => \N__24758\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24755\,
            in2 => \_gnd_net_\,
            in3 => \N__24743\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24740\,
            in2 => \_gnd_net_\,
            in3 => \N__24731\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24728\,
            in2 => \_gnd_net_\,
            in3 => \N__24722\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24890\,
            in2 => \_gnd_net_\,
            in3 => \N__24884\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24959\,
            in2 => \_gnd_net_\,
            in3 => \N__24881\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24839\,
            in2 => \_gnd_net_\,
            in3 => \N__24878\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24875\,
            in2 => \_gnd_net_\,
            in3 => \N__24869\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24866\,
            in2 => \_gnd_net_\,
            in3 => \N__24854\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24851\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__33548\,
            in1 => \N__33292\,
            in2 => \N__24848\,
            in3 => \N__31982\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30005\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33848\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26642\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_27_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28178\,
            in1 => \N__28126\,
            in2 => \_gnd_net_\,
            in3 => \N__41897\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48788\,
            ce => \N__36596\,
            sr => \N__48131\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25123\,
            in1 => \N__25172\,
            in2 => \_gnd_net_\,
            in3 => \N__41896\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48788\,
            ce => \N__36596\,
            sr => \N__48131\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101100100010"
        )
    port map (
            in0 => \N__24952\,
            in1 => \N__27931\,
            in2 => \N__27677\,
            in3 => \N__27341\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__27340\,
            in1 => \N__27676\,
            in2 => \N__27932\,
            in3 => \N__24953\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41781\,
            in1 => \N__28534\,
            in2 => \_gnd_net_\,
            in3 => \N__28592\,
            lcout => \elapsed_time_ns_1_RNI47DN9_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24922\,
            in1 => \N__41780\,
            in2 => \_gnd_net_\,
            in3 => \N__24937\,
            lcout => \elapsed_time_ns_1_RNII43T9_0_6\,
            ltout => \elapsed_time_ns_1_RNII43T9_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__41782\,
            in1 => \_gnd_net_\,
            in2 => \N__24926\,
            in3 => \N__24923\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48781\,
            ce => \N__36607\,
            sr => \N__48136\
        );

    \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__27897\,
            in1 => \N__25035\,
            in2 => \N__27871\,
            in3 => \N__25020\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41769\,
            in1 => \N__28174\,
            in2 => \_gnd_net_\,
            in3 => \N__28125\,
            lcout => \elapsed_time_ns_1_RNI58DN9_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__25037\,
            in1 => \N__27870\,
            in2 => \N__25025\,
            in3 => \N__27899\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25122\,
            in1 => \N__25164\,
            in2 => \_gnd_net_\,
            in3 => \N__41768\,
            lcout => \elapsed_time_ns_1_RNI46CN9_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__41770\,
            in1 => \N__25057\,
            in2 => \N__25103\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIJ53T9_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__27898\,
            in1 => \N__25036\,
            in2 => \N__27872\,
            in3 => \N__25021\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101011101"
        )
    port map (
            in0 => \N__42355\,
            in1 => \N__25459\,
            in2 => \N__25010\,
            in3 => \N__25448\,
            lcout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27814\,
            in1 => \N__25007\,
            in2 => \N__25001\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27529\,
            in1 => \N__24992\,
            in2 => \N__24986\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27502\,
            in1 => \N__24974\,
            in2 => \N__24968\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25307\,
            in2 => \N__25301\,
            in3 => \N__27487\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25283\,
            in2 => \N__25292\,
            in3 => \N__27472\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25277\,
            in2 => \N__25268\,
            in3 => \N__27457\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25259\,
            in2 => \N__25250\,
            in3 => \N__27442\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25229\,
            in2 => \N__25241\,
            in3 => \N__27427\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25223\,
            in2 => \N__25217\,
            in3 => \N__27412\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25208\,
            in2 => \N__25202\,
            in3 => \N__27649\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25193\,
            in2 => \N__25184\,
            in3 => \N__27634\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27619\,
            in1 => \N__25400\,
            in2 => \N__25388\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25376\,
            in2 => \N__25364\,
            in3 => \N__27604\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27589\,
            in1 => \N__27353\,
            in2 => \N__25355\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27574\,
            in1 => \N__25331\,
            in2 => \N__25346\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30782\,
            in2 => \N__31142\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25322\,
            in2 => \N__25316\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31457\,
            in2 => \N__31409\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31625\,
            in2 => \N__31028\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25523\,
            in2 => \N__25511\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25502\,
            in2 => \N__25493\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25433\,
            in2 => \N__31247\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25478\,
            in2 => \N__25469\,
            in3 => \N__25439\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25436\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__31859\,
            in1 => \N__31303\,
            in2 => \N__31285\,
            in3 => \N__31264\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41784\,
            in1 => \N__28701\,
            in2 => \_gnd_net_\,
            in3 => \N__28745\,
            lcout => \elapsed_time_ns_1_RNIV0CN9_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28666\,
            in1 => \N__28641\,
            in2 => \_gnd_net_\,
            in3 => \N__41785\,
            lcout => \elapsed_time_ns_1_RNI36DN9_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25427\,
            in2 => \N__25421\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26153\,
            in1 => \N__25681\,
            in2 => \_gnd_net_\,
            in3 => \N__25667\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__48717\,
            ce => 'H',
            sr => \N__48185\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__26196\,
            in1 => \N__25654\,
            in2 => \N__25664\,
            in3 => \N__25640\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__48717\,
            ce => 'H',
            sr => \N__48185\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26154\,
            in1 => \N__25633\,
            in2 => \_gnd_net_\,
            in3 => \N__25619\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__48717\,
            ce => 'H',
            sr => \N__48185\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26197\,
            in1 => \N__25615\,
            in2 => \_gnd_net_\,
            in3 => \N__25601\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__48717\,
            ce => 'H',
            sr => \N__48185\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26155\,
            in1 => \N__25597\,
            in2 => \_gnd_net_\,
            in3 => \N__25583\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__48717\,
            ce => 'H',
            sr => \N__48185\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26198\,
            in1 => \N__25576\,
            in2 => \_gnd_net_\,
            in3 => \N__25562\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__48717\,
            ce => 'H',
            sr => \N__48185\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26156\,
            in1 => \N__25558\,
            in2 => \_gnd_net_\,
            in3 => \N__25544\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__48717\,
            ce => 'H',
            sr => \N__48185\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26202\,
            in1 => \N__25540\,
            in2 => \_gnd_net_\,
            in3 => \N__25526\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__48707\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26192\,
            in1 => \N__25825\,
            in2 => \_gnd_net_\,
            in3 => \N__25811\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__48707\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26199\,
            in1 => \N__25807\,
            in2 => \_gnd_net_\,
            in3 => \N__25793\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__48707\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26193\,
            in1 => \N__25789\,
            in2 => \_gnd_net_\,
            in3 => \N__25775\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__48707\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26200\,
            in1 => \N__25771\,
            in2 => \_gnd_net_\,
            in3 => \N__25757\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__48707\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26194\,
            in1 => \N__25753\,
            in2 => \_gnd_net_\,
            in3 => \N__25739\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__48707\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26201\,
            in1 => \N__25735\,
            in2 => \_gnd_net_\,
            in3 => \N__25721\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__48707\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26195\,
            in1 => \N__25718\,
            in2 => \_gnd_net_\,
            in3 => \N__25703\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__48707\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26145\,
            in1 => \N__25700\,
            in2 => \_gnd_net_\,
            in3 => \N__25685\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__48698\,
            ce => 'H',
            sr => \N__48204\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26157\,
            in1 => \N__25983\,
            in2 => \_gnd_net_\,
            in3 => \N__25967\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__48698\,
            ce => 'H',
            sr => \N__48204\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26146\,
            in1 => \N__25956\,
            in2 => \_gnd_net_\,
            in3 => \N__25940\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__48698\,
            ce => 'H',
            sr => \N__48204\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26158\,
            in1 => \N__25930\,
            in2 => \_gnd_net_\,
            in3 => \N__25916\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__48698\,
            ce => 'H',
            sr => \N__48204\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26147\,
            in1 => \N__25903\,
            in2 => \_gnd_net_\,
            in3 => \N__25889\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__48698\,
            ce => 'H',
            sr => \N__48204\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26159\,
            in1 => \N__25876\,
            in2 => \_gnd_net_\,
            in3 => \N__25862\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__48698\,
            ce => 'H',
            sr => \N__48204\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26148\,
            in1 => \N__25852\,
            in2 => \_gnd_net_\,
            in3 => \N__25838\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__48698\,
            ce => 'H',
            sr => \N__48204\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26160\,
            in1 => \N__27989\,
            in2 => \_gnd_net_\,
            in3 => \N__25835\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__48698\,
            ce => 'H',
            sr => \N__48204\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26149\,
            in1 => \N__27969\,
            in2 => \_gnd_net_\,
            in3 => \N__25832\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__48690\,
            ce => 'H',
            sr => \N__48211\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26142\,
            in1 => \N__28422\,
            in2 => \_gnd_net_\,
            in3 => \N__25829\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__48690\,
            ce => 'H',
            sr => \N__48211\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26150\,
            in1 => \N__28450\,
            in2 => \_gnd_net_\,
            in3 => \N__26246\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__48690\,
            ce => 'H',
            sr => \N__48211\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26143\,
            in1 => \N__28042\,
            in2 => \_gnd_net_\,
            in3 => \N__26243\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__48690\,
            ce => 'H',
            sr => \N__48211\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26151\,
            in1 => \N__28089\,
            in2 => \_gnd_net_\,
            in3 => \N__26240\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__48690\,
            ce => 'H',
            sr => \N__48211\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26144\,
            in1 => \N__26221\,
            in2 => \_gnd_net_\,
            in3 => \N__26207\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__48690\,
            ce => 'H',
            sr => \N__48211\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26152\,
            in1 => \N__26032\,
            in2 => \_gnd_net_\,
            in3 => \N__26048\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48690\,
            ce => 'H',
            sr => \N__48211\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28366\,
            in2 => \N__29447\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28326\,
            in2 => \N__26018\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32612\,
            in2 => \N__33121\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32916\,
            in2 => \N__26006\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26300\,
            in2 => \N__33122\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32920\,
            in2 => \N__26294\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26285\,
            in2 => \N__33123\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32924\,
            in2 => \N__26279\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26270\,
            in2 => \N__33124\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32928\,
            in2 => \N__26264\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26471\,
            in2 => \N__33125\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32932\,
            in2 => \N__26255\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26342\,
            in2 => \N__33126\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32936\,
            in2 => \N__32084\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32165\,
            in2 => \N__33127\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32940\,
            in2 => \N__26336\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26729\,
            in2 => \N__33259\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33135\,
            in2 => \N__29825\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26720\,
            in2 => \N__33260\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33139\,
            in2 => \N__26327\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26711\,
            in2 => \N__33261\,
            in3 => \N__26303\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33143\,
            in2 => \N__26462\,
            in3 => \N__26438\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26738\,
            in2 => \N__33262\,
            in3 => \N__26423\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33147\,
            in2 => \N__26507\,
            in3 => \N__26408\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33148\,
            in2 => \N__26483\,
            in3 => \N__26393\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27137\,
            in2 => \N__33263\,
            in3 => \N__26378\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33152\,
            in2 => \N__27203\,
            in3 => \N__26363\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33788\,
            in2 => \N__33264\,
            in3 => \N__26348\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33156\,
            in2 => \N__26672\,
            in3 => \N__26345\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26843\,
            in2 => \N__33265\,
            in3 => \N__26591\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33160\,
            in2 => \N__26588\,
            in3 => \N__26573\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__33161\,
            in1 => \N__33492\,
            in2 => \_gnd_net_\,
            in3 => \N__26570\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33186\,
            in1 => \N__33567\,
            in2 => \N__26567\,
            in3 => \N__26527\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__33571\,
            in1 => \N__33180\,
            in2 => \N__30073\,
            in3 => \N__30094\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30491\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32234\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__27011\,
            in1 => \N__33572\,
            in2 => \N__33270\,
            in3 => \N__27055\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__33568\,
            in1 => \N__33184\,
            in2 => \N__30416\,
            in3 => \N__30370\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__33179\,
            in1 => \N__33570\,
            in2 => \N__30337\,
            in3 => \N__30311\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__33569\,
            in1 => \N__33185\,
            in2 => \N__29488\,
            in3 => \N__29533\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__33590\,
            in1 => \N__29965\,
            in2 => \N__33271\,
            in3 => \N__30006\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__30130\,
            in1 => \N__33591\,
            in2 => \N__33293\,
            in3 => \N__30169\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__30303\,
            in1 => \N__26988\,
            in2 => \_gnd_net_\,
            in3 => \N__30327\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__26987\,
            in1 => \N__30168\,
            in2 => \_gnd_net_\,
            in3 => \N__30126\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__33594\,
            in1 => \N__27128\,
            in2 => \N__27085\,
            in3 => \N__33281\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__26986\,
            in1 => \N__30249\,
            in2 => \_gnd_net_\,
            in3 => \N__30195\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__33592\,
            in1 => \N__26605\,
            in2 => \N__26648\,
            in3 => \N__33285\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__26647\,
            in1 => \N__33593\,
            in2 => \N__26609\,
            in3 => \N__33187\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__33290\,
            in1 => \N__33596\,
            in2 => \N__27158\,
            in3 => \N__27190\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__27191\,
            in1 => \N__33291\,
            in2 => \N__33616\,
            in3 => \N__27154\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \N__33287\,
            in1 => \N__27127\,
            in2 => \N__27084\,
            in3 => \N__33602\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__33595\,
            in1 => \N__33289\,
            in2 => \N__27056\,
            in3 => \N__27010\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__26992\,
            in1 => \N__32460\,
            in2 => \_gnd_net_\,
            in3 => \N__32499\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33286\,
            in1 => \N__33600\,
            in2 => \N__33859\,
            in3 => \N__33810\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__33601\,
            in1 => \N__30580\,
            in2 => \N__30539\,
            in3 => \N__33288\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26818\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48656\,
            ce => 'H',
            sr => \N__48258\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34337\,
            in1 => \N__27257\,
            in2 => \N__31004\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_11_23_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27251\,
            in2 => \N__31013\,
            in3 => \N__34271\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34313\,
            in1 => \N__27245\,
            in2 => \N__30992\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27239\,
            in2 => \N__30656\,
            in3 => \N__34247\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27233\,
            in2 => \N__30647\,
            in3 => \N__34292\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34004\,
            in1 => \N__27227\,
            in2 => \N__30638\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27221\,
            in2 => \N__30629\,
            in3 => \N__34025\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34046\,
            in1 => \N__27215\,
            in2 => \N__30617\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34067\,
            in1 => \N__27209\,
            in2 => \N__30983\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_11_24_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27398\,
            in2 => \N__30806\,
            in3 => \N__34088\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27392\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48650\,
            ce => 'H',
            sr => \N__48267\
        );

    \phase_controller_inst2.S1_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31085\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48646\,
            ce => 'H',
            sr => \N__48280\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30714\,
            in1 => \N__30770\,
            in2 => \_gnd_net_\,
            in3 => \N__41893\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48779\,
            ce => \N__36593\,
            sr => \N__48127\
        );

    \phase_controller_inst1.stoper_hc.target_time_26_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41892\,
            in1 => \N__28530\,
            in2 => \_gnd_net_\,
            in3 => \N__28591\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48779\,
            ce => \N__36593\,
            sr => \N__48127\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27332\,
            in1 => \N__27305\,
            in2 => \_gnd_net_\,
            in3 => \N__41894\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48779\,
            ce => \N__36593\,
            sr => \N__48127\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35075\,
            in2 => \_gnd_net_\,
            in3 => \N__27834\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35076\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27835\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27818\,
            in2 => \N__27266\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36542\,
            in1 => \N__27530\,
            in2 => \_gnd_net_\,
            in3 => \N__27518\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__48761\,
            ce => 'H',
            sr => \N__48137\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__36546\,
            in1 => \N__27503\,
            in2 => \N__27515\,
            in3 => \N__27491\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__48761\,
            ce => 'H',
            sr => \N__48137\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36543\,
            in1 => \N__27488\,
            in2 => \_gnd_net_\,
            in3 => \N__27476\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__48761\,
            ce => 'H',
            sr => \N__48137\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36547\,
            in1 => \N__27473\,
            in2 => \_gnd_net_\,
            in3 => \N__27461\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__48761\,
            ce => 'H',
            sr => \N__48137\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36544\,
            in1 => \N__27458\,
            in2 => \_gnd_net_\,
            in3 => \N__27446\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__48761\,
            ce => 'H',
            sr => \N__48137\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36548\,
            in1 => \N__27443\,
            in2 => \_gnd_net_\,
            in3 => \N__27431\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__48761\,
            ce => 'H',
            sr => \N__48137\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36545\,
            in1 => \N__27428\,
            in2 => \_gnd_net_\,
            in3 => \N__27416\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__48761\,
            ce => 'H',
            sr => \N__48137\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36573\,
            in1 => \N__27413\,
            in2 => \_gnd_net_\,
            in3 => \N__27401\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__48747\,
            ce => 'H',
            sr => \N__48142\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36558\,
            in1 => \N__27650\,
            in2 => \_gnd_net_\,
            in3 => \N__27638\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__48747\,
            ce => 'H',
            sr => \N__48142\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36570\,
            in1 => \N__27635\,
            in2 => \_gnd_net_\,
            in3 => \N__27623\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__48747\,
            ce => 'H',
            sr => \N__48142\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36559\,
            in1 => \N__27620\,
            in2 => \_gnd_net_\,
            in3 => \N__27608\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__48747\,
            ce => 'H',
            sr => \N__48142\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36571\,
            in1 => \N__27605\,
            in2 => \_gnd_net_\,
            in3 => \N__27593\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__48747\,
            ce => 'H',
            sr => \N__48142\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36560\,
            in1 => \N__27590\,
            in2 => \_gnd_net_\,
            in3 => \N__27578\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__48747\,
            ce => 'H',
            sr => \N__48142\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36572\,
            in1 => \N__27575\,
            in2 => \_gnd_net_\,
            in3 => \N__27563\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__48747\,
            ce => 'H',
            sr => \N__48142\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36561\,
            in1 => \N__31164\,
            in2 => \_gnd_net_\,
            in3 => \N__27560\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__48747\,
            ce => 'H',
            sr => \N__48142\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36562\,
            in1 => \N__31218\,
            in2 => \_gnd_net_\,
            in3 => \N__27557\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__48735\,
            ce => 'H',
            sr => \N__48151\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36577\,
            in1 => \N__27549\,
            in2 => \_gnd_net_\,
            in3 => \N__27533\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__48735\,
            ce => 'H',
            sr => \N__48151\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36563\,
            in1 => \N__27774\,
            in2 => \_gnd_net_\,
            in3 => \N__27758\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__48735\,
            ce => 'H',
            sr => \N__48151\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36578\,
            in1 => \N__31425\,
            in2 => \_gnd_net_\,
            in3 => \N__27755\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__48735\,
            ce => 'H',
            sr => \N__48151\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36564\,
            in1 => \N__31445\,
            in2 => \_gnd_net_\,
            in3 => \N__27752\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__48735\,
            ce => 'H',
            sr => \N__48151\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36579\,
            in1 => \N__31660\,
            in2 => \_gnd_net_\,
            in3 => \N__27749\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__48735\,
            ce => 'H',
            sr => \N__48151\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36565\,
            in1 => \N__31642\,
            in2 => \_gnd_net_\,
            in3 => \N__27746\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__48735\,
            ce => 'H',
            sr => \N__48151\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36580\,
            in1 => \N__27735\,
            in2 => \_gnd_net_\,
            in3 => \N__27713\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__48735\,
            ce => 'H',
            sr => \N__48151\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36566\,
            in1 => \N__27702\,
            in2 => \_gnd_net_\,
            in3 => \N__27680\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__48725\,
            ce => 'H',
            sr => \N__48159\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36574\,
            in1 => \N__27667\,
            in2 => \_gnd_net_\,
            in3 => \N__27653\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__48725\,
            ce => 'H',
            sr => \N__48159\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36567\,
            in1 => \N__27922\,
            in2 => \_gnd_net_\,
            in3 => \N__27908\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__48725\,
            ce => 'H',
            sr => \N__48159\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36575\,
            in1 => \N__31265\,
            in2 => \_gnd_net_\,
            in3 => \N__27905\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__48725\,
            ce => 'H',
            sr => \N__48159\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36568\,
            in1 => \N__31304\,
            in2 => \_gnd_net_\,
            in3 => \N__27902\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__48725\,
            ce => 'H',
            sr => \N__48159\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36576\,
            in1 => \N__27896\,
            in2 => \_gnd_net_\,
            in3 => \N__27878\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__48725\,
            ce => 'H',
            sr => \N__48159\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36569\,
            in1 => \N__27856\,
            in2 => \_gnd_net_\,
            in3 => \N__27875\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48725\,
            ce => 'H',
            sr => \N__48159\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__46202\,
            in1 => \N__42284\,
            in2 => \N__44733\,
            in3 => \N__46701\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48715\,
            ce => 'H',
            sr => \N__48167\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__36469\,
            in1 => \N__27842\,
            in2 => \N__35093\,
            in3 => \N__27813\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48715\,
            ce => 'H',
            sr => \N__48167\
        );

    \phase_controller_inst2.start_timer_hc_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__28278\,
            in1 => \N__31097\,
            in2 => \N__42968\,
            in3 => \N__27794\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48715\,
            ce => 'H',
            sr => \N__48167\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28279\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48715\,
            ce => 'H',
            sr => \N__48167\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__28196\,
            in1 => \N__28301\,
            in2 => \_gnd_net_\,
            in3 => \N__28277\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000001010"
        )
    port map (
            in0 => \N__31800\,
            in1 => \N__28238\,
            in2 => \N__28214\,
            in3 => \N__28197\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48715\,
            ce => 'H',
            sr => \N__48167\
        );

    \phase_controller_inst2.stoper_hc.target_time_27_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28173\,
            in1 => \N__28130\,
            in2 => \_gnd_net_\,
            in3 => \N__41854\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48705\,
            ce => \N__28510\,
            sr => \N__48176\
        );

    \phase_controller_inst2.stoper_hc.target_time_28_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41853\,
            in1 => \N__31890\,
            in2 => \_gnd_net_\,
            in3 => \N__31910\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48705\,
            ce => \N__28510\,
            sr => \N__48176\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__28027\,
            in1 => \N__28090\,
            in2 => \N__28073\,
            in3 => \N__28051\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__28091\,
            in1 => \N__28069\,
            in2 => \N__28052\,
            in3 => \N__28028\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__27987\,
            in1 => \N__27970\,
            in2 => \N__28604\,
            in3 => \N__27941\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__27940\,
            in1 => \N__27988\,
            in2 => \N__27974\,
            in3 => \N__28600\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_24_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38204\,
            in1 => \N__38256\,
            in2 => \_gnd_net_\,
            in3 => \N__41857\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48697\,
            ce => \N__28507\,
            sr => \N__48186\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28743\,
            in1 => \N__28705\,
            in2 => \_gnd_net_\,
            in3 => \N__41856\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48697\,
            ce => \N__28507\,
            sr => \N__48186\
        );

    \phase_controller_inst2.stoper_hc.target_time_25_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41855\,
            in1 => \N__28667\,
            in2 => \_gnd_net_\,
            in3 => \N__28646\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48697\,
            ce => \N__28507\,
            sr => \N__48186\
        );

    \phase_controller_inst2.stoper_hc.target_time_26_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28584\,
            in1 => \N__28538\,
            in2 => \_gnd_net_\,
            in3 => \N__41858\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48697\,
            ce => \N__28507\,
            sr => \N__48186\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__28462\,
            in1 => \N__28451\,
            in2 => \N__28430\,
            in3 => \N__28393\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28367\,
            in2 => \N__33632\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28317\,
            in2 => \N__28343\,
            in3 => \N__31983\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31984\,
            in1 => \N__32756\,
            in2 => \N__29735\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29744\,
            in2 => \N__32910\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32760\,
            in2 => \N__32351\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28784\,
            in2 => \N__32911\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32764\,
            in2 => \N__29552\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29648\,
            in2 => \N__32912\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32851\,
            in2 => \N__28772\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28754\,
            in2 => \N__33065\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32855\,
            in2 => \N__30353\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30425\,
            in2 => \N__33066\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32859\,
            in2 => \N__32267\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32522\,
            in2 => \N__33067\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32863\,
            in2 => \N__32531\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28805\,
            in2 => \N__33068\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32941\,
            in2 => \N__29462\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32432\,
            in2 => \N__33128\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32945\,
            in2 => \N__29948\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30182\,
            in2 => \N__33129\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32949\,
            in2 => \N__30110\,
            in3 => \N__28787\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28991\,
            in2 => \N__33130\,
            in3 => \N__28970\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32953\,
            in2 => \N__30275\,
            in3 => \N__28958\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30026\,
            in2 => \N__33131\,
            in3 => \N__28946\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33029\,
            in2 => \N__28943\,
            in3 => \N__28913\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28910\,
            in2 => \N__33191\,
            in3 => \N__28883\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33033\,
            in2 => \N__28880\,
            in3 => \N__28853\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28850\,
            in2 => \N__33192\,
            in3 => \N__28826\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33037\,
            in2 => \N__28823\,
            in3 => \N__28808\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30509\,
            in2 => \N__33193\,
            in3 => \N__29420\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33041\,
            in2 => \N__32540\,
            in3 => \N__29417\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101010011"
        )
    port map (
            in0 => \N__29414\,
            in1 => \N__29402\,
            in2 => \N__29318\,
            in3 => \N__29393\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__29378\,
            in1 => \N__29372\,
            in2 => \_gnd_net_\,
            in3 => \N__29312\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__29313\,
            in1 => \N__29354\,
            in2 => \_gnd_net_\,
            in3 => \N__29348\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__29330\,
            in1 => \N__29324\,
            in2 => \_gnd_net_\,
            in3 => \N__29314\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29928\,
            in2 => \N__29915\,
            in3 => \N__29158\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_199_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111010"
        )
    port map (
            in0 => \N__29159\,
            in1 => \_gnd_net_\,
            in2 => \N__29933\,
            in3 => \N__29914\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48671\,
            ce => 'H',
            sr => \N__48223\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29927\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29929\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29910\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_198_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33166\,
            in1 => \N__33406\,
            in2 => \N__32482\,
            in3 => \N__32515\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__33401\,
            in1 => \N__33167\,
            in2 => \N__29815\,
            in3 => \N__29767\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__32632\,
            in1 => \N__33400\,
            in2 => \N__33266\,
            in3 => \N__32674\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__33404\,
            in1 => \N__33169\,
            in2 => \N__29720\,
            in3 => \N__29692\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33168\,
            in1 => \N__33403\,
            in2 => \N__29635\,
            in3 => \N__29575\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__33405\,
            in1 => \N__33165\,
            in2 => \N__29537\,
            in3 => \N__29489\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__33668\,
            in1 => \N__33402\,
            in2 => \_gnd_net_\,
            in3 => \N__33677\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33435\,
            in1 => \N__30581\,
            in2 => \N__33267\,
            in3 => \N__30538\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33434\,
            in1 => \N__30499\,
            in2 => \N__33269\,
            in3 => \N__30451\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33433\,
            in1 => \N__30412\,
            in2 => \N__33268\,
            in3 => \N__30374\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__33453\,
            in1 => \N__33114\,
            in2 => \N__30338\,
            in3 => \N__30310\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33120\,
            in1 => \N__33451\,
            in2 => \N__30260\,
            in3 => \N__30202\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__33452\,
            in1 => \N__33118\,
            in2 => \N__30170\,
            in3 => \N__30131\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__30095\,
            in1 => \N__33454\,
            in2 => \N__33258\,
            in3 => \N__30074\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__33450\,
            in1 => \N__33119\,
            in2 => \N__30014\,
            in3 => \N__29969\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33971\,
            in1 => \N__34333\,
            in2 => \_gnd_net_\,
            in3 => \N__30608\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_12_21_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__48655\,
            ce => 'H',
            sr => \N__48244\
        );

    \pwm_generator_inst.counter_1_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33965\,
            in1 => \N__34270\,
            in2 => \_gnd_net_\,
            in3 => \N__30605\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__48655\,
            ce => 'H',
            sr => \N__48244\
        );

    \pwm_generator_inst.counter_2_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33972\,
            in1 => \N__34312\,
            in2 => \_gnd_net_\,
            in3 => \N__30602\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__48655\,
            ce => 'H',
            sr => \N__48244\
        );

    \pwm_generator_inst.counter_3_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33966\,
            in1 => \N__34246\,
            in2 => \_gnd_net_\,
            in3 => \N__30599\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__48655\,
            ce => 'H',
            sr => \N__48244\
        );

    \pwm_generator_inst.counter_4_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33973\,
            in1 => \N__34291\,
            in2 => \_gnd_net_\,
            in3 => \N__30596\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__48655\,
            ce => 'H',
            sr => \N__48244\
        );

    \pwm_generator_inst.counter_5_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33967\,
            in1 => \N__34002\,
            in2 => \_gnd_net_\,
            in3 => \N__30593\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__48655\,
            ce => 'H',
            sr => \N__48244\
        );

    \pwm_generator_inst.counter_6_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33974\,
            in1 => \N__34023\,
            in2 => \_gnd_net_\,
            in3 => \N__30590\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__48655\,
            ce => 'H',
            sr => \N__48244\
        );

    \pwm_generator_inst.counter_7_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33968\,
            in1 => \N__34045\,
            in2 => \_gnd_net_\,
            in3 => \N__30587\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__48655\,
            ce => 'H',
            sr => \N__48244\
        );

    \pwm_generator_inst.counter_8_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33970\,
            in1 => \N__34066\,
            in2 => \_gnd_net_\,
            in3 => \N__30584\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_12_22_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__48652\,
            ce => 'H',
            sr => \N__48251\
        );

    \pwm_generator_inst.counter_9_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__34087\,
            in1 => \N__33969\,
            in2 => \_gnd_net_\,
            in3 => \N__30698\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48652\,
            ce => 'H',
            sr => \N__48251\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48958\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48649\,
            ce => 'H',
            sr => \N__48259\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__35321\,
            in1 => \N__30679\,
            in2 => \_gnd_net_\,
            in3 => \N__30859\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__30695\,
            in1 => \N__30680\,
            in2 => \N__30895\,
            in3 => \N__35320\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__47463\,
            in1 => \N__47537\,
            in2 => \N__30896\,
            in3 => \N__34397\,
            lcout => \pwm_generator_inst.threshold_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__47472\,
            in1 => \N__47541\,
            in2 => \N__30899\,
            in3 => \N__34388\,
            lcout => \pwm_generator_inst.threshold_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__47542\,
            in1 => \N__47473\,
            in2 => \N__34379\,
            in3 => \N__30877\,
            lcout => \pwm_generator_inst.threshold_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__47474\,
            in1 => \N__47543\,
            in2 => \N__30898\,
            in3 => \N__34367\,
            lcout => \pwm_generator_inst.un14_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110101"
        )
    port map (
            in0 => \N__47544\,
            in1 => \N__47475\,
            in2 => \N__30900\,
            in3 => \N__34358\,
            lcout => \pwm_generator_inst.un14_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110101"
        )
    port map (
            in0 => \N__47539\,
            in1 => \N__47470\,
            in2 => \N__34421\,
            in3 => \N__30869\,
            lcout => \pwm_generator_inst.un14_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__47469\,
            in1 => \N__47538\,
            in2 => \N__30897\,
            in3 => \N__33869\,
            lcout => \pwm_generator_inst.threshold_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__47540\,
            in1 => \N__47471\,
            in2 => \N__34409\,
            in3 => \N__30870\,
            lcout => \pwm_generator_inst.threshold_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__47545\,
            in1 => \N__30891\,
            in2 => \N__34349\,
            in3 => \N__47477\,
            lcout => \pwm_generator_inst.un14_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__47476\,
            in1 => \N__47546\,
            in2 => \N__30939\,
            in3 => \N__34472\,
            lcout => \pwm_generator_inst.threshold_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48308\,
            lcout => \pll_inst.red_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__31234\,
            in1 => \N__31223\,
            in2 => \N__31195\,
            in3 => \N__31169\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30718\,
            in1 => \N__30768\,
            in2 => \_gnd_net_\,
            in3 => \N__41889\,
            lcout => \elapsed_time_ns_1_RNI13CN9_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__31235\,
            in1 => \N__31222\,
            in2 => \N__31196\,
            in3 => \N__31168\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__31733\,
            in1 => \N__31837\,
            in2 => \N__31115\,
            in3 => \N__31127\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48770\,
            ce => 'H',
            sr => \N__48132\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000010101010"
        )
    port map (
            in0 => \N__31126\,
            in1 => \N__35603\,
            in2 => \N__35237\,
            in3 => \N__35174\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48770\,
            ce => 'H',
            sr => \N__48132\
        );

    \phase_controller_inst2.state_RNI9M3O_0_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31125\,
            in2 => \_gnd_net_\,
            in3 => \N__31111\,
            lcout => \phase_controller_inst2.state_RNI9M3OZ0Z_0\,
            ltout => \phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_3_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__31069\,
            in1 => \N__31052\,
            in2 => \N__31100\,
            in3 => \N__36283\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48770\,
            ce => 'H',
            sr => \N__48132\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31050\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31067\,
            lcout => \phase_controller_inst2.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_ns_i_a3_1_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43006\,
            in2 => \_gnd_net_\,
            in3 => \N__42941\,
            lcout => state_ns_i_a3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_2_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__31068\,
            in1 => \N__31051\,
            in2 => \N__31761\,
            in3 => \N__31805\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48770\,
            ce => 'H',
            sr => \N__48132\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__31550\,
            in1 => \N__31466\,
            in2 => \N__31661\,
            in3 => \N__31641\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__31465\,
            in1 => \N__31659\,
            in2 => \N__31643\,
            in3 => \N__31549\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_23_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31613\,
            in1 => \N__31589\,
            in2 => \_gnd_net_\,
            in3 => \N__41860\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48762\,
            ce => \N__36531\,
            sr => \N__48138\
        );

    \phase_controller_inst1.stoper_hc.target_time_22_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31541\,
            in1 => \N__31511\,
            in2 => \_gnd_net_\,
            in3 => \N__41859\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48762\,
            ce => \N__36531\,
            sr => \N__48138\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__31444\,
            in1 => \N__31426\,
            in2 => \N__31394\,
            in3 => \N__31313\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__31312\,
            in1 => \N__31443\,
            in2 => \N__31430\,
            in3 => \N__31390\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_21_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41420\,
            in1 => \N__41945\,
            in2 => \_gnd_net_\,
            in3 => \N__41821\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48749\,
            ce => \N__36538\,
            sr => \N__48143\
        );

    \phase_controller_inst1.stoper_hc.target_time_20_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31382\,
            in1 => \N__31358\,
            in2 => \_gnd_net_\,
            in3 => \N__41820\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48749\,
            ce => \N__36538\,
            sr => \N__48143\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__31852\,
            in1 => \N__31302\,
            in2 => \N__31286\,
            in3 => \N__31263\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31891\,
            in1 => \N__31906\,
            in2 => \_gnd_net_\,
            in3 => \N__41851\,
            lcout => \elapsed_time_ns_1_RNI69DN9_0_28\,
            ltout => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_28_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__41852\,
            in1 => \_gnd_net_\,
            in2 => \N__31895\,
            in3 => \N__31892\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48737\,
            ce => \N__36594\,
            sr => \N__48152\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__31841\,
            in1 => \N__31799\,
            in2 => \N__31772\,
            in3 => \N__31731\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__35190\,
            in1 => \N__31685\,
            in2 => \N__31676\,
            in3 => \N__42966\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48727\,
            ce => 'H',
            sr => \N__48160\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__35216\,
            in1 => \N__31672\,
            in2 => \_gnd_net_\,
            in3 => \N__35189\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101011111010"
        )
    port map (
            in0 => \N__31673\,
            in1 => \N__35599\,
            in2 => \N__35172\,
            in3 => \N__35218\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48727\,
            ce => 'H',
            sr => \N__48160\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101110101"
        )
    port map (
            in0 => \N__35217\,
            in1 => \N__32033\,
            in2 => \N__35638\,
            in3 => \N__35615\,
            lcout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31664\,
            in3 => \N__35156\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35191\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48727\,
            ce => 'H',
            sr => \N__48160\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35157\,
            in2 => \_gnd_net_\,
            in3 => \N__35131\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__31921\,
            in1 => \N__31934\,
            in2 => \N__35885\,
            in3 => \N__35863\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__31933\,
            in1 => \N__35862\,
            in2 => \N__31925\,
            in3 => \N__35883\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42266\,
            in1 => \N__42170\,
            in2 => \_gnd_net_\,
            in3 => \N__47120\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48718\,
            ce => \N__46110\,
            sr => \N__48168\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43622\,
            in1 => \N__43592\,
            in2 => \_gnd_net_\,
            in3 => \N__47121\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48718\,
            ce => \N__46110\,
            sr => \N__48168\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47116\,
            in1 => \N__42224\,
            in2 => \_gnd_net_\,
            in3 => \N__42527\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48708\,
            ce => \N__46112\,
            sr => \N__48177\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43409\,
            in1 => \N__43383\,
            in2 => \_gnd_net_\,
            in3 => \N__47117\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48708\,
            ce => \N__46112\,
            sr => \N__48177\
        );

    \phase_controller_inst2.stoper_tr.target_time_29_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42449\,
            in1 => \N__42425\,
            in2 => \_gnd_net_\,
            in3 => \N__47119\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48708\,
            ce => \N__46112\,
            sr => \N__48177\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44813\,
            in1 => \N__44787\,
            in2 => \_gnd_net_\,
            in3 => \N__47118\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48708\,
            ce => \N__46112\,
            sr => \N__48177\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__35958\,
            in1 => \N__32054\,
            in2 => \N__35984\,
            in3 => \N__32042\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__32041\,
            in1 => \N__35982\,
            in2 => \N__35963\,
            in3 => \N__32053\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_28_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44232\,
            in1 => \N__43808\,
            in2 => \_gnd_net_\,
            in3 => \N__47122\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48699\,
            ce => \N__46113\,
            sr => \N__48187\
        );

    \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100000100"
        )
    port map (
            in0 => \N__36213\,
            in1 => \N__32023\,
            in2 => \N__44138\,
            in3 => \N__36041\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__32022\,
            in1 => \N__44136\,
            in2 => \N__36046\,
            in3 => \N__36212\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_30_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45788\,
            in1 => \N__45806\,
            in2 => \_gnd_net_\,
            in3 => \N__47115\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48691\,
            ce => \N__46115\,
            sr => \N__48196\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__32024\,
            in1 => \N__44137\,
            in2 => \N__36047\,
            in3 => \N__36214\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42199\,
            in1 => \N__38584\,
            in2 => \_gnd_net_\,
            in3 => \N__47112\,
            lcout => \elapsed_time_ns_1_RNI0AOBB_0_13\,
            ltout => \elapsed_time_ns_1_RNI0AOBB_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__47113\,
            in1 => \_gnd_net_\,
            in2 => \N__32012\,
            in3 => \N__42200\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48691\,
            ce => \N__46115\,
            sr => \N__48196\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47114\,
            in1 => \N__46298\,
            in2 => \_gnd_net_\,
            in3 => \N__46337\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48691\,
            ce => \N__46115\,
            sr => \N__48196\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__32009\,
            in1 => \N__33079\,
            in2 => \N__31988\,
            in3 => \N__33470\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33468\,
            in1 => \N__32248\,
            in2 => \N__33219\,
            in3 => \N__32194\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33467\,
            in1 => \N__32156\,
            in2 => \N__33218\,
            in3 => \N__32117\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__32516\,
            in1 => \N__33075\,
            in2 => \N__32483\,
            in3 => \N__33469\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33466\,
            in1 => \N__32422\,
            in2 => \N__33220\,
            in3 => \N__32374\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33515\,
            in1 => \N__32339\,
            in2 => \N__33221\,
            in3 => \N__32294\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33086\,
            in1 => \N__33517\,
            in2 => \N__32252\,
            in3 => \N__32195\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__33516\,
            in1 => \N__32155\,
            in2 => \N__33222\,
            in3 => \N__32113\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32072\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48681\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011001100"
        )
    port map (
            in0 => \N__35120\,
            in1 => \N__42699\,
            in2 => \N__42340\,
            in3 => \N__35092\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48677\,
            ce => 'H',
            sr => \N__48218\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__33223\,
            in1 => \N__33385\,
            in2 => \N__33863\,
            in3 => \N__33815\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33779\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48672\,
            ce => \N__33736\,
            sr => \N__48224\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33713\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33383\,
            in2 => \N__33671\,
            in3 => \N__33667\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__33384\,
            in1 => \N__33224\,
            in2 => \N__32678\,
            in3 => \N__32636\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36845\,
            in2 => \_gnd_net_\,
            in3 => \N__36866\,
            lcout => \current_shift_inst.timer_s1.N_162_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__36847\,
            in1 => \N__36867\,
            in2 => \_gnd_net_\,
            in3 => \N__39335\,
            lcout => \current_shift_inst.timer_s1.N_163_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34332\,
            in2 => \_gnd_net_\,
            in3 => \N__34308\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__34290\,
            in1 => \N__34269\,
            in2 => \N__34250\,
            in3 => \N__34245\,
            lcout => \pwm_generator_inst.un1_counterlt9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36846\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__34086\,
            in1 => \N__34062\,
            in2 => \_gnd_net_\,
            in3 => \N__34044\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__34024\,
            in1 => \N__34003\,
            in2 => \N__33983\,
            in3 => \N__33980\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33935\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48653\,
            ce => 'H',
            sr => \N__48252\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39893\,
            in2 => \_gnd_net_\,
            in3 => \N__39873\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48653\,
            ce => 'H',
            sr => \N__48252\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33902\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48653\,
            ce => 'H',
            sr => \N__48252\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34442\,
            in2 => \N__37310\,
            in3 => \N__37305\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37223\,
            in2 => \_gnd_net_\,
            in3 => \N__34412\,
            lcout => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34430\,
            in2 => \_gnd_net_\,
            in3 => \N__34400\,
            lcout => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34460\,
            in2 => \_gnd_net_\,
            in3 => \N__34391\,
            lcout => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34448\,
            in2 => \_gnd_net_\,
            in3 => \N__34382\,
            lcout => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34466\,
            in2 => \_gnd_net_\,
            in3 => \N__34370\,
            lcout => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34454\,
            in2 => \_gnd_net_\,
            in3 => \N__34361\,
            lcout => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34763\,
            in2 => \_gnd_net_\,
            in3 => \N__34352\,
            lcout => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34436\,
            in2 => \_gnd_net_\,
            in3 => \N__34340\,
            lcout => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\,
            ltout => OPEN,
            carryin => \bfn_13_25_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__37481\,
            in1 => \N__37514\,
            in2 => \N__37309\,
            in3 => \N__34475\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100001110100"
        )
    port map (
            in0 => \N__37439\,
            in1 => \N__37298\,
            in2 => \N__37985\,
            in3 => \N__37184\,
            lcout => \pwm_generator_inst.un19_threshold_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__37202\,
            in1 => \N__40778\,
            in2 => \N__40763\,
            in3 => \N__37288\,
            lcout => \pwm_generator_inst.un19_threshold_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__37952\,
            in1 => \N__37154\,
            in2 => \N__37307\,
            in3 => \N__37175\,
            lcout => \pwm_generator_inst.un19_threshold_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__37193\,
            in1 => \N__41375\,
            in2 => \N__37306\,
            in3 => \N__41393\,
            lcout => \pwm_generator_inst.un19_threshold_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__44423\,
            in1 => \N__37319\,
            in2 => \N__44402\,
            in3 => \N__37284\,
            lcout => \pwm_generator_inst.un19_threshold_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__37538\,
            in1 => \N__37297\,
            in2 => \N__37472\,
            in3 => \N__37133\,
            lcout => \pwm_generator_inst.un19_threshold_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__37358\,
            in1 => \N__37211\,
            in2 => \N__37418\,
            in3 => \N__37296\,
            lcout => \pwm_generator_inst.un19_threshold_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37948\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37174\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__37142\,
            in1 => \N__37928\,
            in2 => \N__37308\,
            in3 => \N__37454\,
            lcout => \pwm_generator_inst.un19_threshold_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_axb_4_LC_13_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34754\,
            in2 => \N__34733\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_13_28_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_13_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34715\,
            in2 => \N__34697\,
            in3 => \N__34679\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_13_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34676\,
            in2 => \N__34655\,
            in3 => \N__34637\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_13_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34634\,
            in2 => \N__34616\,
            in3 => \N__34595\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_13_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34592\,
            in2 => \N__34574\,
            in3 => \N__34559\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_13_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34556\,
            in2 => \N__34541\,
            in3 => \N__34520\,
            lcout => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34517\,
            in2 => \N__34499\,
            in3 => \N__34478\,
            lcout => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_13_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34994\,
            in2 => \N__34976\,
            in3 => \N__34958\,
            lcout => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34955\,
            in2 => \N__34934\,
            in3 => \N__34916\,
            lcout => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \bfn_13_29_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_13_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34913\,
            in2 => \N__34892\,
            in3 => \N__34874\,
            lcout => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_13_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34871\,
            in2 => \N__35322\,
            in3 => \N__34853\,
            lcout => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_13_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35311\,
            in2 => \N__34850\,
            in3 => \N__34829\,
            lcout => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_13_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34826\,
            in2 => \N__35323\,
            in3 => \N__34808\,
            lcout => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_13_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35315\,
            in2 => \N__34805\,
            in3 => \N__34787\,
            lcout => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_13_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34784\,
            in2 => \N__35324\,
            in3 => \N__34766\,
            lcout => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_13_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35319\,
            in2 => \N__35273\,
            in3 => \N__35255\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_13_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__38267\,
            in1 => \N__35252\,
            in2 => \_gnd_net_\,
            in3 => \N__35240\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35236\,
            in2 => \_gnd_net_\,
            in3 => \N__35201\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__42392\,
            in1 => \N__42348\,
            in2 => \_gnd_net_\,
            in3 => \N__35041\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__35173\,
            in1 => \N__35138\,
            in2 => \N__35578\,
            in3 => \N__36120\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48782\,
            ce => 'H',
            sr => \N__48128\
        );

    \phase_controller_inst1.stoper_hc.running_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111110000"
        )
    port map (
            in0 => \N__42356\,
            in1 => \N__35116\,
            in2 => \N__35045\,
            in3 => \N__35074\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48782\,
            ce => 'H',
            sr => \N__48128\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38150\,
            in2 => \N__35030\,
            in3 => \N__35568\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35021\,
            in2 => \N__35009\,
            in3 => \N__35552\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35000\,
            in2 => \N__41327\,
            in3 => \N__35525\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38351\,
            in2 => \N__35393\,
            in3 => \N__35507\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38345\,
            in2 => \N__35384\,
            in3 => \N__35828\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35807\,
            in1 => \N__35375\,
            in2 => \N__38339\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35369\,
            in2 => \N__38171\,
            in3 => \N__35789\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38156\,
            in2 => \N__35363\,
            in3 => \N__35771\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38162\,
            in2 => \N__35354\,
            in3 => \N__35753\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38435\,
            in2 => \N__35345\,
            in3 => \N__35735\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38618\,
            in2 => \N__35333\,
            in3 => \N__35717\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38630\,
            in2 => \N__35492\,
            in3 => \N__35699\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35939\,
            in1 => \N__35483\,
            in2 => \N__35468\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35921\,
            in1 => \N__35459\,
            in2 => \N__35447\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35438\,
            in2 => \N__35426\,
            in3 => \N__35903\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35417\,
            in2 => \N__35408\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38069\,
            in2 => \N__38144\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38516\,
            in2 => \N__38468\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38369\,
            in2 => \N__38423\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38276\,
            in2 => \N__38330\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41960\,
            in2 => \N__42038\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35681\,
            in2 => \N__35669\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35654\,
            in2 => \N__35642\,
            in3 => \N__35609\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35606\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35585\,
            in2 => \N__35579\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36169\,
            in1 => \N__35551\,
            in2 => \_gnd_net_\,
            in3 => \N__35537\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__48738\,
            ce => 'H',
            sr => \N__48153\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__36173\,
            in1 => \N__35524\,
            in2 => \N__35534\,
            in3 => \N__35510\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__48738\,
            ce => 'H',
            sr => \N__48153\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36170\,
            in1 => \N__35506\,
            in2 => \_gnd_net_\,
            in3 => \N__35831\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__48738\,
            ce => 'H',
            sr => \N__48153\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36174\,
            in1 => \N__35824\,
            in2 => \_gnd_net_\,
            in3 => \N__35810\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__48738\,
            ce => 'H',
            sr => \N__48153\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36171\,
            in1 => \N__35806\,
            in2 => \_gnd_net_\,
            in3 => \N__35792\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__48738\,
            ce => 'H',
            sr => \N__48153\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36175\,
            in1 => \N__35788\,
            in2 => \_gnd_net_\,
            in3 => \N__35774\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__48738\,
            ce => 'H',
            sr => \N__48153\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36172\,
            in1 => \N__35770\,
            in2 => \_gnd_net_\,
            in3 => \N__35756\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__48738\,
            ce => 'H',
            sr => \N__48153\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36124\,
            in1 => \N__35752\,
            in2 => \_gnd_net_\,
            in3 => \N__35738\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__48728\,
            ce => 'H',
            sr => \N__48161\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36183\,
            in1 => \N__35734\,
            in2 => \_gnd_net_\,
            in3 => \N__35720\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__48728\,
            ce => 'H',
            sr => \N__48161\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36121\,
            in1 => \N__35716\,
            in2 => \_gnd_net_\,
            in3 => \N__35702\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__48728\,
            ce => 'H',
            sr => \N__48161\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36184\,
            in1 => \N__35698\,
            in2 => \_gnd_net_\,
            in3 => \N__35684\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__48728\,
            ce => 'H',
            sr => \N__48161\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36122\,
            in1 => \N__35938\,
            in2 => \_gnd_net_\,
            in3 => \N__35924\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__48728\,
            ce => 'H',
            sr => \N__48161\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36185\,
            in1 => \N__35920\,
            in2 => \_gnd_net_\,
            in3 => \N__35906\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__48728\,
            ce => 'H',
            sr => \N__48161\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36123\,
            in1 => \N__35902\,
            in2 => \_gnd_net_\,
            in3 => \N__35888\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__48728\,
            ce => 'H',
            sr => \N__48161\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36186\,
            in1 => \N__35884\,
            in2 => \_gnd_net_\,
            in3 => \N__35867\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__48728\,
            ce => 'H',
            sr => \N__48161\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36187\,
            in1 => \N__35864\,
            in2 => \_gnd_net_\,
            in3 => \N__35846\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__48719\,
            ce => 'H',
            sr => \N__48169\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36191\,
            in1 => \N__38083\,
            in2 => \_gnd_net_\,
            in3 => \N__35843\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__48719\,
            ce => 'H',
            sr => \N__48169\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36188\,
            in1 => \N__38128\,
            in2 => \_gnd_net_\,
            in3 => \N__35840\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__48719\,
            ce => 'H',
            sr => \N__48169\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36192\,
            in1 => \N__38503\,
            in2 => \_gnd_net_\,
            in3 => \N__35837\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__48719\,
            ce => 'H',
            sr => \N__48169\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36189\,
            in1 => \N__38485\,
            in2 => \_gnd_net_\,
            in3 => \N__35834\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__48719\,
            ce => 'H',
            sr => \N__48169\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36193\,
            in1 => \N__38389\,
            in2 => \_gnd_net_\,
            in3 => \N__36002\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__48719\,
            ce => 'H',
            sr => \N__48169\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36190\,
            in1 => \N__38408\,
            in2 => \_gnd_net_\,
            in3 => \N__35999\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__48719\,
            ce => 'H',
            sr => \N__48169\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36194\,
            in1 => \N__38290\,
            in2 => \_gnd_net_\,
            in3 => \N__35996\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__48719\,
            ce => 'H',
            sr => \N__48169\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36176\,
            in1 => \N__38314\,
            in2 => \_gnd_net_\,
            in3 => \N__35993\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__48709\,
            ce => 'H',
            sr => \N__48178\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36180\,
            in1 => \N__41986\,
            in2 => \_gnd_net_\,
            in3 => \N__35990\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__48709\,
            ce => 'H',
            sr => \N__48178\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36177\,
            in1 => \N__42019\,
            in2 => \_gnd_net_\,
            in3 => \N__35987\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__48709\,
            ce => 'H',
            sr => \N__48178\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36181\,
            in1 => \N__35983\,
            in2 => \_gnd_net_\,
            in3 => \N__35966\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__48709\,
            ce => 'H',
            sr => \N__48178\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36178\,
            in1 => \N__35962\,
            in2 => \_gnd_net_\,
            in3 => \N__35942\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__48709\,
            ce => 'H',
            sr => \N__48178\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36182\,
            in1 => \N__36215\,
            in2 => \_gnd_net_\,
            in3 => \N__36197\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__48709\,
            ce => 'H',
            sr => \N__48178\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36179\,
            in1 => \N__36045\,
            in2 => \_gnd_net_\,
            in3 => \N__36050\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48709\,
            ce => 'H',
            sr => \N__48178\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36717\,
            in1 => \N__38562\,
            in2 => \_gnd_net_\,
            in3 => \N__36023\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__48700\,
            ce => \N__43940\,
            sr => \N__48188\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36709\,
            in1 => \N__38535\,
            in2 => \_gnd_net_\,
            in3 => \N__36020\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__48700\,
            ce => \N__43940\,
            sr => \N__48188\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36718\,
            in1 => \N__38833\,
            in2 => \_gnd_net_\,
            in3 => \N__36017\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__48700\,
            ce => \N__43940\,
            sr => \N__48188\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36710\,
            in1 => \N__38809\,
            in2 => \_gnd_net_\,
            in3 => \N__36014\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__48700\,
            ce => \N__43940\,
            sr => \N__48188\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36719\,
            in1 => \N__38785\,
            in2 => \_gnd_net_\,
            in3 => \N__36011\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__48700\,
            ce => \N__43940\,
            sr => \N__48188\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36711\,
            in1 => \N__38761\,
            in2 => \_gnd_net_\,
            in3 => \N__36008\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__48700\,
            ce => \N__43940\,
            sr => \N__48188\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36720\,
            in1 => \N__38737\,
            in2 => \_gnd_net_\,
            in3 => \N__36005\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__48700\,
            ce => \N__43940\,
            sr => \N__48188\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36712\,
            in1 => \N__38713\,
            in2 => \_gnd_net_\,
            in3 => \N__36242\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__48700\,
            ce => \N__43940\,
            sr => \N__48188\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36716\,
            in1 => \N__38689\,
            in2 => \_gnd_net_\,
            in3 => \N__36239\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__48692\,
            ce => \N__43939\,
            sr => \N__48197\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36724\,
            in1 => \N__38665\,
            in2 => \_gnd_net_\,
            in3 => \N__36236\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__48692\,
            ce => \N__43939\,
            sr => \N__48197\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36713\,
            in1 => \N__39023\,
            in2 => \_gnd_net_\,
            in3 => \N__36233\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__48692\,
            ce => \N__43939\,
            sr => \N__48197\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36721\,
            in1 => \N__39001\,
            in2 => \_gnd_net_\,
            in3 => \N__36230\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__48692\,
            ce => \N__43939\,
            sr => \N__48197\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36714\,
            in1 => \N__38979\,
            in2 => \_gnd_net_\,
            in3 => \N__36227\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__48692\,
            ce => \N__43939\,
            sr => \N__48197\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36722\,
            in1 => \N__38953\,
            in2 => \_gnd_net_\,
            in3 => \N__36224\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__48692\,
            ce => \N__43939\,
            sr => \N__48197\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36715\,
            in1 => \N__38929\,
            in2 => \_gnd_net_\,
            in3 => \N__36221\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__48692\,
            ce => \N__43939\,
            sr => \N__48197\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36723\,
            in1 => \N__38905\,
            in2 => \_gnd_net_\,
            in3 => \N__36218\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__48692\,
            ce => \N__43939\,
            sr => \N__48197\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36703\,
            in1 => \N__38881\,
            in2 => \_gnd_net_\,
            in3 => \N__36269\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__48686\,
            ce => \N__43938\,
            sr => \N__48205\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36725\,
            in1 => \N__38857\,
            in2 => \_gnd_net_\,
            in3 => \N__36266\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__48686\,
            ce => \N__43938\,
            sr => \N__48205\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36704\,
            in1 => \N__39244\,
            in2 => \_gnd_net_\,
            in3 => \N__36263\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__48686\,
            ce => \N__43938\,
            sr => \N__48205\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36726\,
            in1 => \N__39220\,
            in2 => \_gnd_net_\,
            in3 => \N__36260\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__48686\,
            ce => \N__43938\,
            sr => \N__48205\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36705\,
            in1 => \N__39196\,
            in2 => \_gnd_net_\,
            in3 => \N__36257\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__48686\,
            ce => \N__43938\,
            sr => \N__48205\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36727\,
            in1 => \N__39172\,
            in2 => \_gnd_net_\,
            in3 => \N__36254\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__48686\,
            ce => \N__43938\,
            sr => \N__48205\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36706\,
            in1 => \N__39148\,
            in2 => \_gnd_net_\,
            in3 => \N__36251\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__48686\,
            ce => \N__43938\,
            sr => \N__48205\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36728\,
            in1 => \N__39124\,
            in2 => \_gnd_net_\,
            in3 => \N__36248\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__48686\,
            ce => \N__43938\,
            sr => \N__48205\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36699\,
            in1 => \N__39100\,
            in2 => \_gnd_net_\,
            in3 => \N__36245\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__48682\,
            ce => \N__43934\,
            sr => \N__48212\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36707\,
            in1 => \N__39076\,
            in2 => \_gnd_net_\,
            in3 => \N__36743\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__48682\,
            ce => \N__43934\,
            sr => \N__48212\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36700\,
            in1 => \N__39056\,
            in2 => \_gnd_net_\,
            in3 => \N__36740\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__48682\,
            ce => \N__43934\,
            sr => \N__48212\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36708\,
            in1 => \N__39418\,
            in2 => \_gnd_net_\,
            in3 => \N__36737\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__48682\,
            ce => \N__43934\,
            sr => \N__48212\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36701\,
            in1 => \N__39040\,
            in2 => \_gnd_net_\,
            in3 => \N__36734\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__48682\,
            ce => \N__43934\,
            sr => \N__48212\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__39434\,
            in1 => \N__36702\,
            in2 => \_gnd_net_\,
            in3 => \N__36731\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48682\,
            ce => \N__43934\,
            sr => \N__48212\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43985\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42344\,
            in2 => \_gnd_net_\,
            in3 => \N__42380\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39294\,
            in2 => \_gnd_net_\,
            in3 => \N__36954\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36323\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48673\,
            ce => 'H',
            sr => \N__48225\
        );

    \phase_controller_inst1.state_3_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__39307\,
            in1 => \N__44564\,
            in2 => \N__36959\,
            in3 => \N__36293\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48673\,
            ce => 'H',
            sr => \N__48225\
        );

    \phase_controller_inst1.state_2_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__36958\,
            in1 => \N__44631\,
            in2 => \N__42710\,
            in3 => \N__39306\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48673\,
            ce => 'H',
            sr => \N__48225\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36935\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48666\,
            ce => 'H',
            sr => \N__48229\
        );

    \current_shift_inst.stop_timer_s1_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__39311\,
            in1 => \N__39333\,
            in2 => \N__36872\,
            in3 => \N__39352\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48662\,
            ce => 'H',
            sr => \N__48234\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36905\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48662\,
            ce => 'H',
            sr => \N__48234\
        );

    \current_shift_inst.timer_s1.running_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__39334\,
            in1 => \N__36868\,
            in2 => \_gnd_net_\,
            in3 => \N__36848\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48662\,
            ce => 'H',
            sr => \N__48234\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36829\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48659\,
            ce => 'H',
            sr => \N__48239\
        );

    \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36785\,
            in2 => \_gnd_net_\,
            in3 => \N__36803\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_14_25_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36761\,
            in2 => \_gnd_net_\,
            in3 => \N__36779\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37127\,
            in2 => \_gnd_net_\,
            in3 => \N__36755\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37103\,
            in2 => \_gnd_net_\,
            in3 => \N__37121\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37079\,
            in2 => \_gnd_net_\,
            in3 => \N__37097\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37055\,
            in2 => \_gnd_net_\,
            in3 => \N__37073\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37031\,
            in2 => \_gnd_net_\,
            in3 => \N__37049\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37013\,
            in2 => \_gnd_net_\,
            in3 => \N__37025\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36989\,
            in2 => \_gnd_net_\,
            in3 => \N__37007\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_14_26_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36965\,
            in2 => \_gnd_net_\,
            in3 => \N__36983\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44395\,
            in2 => \_gnd_net_\,
            in3 => \N__37313\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__37295\,
            in1 => \N__37397\,
            in2 => \_gnd_net_\,
            in3 => \N__37214\,
            lcout => \pwm_generator_inst.un19_threshold_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37413\,
            in2 => \_gnd_net_\,
            in3 => \N__37205\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40749\,
            in2 => \_gnd_net_\,
            in3 => \N__37196\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41367\,
            in2 => \_gnd_net_\,
            in3 => \N__37187\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37434\,
            in2 => \_gnd_net_\,
            in3 => \N__37178\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37170\,
            in2 => \_gnd_net_\,
            in3 => \N__37145\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_14_27_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37452\,
            in2 => \_gnd_net_\,
            in3 => \N__37136\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37467\,
            in2 => \_gnd_net_\,
            in3 => \N__37487\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_14_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37484\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37534\,
            in2 => \_gnd_net_\,
            in3 => \N__37468\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37927\,
            in2 => \_gnd_net_\,
            in3 => \N__37453\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37978\,
            in2 => \_gnd_net_\,
            in3 => \N__37438\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_14_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37354\,
            in2 => \_gnd_net_\,
            in3 => \N__37417\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_LC_14_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37393\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_28_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_14_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37370\,
            in2 => \_gnd_net_\,
            in3 => \N__37343\,
            lcout => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37340\,
            in2 => \_gnd_net_\,
            in3 => \N__37322\,
            lcout => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38009\,
            in2 => \_gnd_net_\,
            in3 => \N__37994\,
            lcout => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_14_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37991\,
            in2 => \_gnd_net_\,
            in3 => \N__37967\,
            lcout => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_14_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37632\,
            in2 => \N__37964\,
            in3 => \N__37937\,
            lcout => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_14_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37934\,
            in2 => \N__37716\,
            in3 => \N__37916\,
            lcout => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_14_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37636\,
            in2 => \N__37547\,
            in3 => \N__37523\,
            lcout => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_14_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37520\,
            in2 => \_gnd_net_\,
            in3 => \N__37502\,
            lcout => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\,
            ltout => OPEN,
            carryin => \bfn_14_29_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_LC_14_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37499\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_LC_14_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37493\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_LC_14_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38063\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_LC_14_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38057\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_LC_14_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38051\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_LC_14_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38045\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_LC_14_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38039\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_LC_14_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38033\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_30_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_LC_14_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38027\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_LC_14_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38021\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_LC_14_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38015\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_14_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38270\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38196\,
            in1 => \N__38261\,
            in2 => \_gnd_net_\,
            in3 => \N__41880\,
            lcout => \elapsed_time_ns_1_RNI25DN9_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47062\,
            in1 => \N__44882\,
            in2 => \_gnd_net_\,
            in3 => \N__44853\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48783\,
            ce => \N__46107\,
            sr => \N__48129\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44372\,
            in1 => \N__44350\,
            in2 => \_gnd_net_\,
            in3 => \N__47064\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48783\,
            ce => \N__46107\,
            sr => \N__48129\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47063\,
            in1 => \N__44937\,
            in2 => \_gnd_net_\,
            in3 => \N__44920\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48783\,
            ce => \N__46107\,
            sr => \N__48129\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47061\,
            in1 => \N__43173\,
            in2 => \_gnd_net_\,
            in3 => \N__43157\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48783\,
            ce => \N__46107\,
            sr => \N__48129\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__38135\,
            in1 => \N__41351\,
            in2 => \N__38093\,
            in3 => \N__38113\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__41350\,
            in1 => \N__38134\,
            in2 => \N__38114\,
            in3 => \N__38092\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47058\,
            in1 => \N__43498\,
            in2 => \_gnd_net_\,
            in3 => \N__43473\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48771\,
            ce => \N__46108\,
            sr => \N__48133\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45004\,
            in1 => \N__44964\,
            in2 => \_gnd_net_\,
            in3 => \N__47060\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48771\,
            ce => \N__46108\,
            sr => \N__48133\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47059\,
            in1 => \N__44302\,
            in2 => \_gnd_net_\,
            in3 => \N__44253\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48771\,
            ce => \N__46108\,
            sr => \N__48133\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__38321\,
            in1 => \N__38296\,
            in2 => \N__41342\,
            in3 => \N__38606\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__38605\,
            in1 => \N__38320\,
            in2 => \N__38300\,
            in3 => \N__41338\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_27_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46935\,
            in1 => \N__43868\,
            in2 => \_gnd_net_\,
            in3 => \N__43824\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48763\,
            ce => \N__46111\,
            sr => \N__48139\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43472\,
            in1 => \N__43580\,
            in2 => \N__43559\,
            in3 => \N__43145\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38573\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48750\,
            ce => \N__44117\,
            sr => \N__48144\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38546\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48750\,
            ce => \N__44117\,
            sr => \N__48144\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43581\,
            in1 => \N__43618\,
            in2 => \_gnd_net_\,
            in3 => \N__46841\,
            lcout => \elapsed_time_ns_1_RNIED91B_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__38444\,
            in1 => \N__38453\,
            in2 => \N__38504\,
            in3 => \N__38484\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__38452\,
            in1 => \N__38502\,
            in2 => \N__38486\,
            in3 => \N__38443\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_20_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46932\,
            in1 => \N__43274\,
            in2 => \_gnd_net_\,
            in3 => \N__43245\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48739\,
            ce => \N__46114\,
            sr => \N__48154\
        );

    \phase_controller_inst2.stoper_tr.target_time_21_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42552\,
            in1 => \N__42487\,
            in2 => \_gnd_net_\,
            in3 => \N__46934\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48739\,
            ce => \N__46114\,
            sr => \N__48154\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42104\,
            in1 => \N__42116\,
            in2 => \_gnd_net_\,
            in3 => \N__46933\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48739\,
            ce => \N__46114\,
            sr => \N__48154\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__38385\,
            in1 => \N__38406\,
            in2 => \N__38645\,
            in3 => \N__38360\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__38359\,
            in1 => \N__38407\,
            in2 => \N__38390\,
            in3 => \N__38641\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_22_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47231\,
            in1 => \N__47209\,
            in2 => \_gnd_net_\,
            in3 => \N__47144\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48729\,
            ce => \N__46116\,
            sr => \N__48162\
        );

    \phase_controller_inst2.stoper_tr.target_time_23_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47348\,
            in1 => \N__47319\,
            in2 => \_gnd_net_\,
            in3 => \N__47110\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48729\,
            ce => \N__46116\,
            sr => \N__48162\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42071\,
            in1 => \N__42049\,
            in2 => \_gnd_net_\,
            in3 => \N__47141\,
            lcout => \elapsed_time_ns_1_RNIV8OBB_0_12\,
            ltout => \elapsed_time_ns_1_RNIV8OBB_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47111\,
            in2 => \N__38633\,
            in3 => \N__42072\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48729\,
            ce => \N__46116\,
            sr => \N__48162\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45996\,
            in1 => \N__45974\,
            in2 => \_gnd_net_\,
            in3 => \N__47143\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48729\,
            ce => \N__46116\,
            sr => \N__48162\
        );

    \phase_controller_inst2.stoper_tr.target_time_24_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47142\,
            in1 => \N__45540\,
            in2 => \_gnd_net_\,
            in3 => \N__45522\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48729\,
            ce => \N__46116\,
            sr => \N__48162\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42193\,
            in1 => \N__38591\,
            in2 => \_gnd_net_\,
            in3 => \N__47109\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48720\,
            ce => \N__46677\,
            sr => \N__48170\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47107\,
            in1 => \N__42169\,
            in2 => \_gnd_net_\,
            in3 => \N__42258\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48720\,
            ce => \N__46677\,
            sr => \N__48170\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47108\,
            in1 => \N__42216\,
            in2 => \_gnd_net_\,
            in3 => \N__42523\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48720\,
            ce => \N__46677\,
            sr => \N__48170\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38832\,
            in2 => \N__38569\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__48710\,
            ce => \N__44112\,
            sr => \N__48179\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38808\,
            in2 => \N__38542\,
            in3 => \N__38519\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__48710\,
            ce => \N__44112\,
            sr => \N__48179\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38784\,
            in2 => \N__38837\,
            in3 => \N__38816\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__48710\,
            ce => \N__44112\,
            sr => \N__48179\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38760\,
            in2 => \N__38813\,
            in3 => \N__38792\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__48710\,
            ce => \N__44112\,
            sr => \N__48179\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38736\,
            in2 => \N__38789\,
            in3 => \N__38768\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__48710\,
            ce => \N__44112\,
            sr => \N__48179\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38712\,
            in2 => \N__38765\,
            in3 => \N__38744\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__48710\,
            ce => \N__44112\,
            sr => \N__48179\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38688\,
            in2 => \N__38741\,
            in3 => \N__38720\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__48710\,
            ce => \N__44112\,
            sr => \N__48179\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38664\,
            in2 => \N__38717\,
            in3 => \N__38696\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__48710\,
            ce => \N__44112\,
            sr => \N__48179\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39021\,
            in2 => \N__38693\,
            in3 => \N__38672\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__48701\,
            ce => \N__44116\,
            sr => \N__48189\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39000\,
            in2 => \N__38669\,
            in3 => \N__38648\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__48701\,
            ce => \N__44116\,
            sr => \N__48189\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39022\,
            in2 => \N__38980\,
            in3 => \N__39008\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__48701\,
            ce => \N__44116\,
            sr => \N__48189\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38952\,
            in2 => \N__39005\,
            in3 => \N__38984\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__48701\,
            ce => \N__44116\,
            sr => \N__48189\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38928\,
            in2 => \N__38981\,
            in3 => \N__38960\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__48701\,
            ce => \N__44116\,
            sr => \N__48189\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38904\,
            in2 => \N__38957\,
            in3 => \N__38936\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__48701\,
            ce => \N__44116\,
            sr => \N__48189\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38880\,
            in2 => \N__38933\,
            in3 => \N__38912\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__48701\,
            ce => \N__44116\,
            sr => \N__48189\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38856\,
            in2 => \N__38909\,
            in3 => \N__38888\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__48701\,
            ce => \N__44116\,
            sr => \N__48189\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39243\,
            in2 => \N__38885\,
            in3 => \N__38864\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__48693\,
            ce => \N__44108\,
            sr => \N__48198\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39219\,
            in2 => \N__38861\,
            in3 => \N__38840\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__48693\,
            ce => \N__44108\,
            sr => \N__48198\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39195\,
            in2 => \N__39248\,
            in3 => \N__39227\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__48693\,
            ce => \N__44108\,
            sr => \N__48198\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39171\,
            in2 => \N__39224\,
            in3 => \N__39203\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__48693\,
            ce => \N__44108\,
            sr => \N__48198\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39147\,
            in2 => \N__39200\,
            in3 => \N__39179\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__48693\,
            ce => \N__44108\,
            sr => \N__48198\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39123\,
            in2 => \N__39176\,
            in3 => \N__39155\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__48693\,
            ce => \N__44108\,
            sr => \N__48198\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39099\,
            in2 => \N__39152\,
            in3 => \N__39131\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__48693\,
            ce => \N__44108\,
            sr => \N__48198\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39075\,
            in2 => \N__39128\,
            in3 => \N__39107\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__48693\,
            ce => \N__44108\,
            sr => \N__48198\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39054\,
            in2 => \N__39104\,
            in3 => \N__39083\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__48687\,
            ce => \N__44095\,
            sr => \N__48206\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39417\,
            in2 => \N__39080\,
            in3 => \N__39059\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__48687\,
            ce => \N__44095\,
            sr => \N__48206\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39055\,
            in2 => \N__39041\,
            in3 => \N__39026\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__48687\,
            ce => \N__44095\,
            sr => \N__48206\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39433\,
            in2 => \N__39422\,
            in3 => \N__39401\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__48687\,
            ce => \N__44095\,
            sr => \N__48206\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39398\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48687\,
            ce => \N__44095\,
            sr => \N__48206\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__43999\,
            in1 => \N__43964\,
            in2 => \_gnd_net_\,
            in3 => \N__44018\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48683\,
            ce => 'H',
            sr => \N__48213\
        );

    \phase_controller_inst1.start_timer_hc_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__42967\,
            in1 => \N__42668\,
            in2 => \N__42388\,
            in3 => \N__39395\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48683\,
            ce => 'H',
            sr => \N__48213\
        );

    \delay_measurement_inst.start_timer_tr_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43965\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42721\,
            ce => 'H',
            sr => \N__48219\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39388\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48674\,
            ce => 'H',
            sr => \N__48226\
        );

    \phase_controller_inst1.S1_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__39309\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48667\,
            ce => 'H',
            sr => \N__48230\
        );

    \current_shift_inst.start_timer_s1_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__39351\,
            in1 => \N__39308\,
            in2 => \_gnd_net_\,
            in3 => \N__39332\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48667\,
            ce => 'H',
            sr => \N__48230\
        );

    \phase_controller_inst1.T01_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39259\,
            in2 => \_gnd_net_\,
            in3 => \N__39310\,
            lcout => \T01_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48663\,
            ce => 'H',
            sr => \N__48235\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39892\,
            in2 => \N__39878\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39809\,
            in2 => \N__39800\,
            in3 => \N__39773\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__48660\,
            ce => 'H',
            sr => \N__48240\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39770\,
            in2 => \N__39758\,
            in3 => \N__39710\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__48660\,
            ce => 'H',
            sr => \N__48240\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39707\,
            in2 => \N__39695\,
            in3 => \N__39650\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__48660\,
            ce => 'H',
            sr => \N__48240\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39646\,
            in2 => \N__39605\,
            in3 => \N__39593\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__48660\,
            ce => 'H',
            sr => \N__48240\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39590\,
            in2 => \N__39580\,
            in3 => \N__39542\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__48660\,
            ce => 'H',
            sr => \N__48240\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39539\,
            in2 => \N__39530\,
            in3 => \N__39488\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__48660\,
            ce => 'H',
            sr => \N__48240\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39485\,
            in2 => \N__39476\,
            in3 => \N__39437\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__48660\,
            ce => 'H',
            sr => \N__48240\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40343\,
            in2 => \N__40334\,
            in3 => \N__40283\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_15_24_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__48657\,
            ce => 'H',
            sr => \N__48245\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40280\,
            in2 => \N__40271\,
            in3 => \N__40217\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__48657\,
            ce => 'H',
            sr => \N__48245\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40214\,
            in2 => \N__40202\,
            in3 => \N__40151\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__48657\,
            ce => 'H',
            sr => \N__48245\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40148\,
            in2 => \N__40136\,
            in3 => \N__40085\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__48657\,
            ce => 'H',
            sr => \N__48245\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40082\,
            in2 => \N__40043\,
            in3 => \N__40031\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__48657\,
            ce => 'H',
            sr => \N__48245\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40833\,
            in2 => \N__40028\,
            in3 => \N__39986\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__48657\,
            ce => 'H',
            sr => \N__48245\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39983\,
            in2 => \N__40867\,
            in3 => \N__39941\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__48657\,
            ce => 'H',
            sr => \N__48245\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40837\,
            in2 => \N__39938\,
            in3 => \N__39896\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__48657\,
            ce => 'H',
            sr => \N__48245\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40838\,
            in2 => \N__40736\,
            in3 => \N__40676\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_15_25_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__48654\,
            ce => 'H',
            sr => \N__48253\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40673\,
            in2 => \N__40868\,
            in3 => \N__40628\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__48654\,
            ce => 'H',
            sr => \N__48253\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40842\,
            in2 => \N__40625\,
            in3 => \N__40580\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__48654\,
            ce => 'H',
            sr => \N__48253\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40577\,
            in2 => \N__40869\,
            in3 => \N__40532\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__48654\,
            ce => 'H',
            sr => \N__48253\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40846\,
            in2 => \N__40528\,
            in3 => \N__40487\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__48654\,
            ce => 'H',
            sr => \N__48253\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40484\,
            in2 => \N__40870\,
            in3 => \N__40439\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__48654\,
            ce => 'H',
            sr => \N__48253\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40850\,
            in2 => \N__40436\,
            in3 => \N__40391\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__48654\,
            ce => 'H',
            sr => \N__48253\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40388\,
            in2 => \N__40871\,
            in3 => \N__40346\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__48654\,
            ce => 'H',
            sr => \N__48253\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40854\,
            in2 => \N__41315\,
            in3 => \N__41273\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_15_26_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__48651\,
            ce => 'H',
            sr => \N__48260\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41269\,
            in2 => \N__40872\,
            in3 => \N__41234\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__48651\,
            ce => 'H',
            sr => \N__48260\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40858\,
            in2 => \N__41231\,
            in3 => \N__41183\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__48651\,
            ce => 'H',
            sr => \N__48260\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41180\,
            in2 => \N__40873\,
            in3 => \N__41144\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__48651\,
            ce => 'H',
            sr => \N__48260\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40862\,
            in2 => \N__41141\,
            in3 => \N__41099\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__48651\,
            ce => 'H',
            sr => \N__48260\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41096\,
            in2 => \N__40874\,
            in3 => \N__41054\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__48651\,
            ce => 'H',
            sr => \N__48260\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__41051\,
            in1 => \N__40866\,
            in2 => \_gnd_net_\,
            in3 => \N__40781\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48651\,
            ce => 'H',
            sr => \N__48260\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__40759\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40774\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__41371\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41386\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43317\,
            in1 => \N__43337\,
            in2 => \_gnd_net_\,
            in3 => \N__47056\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48789\,
            ce => \N__46109\,
            sr => \N__48123\
        );

    \phase_controller_inst2.stoper_tr.target_time_25_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47055\,
            in1 => \N__45072\,
            in2 => \_gnd_net_\,
            in3 => \N__45056\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48789\,
            ce => \N__46109\,
            sr => \N__48123\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43520\,
            in1 => \N__43565\,
            in2 => \_gnd_net_\,
            in3 => \N__47057\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48789\,
            ce => \N__46109\,
            sr => \N__48123\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43177\,
            in1 => \N__43155\,
            in2 => \_gnd_net_\,
            in3 => \N__47052\,
            lcout => \elapsed_time_ns_1_RNIDC91B_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__44056\,
            in1 => \N__42907\,
            in2 => \_gnd_net_\,
            in3 => \N__46228\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47054\,
            in1 => \N__44298\,
            in2 => \_gnd_net_\,
            in3 => \N__44257\,
            lcout => \elapsed_time_ns_1_RNIIH91B_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44941\,
            in1 => \N__44919\,
            in2 => \_gnd_net_\,
            in3 => \N__47051\,
            lcout => \elapsed_time_ns_1_RNIKJ91B_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47053\,
            in1 => \N__43272\,
            in2 => \_gnd_net_\,
            in3 => \N__43249\,
            lcout => \elapsed_time_ns_1_RNIU8PBB_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43519\,
            in1 => \N__43560\,
            in2 => \_gnd_net_\,
            in3 => \N__46927\,
            lcout => \elapsed_time_ns_1_RNIFE91B_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__42025\,
            in1 => \N__41972\,
            in2 => \N__42005\,
            in3 => \N__46130\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43874\,
            in1 => \N__43828\,
            in2 => \_gnd_net_\,
            in3 => \N__46926\,
            lcout => \elapsed_time_ns_1_RNI5GPBB_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46928\,
            in1 => \N__45003\,
            in2 => \_gnd_net_\,
            in3 => \N__44965\,
            lcout => \elapsed_time_ns_1_RNIHG91B_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__46129\,
            in1 => \N__42026\,
            in2 => \N__42004\,
            in3 => \N__41971\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46925\,
            in1 => \N__44877\,
            in2 => \_gnd_net_\,
            in3 => \N__44854\,
            lcout => \elapsed_time_ns_1_RNIJI91B_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43499\,
            in1 => \N__43480\,
            in2 => \_gnd_net_\,
            in3 => \N__46929\,
            lcout => \elapsed_time_ns_1_RNIGF91B_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__43869\,
            in1 => \N__44231\,
            in2 => \_gnd_net_\,
            in3 => \N__41951\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41415\,
            in1 => \N__41944\,
            in2 => \_gnd_net_\,
            in3 => \N__41888\,
            lcout => \elapsed_time_ns_1_RNIV1DN9_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44915\,
            in2 => \_gnd_net_\,
            in3 => \N__44849\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__42122\,
            in1 => \N__44297\,
            in2 => \N__42137\,
            in3 => \N__45002\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__46394\,
            in1 => \N__42566\,
            in2 => \N__42134\,
            in3 => \N__42131\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__43405\,
            in1 => \_gnd_net_\,
            in2 => \N__42125\,
            in3 => \N__43384\,
            lcout => \elapsed_time_ns_1_RNI2COBB_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45976\,
            in1 => \N__42101\,
            in2 => \N__42077\,
            in3 => \N__44345\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46930\,
            in1 => \N__42115\,
            in2 => \_gnd_net_\,
            in3 => \N__42102\,
            lcout => \elapsed_time_ns_1_RNIT6OBB_0_10\,
            ltout => \elapsed_time_ns_1_RNIT6OBB_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__42103\,
            in1 => \_gnd_net_\,
            in2 => \N__42080\,
            in3 => \N__46931\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48751\,
            ce => \N__46699\,
            sr => \N__48145\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46936\,
            in1 => \N__42076\,
            in2 => \_gnd_net_\,
            in3 => \N__42050\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48751\,
            ce => \N__46699\,
            sr => \N__48145\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46975\,
            in1 => \N__45550\,
            in2 => \_gnd_net_\,
            in3 => \N__45523\,
            lcout => \elapsed_time_ns_1_RNI2DPBB_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46974\,
            in1 => \N__42553\,
            in2 => \_gnd_net_\,
            in3 => \N__42488\,
            lcout => \elapsed_time_ns_1_RNIV9PBB_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100111011"
        )
    port map (
            in0 => \N__45829\,
            in1 => \N__46246\,
            in2 => \N__45695\,
            in3 => \N__45632\,
            lcout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42287\,
            in3 => \N__46190\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46976\,
            in1 => \N__46000\,
            in2 => \_gnd_net_\,
            in3 => \N__45975\,
            lcout => \elapsed_time_ns_1_RNIU7OBB_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46191\,
            in2 => \_gnd_net_\,
            in3 => \N__42277\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000010"
        )
    port map (
            in0 => \N__42242\,
            in1 => \N__43789\,
            in2 => \N__43772\,
            in3 => \N__42233\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47083\,
            in1 => \N__42262\,
            in2 => \_gnd_net_\,
            in3 => \N__42165\,
            lcout => \elapsed_time_ns_1_RNI3DOBB_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__42241\,
            in1 => \N__43788\,
            in2 => \N__43771\,
            in3 => \N__42232\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47084\,
            in1 => \N__42220\,
            in2 => \_gnd_net_\,
            in3 => \N__42522\,
            lcout => \elapsed_time_ns_1_RNI4EOBB_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42192\,
            in1 => \N__43358\,
            in2 => \N__42164\,
            in3 => \N__46319\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__42533\,
            in1 => \N__42455\,
            in2 => \N__42569\,
            in3 => \N__42494\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_21_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42554\,
            in1 => \N__42486\,
            in2 => \_gnd_net_\,
            in3 => \N__47082\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48721\,
            ce => \N__46614\,
            sr => \N__48171\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__42418\,
            in1 => \_gnd_net_\,
            in2 => \N__47145\,
            in3 => \N__42445\,
            lcout => \elapsed_time_ns_1_RNI7IPBB_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45029\,
            in1 => \N__42417\,
            in2 => \N__45785\,
            in3 => \N__46044\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44766\,
            in1 => \N__43299\,
            in2 => \N__43232\,
            in3 => \N__42512\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47298\,
            in1 => \N__45507\,
            in2 => \N__47195\,
            in3 => \N__42473\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_29_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47081\,
            in1 => \N__42441\,
            in2 => \_gnd_net_\,
            in3 => \N__42413\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48702\,
            ce => \N__46676\,
            sr => \N__48190\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42384\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48694\,
            ce => 'H',
            sr => \N__48199\
        );

    \phase_controller_inst1.start_timer_tr_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__42962\,
            in1 => \N__42677\,
            in2 => \N__44055\,
            in3 => \N__44563\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48694\,
            ce => 'H',
            sr => \N__48199\
        );

    \delay_measurement_inst.stop_timer_tr_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43966\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42722\,
            ce => 'H',
            sr => \N__48207\
        );

    \phase_controller_inst1.state_RNIE87F_2_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__44627\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42709\,
            lcout => \phase_controller_inst1.state_RNIE87FZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__42633\,
            in1 => \N__42708\,
            in2 => \N__44632\,
            in3 => \N__43057\,
            lcout => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_1_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__42634\,
            in1 => \N__43067\,
            in2 => \_gnd_net_\,
            in3 => \N__42667\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48678\,
            ce => 'H',
            sr => \N__48220\
        );

    \phase_controller_inst1.T45_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42652\,
            in2 => \_gnd_net_\,
            in3 => \N__44578\,
            lcout => \T45_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48668\,
            ce => 'H',
            sr => \N__48231\
        );

    \phase_controller_inst1.state_0_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__46163\,
            in1 => \N__44579\,
            in2 => \N__42641\,
            in3 => \N__43069\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48668\,
            ce => 'H',
            sr => \N__48231\
        );

    \phase_controller_inst1.T23_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42586\,
            in2 => \_gnd_net_\,
            in3 => \N__43068\,
            lcout => \T23_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48664\,
            ce => 'H',
            sr => \N__48236\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42869\,
            in1 => \N__42575\,
            in2 => \N__43103\,
            in3 => \N__42881\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42824\,
            in1 => \N__42860\,
            in2 => \N__42812\,
            in3 => \N__42851\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42890\,
            in1 => \N__42842\,
            in2 => \N__42797\,
            in3 => \N__42833\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42889\,
            in2 => \_gnd_net_\,
            in3 => \N__42880\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__42773\,
            in1 => \N__42779\,
            in2 => \N__42872\,
            in3 => \N__42868\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44455\,
            in1 => \N__42859\,
            in2 => \N__44476\,
            in3 => \N__42850\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42841\,
            in2 => \_gnd_net_\,
            in3 => \N__42832\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__42823\,
            in1 => \N__42808\,
            in2 => \N__42755\,
            in3 => \N__42790\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__42740\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42730\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42772\,
            in1 => \N__43093\,
            in2 => \N__42758\,
            in3 => \N__42754\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__42739\,
            in1 => \N__43123\,
            in2 => \N__43115\,
            in3 => \N__42731\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__43124\,
            in1 => \N__43111\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_16_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44491\,
            in1 => \N__44509\,
            in2 => \N__43094\,
            in3 => \N__43079\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S2_LC_16_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43073\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48647\,
            ce => 'H',
            sr => \N__48272\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45076\,
            in1 => \N__45048\,
            in2 => \_gnd_net_\,
            in3 => \N__47065\,
            lcout => \elapsed_time_ns_1_RNI3EPBB_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47066\,
            in1 => \N__44371\,
            in2 => \_gnd_net_\,
            in3 => \N__44349\,
            lcout => \elapsed_time_ns_1_RNILK91B_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44057\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48790\,
            ce => 'H',
            sr => \N__48124\
        );

    \phase_controller_inst1.state_4_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42999\,
            in2 => \_gnd_net_\,
            in3 => \N__42929\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48790\,
            ce => 'H',
            sr => \N__48124\
        );

    \phase_controller_inst1.stoper_tr.running_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111110000"
        )
    port map (
            in0 => \N__46238\,
            in1 => \N__46271\,
            in2 => \N__42908\,
            in3 => \N__46189\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48790\,
            ce => 'H',
            sr => \N__48124\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__43747\,
            in1 => \N__43723\,
            in2 => \N__44750\,
            in3 => \N__43283\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__43282\,
            in1 => \N__43748\,
            in2 => \N__43727\,
            in3 => \N__44746\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44809\,
            in1 => \N__44788\,
            in2 => \_gnd_net_\,
            in3 => \N__46921\,
            lcout => \elapsed_time_ns_1_RNI6GOBB_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43401\,
            in1 => \N__43385\,
            in2 => \_gnd_net_\,
            in3 => \N__46924\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48784\,
            ce => \N__46706\,
            sr => \N__48130\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43318\,
            in1 => \N__43333\,
            in2 => \_gnd_net_\,
            in3 => \N__46922\,
            lcout => \elapsed_time_ns_1_RNI5FOBB_0_18\,
            ltout => \elapsed_time_ns_1_RNI5FOBB_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46923\,
            in1 => \_gnd_net_\,
            in2 => \N__43322\,
            in3 => \N__43319\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48784\,
            ce => \N__46706\,
            sr => \N__48130\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__43703\,
            in1 => \N__43192\,
            in2 => \N__43682\,
            in3 => \N__43205\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_20_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43273\,
            in1 => \N__43250\,
            in2 => \_gnd_net_\,
            in3 => \N__46993\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48772\,
            ce => \N__46675\,
            sr => \N__48134\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__43204\,
            in1 => \N__43681\,
            in2 => \N__43196\,
            in3 => \N__43702\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43178\,
            in1 => \N__43156\,
            in2 => \_gnd_net_\,
            in3 => \N__46992\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48772\,
            ce => \N__46675\,
            sr => \N__48134\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46990\,
            in1 => \N__43617\,
            in2 => \_gnd_net_\,
            in3 => \N__43588\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48772\,
            ce => \N__46675\,
            sr => \N__48134\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43564\,
            in1 => \N__43518\,
            in2 => \_gnd_net_\,
            in3 => \N__46994\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48772\,
            ce => \N__46675\,
            sr => \N__48134\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46991\,
            in1 => \N__43497\,
            in2 => \_gnd_net_\,
            in3 => \N__43481\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48772\,
            ce => \N__46675\,
            sr => \N__48134\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43442\,
            in2 => \N__44738\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46694\,
            in1 => \N__44687\,
            in2 => \_gnd_net_\,
            in3 => \N__43436\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__48764\,
            ce => 'H',
            sr => \N__48140\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__46601\,
            in1 => \N__44651\,
            in2 => \N__43433\,
            in3 => \N__43421\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__48764\,
            ce => 'H',
            sr => \N__48140\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46695\,
            in1 => \N__45284\,
            in2 => \_gnd_net_\,
            in3 => \N__43418\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__48764\,
            ce => 'H',
            sr => \N__48140\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46602\,
            in1 => \N__45266\,
            in2 => \_gnd_net_\,
            in3 => \N__43415\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__48764\,
            ce => 'H',
            sr => \N__48140\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46696\,
            in1 => \N__45230\,
            in2 => \_gnd_net_\,
            in3 => \N__43412\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__48764\,
            ce => 'H',
            sr => \N__48140\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46603\,
            in1 => \N__45203\,
            in2 => \_gnd_net_\,
            in3 => \N__43649\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__48764\,
            ce => 'H',
            sr => \N__48140\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46697\,
            in1 => \N__45176\,
            in2 => \_gnd_net_\,
            in3 => \N__43646\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__48764\,
            ce => 'H',
            sr => \N__48140\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46594\,
            in1 => \N__45145\,
            in2 => \_gnd_net_\,
            in3 => \N__43643\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__48752\,
            ce => 'H',
            sr => \N__48146\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46604\,
            in1 => \N__45122\,
            in2 => \_gnd_net_\,
            in3 => \N__43640\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__48752\,
            ce => 'H',
            sr => \N__48146\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46591\,
            in1 => \N__45089\,
            in2 => \_gnd_net_\,
            in3 => \N__43637\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__48752\,
            ce => 'H',
            sr => \N__48146\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46605\,
            in1 => \N__45476\,
            in2 => \_gnd_net_\,
            in3 => \N__43634\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__48752\,
            ce => 'H',
            sr => \N__48146\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46592\,
            in1 => \N__45455\,
            in2 => \_gnd_net_\,
            in3 => \N__43631\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__48752\,
            ce => 'H',
            sr => \N__48146\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46606\,
            in1 => \N__45422\,
            in2 => \_gnd_net_\,
            in3 => \N__43628\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__48752\,
            ce => 'H',
            sr => \N__48146\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46593\,
            in1 => \N__45392\,
            in2 => \_gnd_net_\,
            in3 => \N__43625\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__48752\,
            ce => 'H',
            sr => \N__48146\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46607\,
            in1 => \N__43790\,
            in2 => \_gnd_net_\,
            in3 => \N__43775\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__48752\,
            ce => 'H',
            sr => \N__48146\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46678\,
            in1 => \N__43770\,
            in2 => \_gnd_net_\,
            in3 => \N__43751\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__48740\,
            ce => 'H',
            sr => \N__48155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46682\,
            in1 => \N__43746\,
            in2 => \_gnd_net_\,
            in3 => \N__43730\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__48740\,
            ce => 'H',
            sr => \N__48155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46679\,
            in1 => \N__43722\,
            in2 => \_gnd_net_\,
            in3 => \N__43706\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__48740\,
            ce => 'H',
            sr => \N__48155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46683\,
            in1 => \N__43701\,
            in2 => \_gnd_net_\,
            in3 => \N__43685\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__48740\,
            ce => 'H',
            sr => \N__48155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46680\,
            in1 => \N__43677\,
            in2 => \_gnd_net_\,
            in3 => \N__43661\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__48740\,
            ce => 'H',
            sr => \N__48155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46684\,
            in1 => \N__47395\,
            in2 => \_gnd_net_\,
            in3 => \N__43658\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__48740\,
            ce => 'H',
            sr => \N__48155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46681\,
            in1 => \N__47371\,
            in2 => \_gnd_net_\,
            in3 => \N__43655\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__48740\,
            ce => 'H',
            sr => \N__48155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46685\,
            in1 => \N__45578\,
            in2 => \_gnd_net_\,
            in3 => \N__43652\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__48740\,
            ce => 'H',
            sr => \N__48155\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46661\,
            in1 => \N__45610\,
            in2 => \_gnd_net_\,
            in3 => \N__43895\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__48730\,
            ce => 'H',
            sr => \N__48163\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46608\,
            in1 => \N__45873\,
            in2 => \_gnd_net_\,
            in3 => \N__43892\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__48730\,
            ce => 'H',
            sr => \N__48163\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46662\,
            in1 => \N__45895\,
            in2 => \_gnd_net_\,
            in3 => \N__43889\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__48730\,
            ce => 'H',
            sr => \N__48163\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46609\,
            in1 => \N__44198\,
            in2 => \_gnd_net_\,
            in3 => \N__43886\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__48730\,
            ce => 'H',
            sr => \N__48163\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46663\,
            in1 => \N__44164\,
            in2 => \_gnd_net_\,
            in3 => \N__43883\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__48730\,
            ce => 'H',
            sr => \N__48163\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46610\,
            in1 => \N__45713\,
            in2 => \_gnd_net_\,
            in3 => \N__43880\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__48730\,
            ce => 'H',
            sr => \N__48163\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46664\,
            in1 => \N__45733\,
            in2 => \_gnd_net_\,
            in3 => \N__43877\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48730\,
            ce => 'H',
            sr => \N__48163\
        );

    \phase_controller_inst1.stoper_tr.target_time_27_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47089\,
            in1 => \N__43873\,
            in2 => \_gnd_net_\,
            in3 => \N__43832\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48722\,
            ce => \N__46657\,
            sr => \N__48172\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44233\,
            in1 => \N__43801\,
            in2 => \_gnd_net_\,
            in3 => \N__47088\,
            lcout => \elapsed_time_ns_1_RNI6HPBB_0_28\,
            ltout => \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_28_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__47090\,
            in1 => \_gnd_net_\,
            in2 => \N__44237\,
            in3 => \N__44234\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48722\,
            ce => \N__46657\,
            sr => \N__48172\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__44146\,
            in1 => \N__44163\,
            in2 => \N__44183\,
            in3 => \N__44197\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__44196\,
            in1 => \N__44179\,
            in2 => \N__44165\,
            in3 => \N__44147\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__45911\,
            in1 => \N__45891\,
            in2 => \N__45874\,
            in3 => \N__45850\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_31_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46396\,
            in1 => \N__46354\,
            in2 => \_gnd_net_\,
            in3 => \N__47106\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48711\,
            ce => \N__46118\,
            sr => \N__48180\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44000\,
            in2 => \_gnd_net_\,
            in3 => \N__44016\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_200_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46242\,
            in2 => \_gnd_net_\,
            in3 => \N__44042\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__44017\,
            in1 => \N__43995\,
            in2 => \_gnd_net_\,
            in3 => \N__43970\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_201_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.T12_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44590\,
            in2 => \_gnd_net_\,
            in3 => \N__44633\,
            lcout => \T12_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48688\,
            ce => 'H',
            sr => \N__48208\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46159\,
            in2 => \_gnd_net_\,
            in3 => \N__44577\,
            lcout => \phase_controller_inst1.state_RNI7NN7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44543\,
            in1 => \N__44537\,
            in2 => \N__44531\,
            in3 => \N__44522\,
            lcout => \current_shift_inst.PI_CTRL.N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_17_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44516\,
            in1 => \N__44498\,
            in2 => \N__44480\,
            in3 => \N__44459\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_17_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44444\,
            in1 => \N__44438\,
            in2 => \N__44432\,
            in3 => \N__44429\,
            lcout => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_17_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44419\,
            in2 => \_gnd_net_\,
            in3 => \N__44394\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44367\,
            in1 => \N__44351\,
            in2 => \_gnd_net_\,
            in3 => \N__47138\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48802\,
            ce => \N__46702\,
            sr => \N__48121\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44303\,
            in1 => \N__44258\,
            in2 => \_gnd_net_\,
            in3 => \N__47137\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48798\,
            ce => \N__46698\,
            sr => \N__48122\
        );

    \phase_controller_inst1.stoper_tr.target_time_25_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45077\,
            in1 => \N__45055\,
            in2 => \_gnd_net_\,
            in3 => \N__47135\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48791\,
            ce => \N__46687\,
            sr => \N__48125\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47132\,
            in1 => \N__45008\,
            in2 => \_gnd_net_\,
            in3 => \N__44966\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48791\,
            ce => \N__46687\,
            sr => \N__48125\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44945\,
            in1 => \N__44921\,
            in2 => \_gnd_net_\,
            in3 => \N__47136\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48791\,
            ce => \N__46687\,
            sr => \N__48125\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47133\,
            in1 => \N__44878\,
            in2 => \_gnd_net_\,
            in3 => \N__44855\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48791\,
            ce => \N__46687\,
            sr => \N__48125\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44805\,
            in1 => \N__44789\,
            in2 => \_gnd_net_\,
            in3 => \N__47134\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48791\,
            ce => \N__46687\,
            sr => \N__48125\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44734\,
            in1 => \N__44702\,
            in2 => \N__44696\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_18_10_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44686\,
            in1 => \N__44666\,
            in2 => \N__44675\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44639\,
            in2 => \N__44660\,
            in3 => \N__44650\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45272\,
            in2 => \N__45293\,
            in3 => \N__45283\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45265\,
            in1 => \N__45245\,
            in2 => \N__45254\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45239\,
            in2 => \N__45218\,
            in3 => \N__45229\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45209\,
            in2 => \N__45191\,
            in3 => \N__45202\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45182\,
            in2 => \N__45164\,
            in3 => \N__45175\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45155\,
            in2 => \N__45131\,
            in3 => \N__45146\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_18_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45121\,
            in1 => \N__45110\,
            in2 => \N__45101\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45491\,
            in2 => \N__45944\,
            in3 => \N__45088\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45485\,
            in2 => \N__45464\,
            in3 => \N__45475\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45454\,
            in1 => \N__45443\,
            in2 => \N__45431\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45680\,
            in2 => \N__45410\,
            in3 => \N__45421\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45401\,
            in2 => \N__45380\,
            in3 => \N__45391\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45368\,
            in2 => \N__45356\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45341\,
            in2 => \N__45329\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45314\,
            in2 => \N__45305\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47357\,
            in2 => \N__45932\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45617\,
            in2 => \N__45563\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45836\,
            in2 => \N__45671\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45656\,
            in2 => \N__45647\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45755\,
            in2 => \N__45830\,
            in3 => \N__45623\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45620\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100000100"
        )
    port map (
            in0 => \N__45577\,
            in1 => \N__45920\,
            in2 => \N__45611\,
            in3 => \N__45592\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__45919\,
            in1 => \N__45606\,
            in2 => \N__45593\,
            in3 => \N__45576\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_24_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47130\,
            in1 => \N__45551\,
            in2 => \_gnd_net_\,
            in3 => \N__45527\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48753\,
            ce => \N__46665\,
            sr => \N__48147\
        );

    \phase_controller_inst1.stoper_tr.target_time_26_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46028\,
            in1 => \N__46068\,
            in2 => \_gnd_net_\,
            in3 => \N__47131\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48753\,
            ce => \N__46665\,
            sr => \N__48147\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__45907\,
            in1 => \N__45896\,
            in2 => \N__45875\,
            in3 => \N__45851\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__45745\,
            in1 => \N__45728\,
            in2 => \N__46414\,
            in3 => \N__45711\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45786\,
            in1 => \N__45802\,
            in2 => \_gnd_net_\,
            in3 => \N__47123\,
            lcout => \elapsed_time_ns_1_RNIVAQBB_0_30\,
            ltout => \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_30_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__47124\,
            in1 => \_gnd_net_\,
            in2 => \N__45791\,
            in3 => \N__45787\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48741\,
            ce => \N__46615\,
            sr => \N__48156\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001101110001"
        )
    port map (
            in0 => \N__45712\,
            in1 => \N__46413\,
            in2 => \N__45734\,
            in3 => \N__45746\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__45744\,
            in1 => \N__45729\,
            in2 => \N__46415\,
            in3 => \N__45710\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46287\,
            in1 => \N__46335\,
            in2 => \_gnd_net_\,
            in3 => \N__47161\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48731\,
            ce => \N__46589\,
            sr => \N__48164\
        );

    \phase_controller_inst1.stoper_tr.target_time_31_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47160\,
            in1 => \N__46397\,
            in2 => \_gnd_net_\,
            in3 => \N__46353\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48731\,
            ce => \N__46589\,
            sr => \N__48164\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46355\,
            in1 => \N__46395\,
            in2 => \_gnd_net_\,
            in3 => \N__47140\,
            lcout => \elapsed_time_ns_1_RNI0CQBB_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47139\,
            in1 => \N__46291\,
            in2 => \_gnd_net_\,
            in3 => \N__46336\,
            lcout => \elapsed_time_ns_1_RNI1BOBB_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011001100"
        )
    port map (
            in0 => \N__46267\,
            in1 => \N__46149\,
            in2 => \N__46253\,
            in3 => \N__46201\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48712\,
            ce => 'H',
            sr => \N__48181\
        );

    \phase_controller_inst2.stoper_tr.target_time_26_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47163\,
            in1 => \N__46020\,
            in2 => \_gnd_net_\,
            in3 => \N__46076\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48803\,
            ce => \N__46117\,
            sr => \N__48126\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46024\,
            in1 => \N__46075\,
            in2 => \_gnd_net_\,
            in3 => \N__46977\,
            lcout => \elapsed_time_ns_1_RNI4FPBB_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47162\,
            in1 => \N__46004\,
            in2 => \_gnd_net_\,
            in3 => \N__45980\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48792\,
            ce => \N__46700\,
            sr => \N__48135\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__47282\,
            in1 => \N__46715\,
            in2 => \N__47405\,
            in3 => \N__47380\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_20_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__46714\,
            in1 => \N__47404\,
            in2 => \N__47381\,
            in3 => \N__47281\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47346\,
            in1 => \N__47323\,
            in2 => \_gnd_net_\,
            in3 => \N__47147\,
            lcout => \elapsed_time_ns_1_RNI1CPBB_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47205\,
            in1 => \N__47230\,
            in2 => \_gnd_net_\,
            in3 => \N__47146\,
            lcout => \elapsed_time_ns_1_RNI0BPBB_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_23_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47347\,
            in1 => \N__47324\,
            in2 => \_gnd_net_\,
            in3 => \N__47165\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48754\,
            ce => \N__46590\,
            sr => \N__48165\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47270\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48713\,
            ce => 'H',
            sr => \N__48200\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47240\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48695\,
            ce => 'H',
            sr => \N__48214\
        );

    \phase_controller_inst1.stoper_tr.target_time_22_LC_21_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47226\,
            in1 => \N__47210\,
            in2 => \_gnd_net_\,
            in3 => \N__47164\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48793\,
            ce => \N__46686\,
            sr => \N__48148\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_22_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__49177\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47691\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_22_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48900\,
            in2 => \_gnd_net_\,
            in3 => \N__49176\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_22_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101011"
        )
    port map (
            in0 => \N__47411\,
            in1 => \N__47573\,
            in2 => \N__49094\,
            in3 => \N__47780\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49234\,
            in1 => \N__47501\,
            in2 => \N__48907\,
            in3 => \N__47758\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => \current_shift_inst.PI_CTRL.N_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_22_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__48962\,
            in1 => \N__47486\,
            in2 => \N__47495\,
            in3 => \N__48851\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_22_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__49233\,
            in1 => \N__47757\,
            in2 => \N__47705\,
            in3 => \N__47492\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_22_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49116\,
            in2 => \_gnd_net_\,
            in3 => \N__47605\,
            lcout => \current_shift_inst.PI_CTRL.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_23_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101110"
        )
    port map (
            in0 => \N__49300\,
            in1 => \N__47620\,
            in2 => \N__49066\,
            in3 => \N__47609\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_23_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47665\,
            in1 => \N__48827\,
            in2 => \N__49208\,
            in3 => \N__47722\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_23_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__49160\,
            in1 => \N__47572\,
            in2 => \N__47480\,
            in3 => \N__49087\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_23_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47721\,
            in2 => \_gnd_net_\,
            in3 => \N__49159\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_23_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__48826\,
            in1 => \N__47664\,
            in2 => \N__47414\,
            in3 => \N__49203\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_23_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__47635\,
            in1 => \N__49345\,
            in2 => \_gnd_net_\,
            in3 => \N__49252\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_23_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__48959\,
            in1 => \N__49125\,
            in2 => \_gnd_net_\,
            in3 => \N__47772\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_23_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__48961\,
            in1 => \N__47774\,
            in2 => \N__49065\,
            in3 => \N__49126\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_23_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__47773\,
            in1 => \N__49050\,
            in2 => \_gnd_net_\,
            in3 => \N__48960\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001010100"
        )
    port map (
            in0 => \N__48980\,
            in1 => \N__49062\,
            in2 => \N__47762\,
            in3 => \N__48872\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48723\,
            ce => 'H',
            sr => \N__48241\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001010100"
        )
    port map (
            in0 => \N__48979\,
            in1 => \N__49064\,
            in2 => \N__47704\,
            in3 => \N__48871\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48714\,
            ce => 'H',
            sr => \N__48246\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_24_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__49329\,
            in1 => \N__49317\,
            in2 => \N__49288\,
            in3 => \N__47648\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48714\,
            ce => 'H',
            sr => \N__48246\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_24_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101010001"
        )
    port map (
            in0 => \N__49316\,
            in1 => \N__47621\,
            in2 => \N__49067\,
            in3 => \N__47604\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48714\,
            ce => 'H',
            sr => \N__48246\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_24_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__49281\,
            in1 => \N__49361\,
            in2 => \N__49319\,
            in3 => \N__49330\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48714\,
            ce => 'H',
            sr => \N__48246\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_24_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__49331\,
            in1 => \N__49318\,
            in2 => \N__49289\,
            in3 => \N__49268\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48714\,
            ce => 'H',
            sr => \N__48246\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010001010100"
        )
    port map (
            in0 => \N__48978\,
            in1 => \N__49063\,
            in2 => \N__49238\,
            in3 => \N__48870\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48714\,
            ce => 'H',
            sr => \N__48246\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_24_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__49054\,
            in1 => \N__48976\,
            in2 => \N__49187\,
            in3 => \N__48867\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48703\,
            ce => 'H',
            sr => \N__48254\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_24_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__49145\,
            in1 => \N__49139\,
            in2 => \N__49130\,
            in3 => \N__48869\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48703\,
            ce => 'H',
            sr => \N__48254\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_24_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__49055\,
            in1 => \N__48977\,
            in2 => \N__48908\,
            in3 => \N__48868\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48703\,
            ce => 'H',
            sr => \N__48254\
        );
end \INTERFACE\;
