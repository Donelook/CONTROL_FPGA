// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 24 2025 22:19:58

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    start_stop,
    s2_phy,
    T23,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    T45,
    T12,
    s4_phy,
    rgb_g,
    T01,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    input start_stop;
    output s2_phy;
    output T23;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output T45;
    output T12;
    output s4_phy;
    output rgb_g;
    output T01;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__47639;
    wire N__47638;
    wire N__47637;
    wire N__47628;
    wire N__47627;
    wire N__47626;
    wire N__47619;
    wire N__47618;
    wire N__47617;
    wire N__47610;
    wire N__47609;
    wire N__47608;
    wire N__47601;
    wire N__47600;
    wire N__47599;
    wire N__47592;
    wire N__47591;
    wire N__47590;
    wire N__47583;
    wire N__47582;
    wire N__47581;
    wire N__47574;
    wire N__47573;
    wire N__47572;
    wire N__47565;
    wire N__47564;
    wire N__47563;
    wire N__47556;
    wire N__47555;
    wire N__47554;
    wire N__47547;
    wire N__47546;
    wire N__47545;
    wire N__47538;
    wire N__47537;
    wire N__47536;
    wire N__47529;
    wire N__47528;
    wire N__47527;
    wire N__47520;
    wire N__47519;
    wire N__47518;
    wire N__47511;
    wire N__47510;
    wire N__47509;
    wire N__47502;
    wire N__47501;
    wire N__47500;
    wire N__47493;
    wire N__47492;
    wire N__47491;
    wire N__47474;
    wire N__47471;
    wire N__47470;
    wire N__47467;
    wire N__47466;
    wire N__47463;
    wire N__47460;
    wire N__47457;
    wire N__47450;
    wire N__47449;
    wire N__47446;
    wire N__47443;
    wire N__47440;
    wire N__47439;
    wire N__47436;
    wire N__47433;
    wire N__47430;
    wire N__47429;
    wire N__47424;
    wire N__47421;
    wire N__47418;
    wire N__47411;
    wire N__47408;
    wire N__47405;
    wire N__47402;
    wire N__47399;
    wire N__47396;
    wire N__47393;
    wire N__47390;
    wire N__47387;
    wire N__47384;
    wire N__47381;
    wire N__47378;
    wire N__47375;
    wire N__47372;
    wire N__47369;
    wire N__47368;
    wire N__47367;
    wire N__47366;
    wire N__47365;
    wire N__47364;
    wire N__47363;
    wire N__47362;
    wire N__47361;
    wire N__47360;
    wire N__47359;
    wire N__47358;
    wire N__47357;
    wire N__47356;
    wire N__47355;
    wire N__47354;
    wire N__47353;
    wire N__47352;
    wire N__47351;
    wire N__47350;
    wire N__47347;
    wire N__47346;
    wire N__47345;
    wire N__47344;
    wire N__47343;
    wire N__47342;
    wire N__47341;
    wire N__47340;
    wire N__47339;
    wire N__47338;
    wire N__47337;
    wire N__47336;
    wire N__47335;
    wire N__47334;
    wire N__47333;
    wire N__47332;
    wire N__47329;
    wire N__47328;
    wire N__47327;
    wire N__47326;
    wire N__47325;
    wire N__47322;
    wire N__47311;
    wire N__47308;
    wire N__47299;
    wire N__47292;
    wire N__47289;
    wire N__47286;
    wire N__47281;
    wire N__47278;
    wire N__47265;
    wire N__47258;
    wire N__47257;
    wire N__47256;
    wire N__47253;
    wire N__47250;
    wire N__47241;
    wire N__47238;
    wire N__47229;
    wire N__47228;
    wire N__47227;
    wire N__47226;
    wire N__47225;
    wire N__47224;
    wire N__47223;
    wire N__47222;
    wire N__47221;
    wire N__47218;
    wire N__47215;
    wire N__47206;
    wire N__47205;
    wire N__47204;
    wire N__47203;
    wire N__47202;
    wire N__47201;
    wire N__47200;
    wire N__47199;
    wire N__47198;
    wire N__47197;
    wire N__47196;
    wire N__47195;
    wire N__47194;
    wire N__47193;
    wire N__47188;
    wire N__47181;
    wire N__47180;
    wire N__47179;
    wire N__47178;
    wire N__47177;
    wire N__47172;
    wire N__47169;
    wire N__47160;
    wire N__47143;
    wire N__47136;
    wire N__47119;
    wire N__47110;
    wire N__47109;
    wire N__47106;
    wire N__47105;
    wire N__47104;
    wire N__47103;
    wire N__47100;
    wire N__47097;
    wire N__47088;
    wire N__47085;
    wire N__47072;
    wire N__47061;
    wire N__47048;
    wire N__47047;
    wire N__47046;
    wire N__47043;
    wire N__47040;
    wire N__47037;
    wire N__47034;
    wire N__47031;
    wire N__47028;
    wire N__47027;
    wire N__47024;
    wire N__47021;
    wire N__47018;
    wire N__47015;
    wire N__47006;
    wire N__47005;
    wire N__47004;
    wire N__47003;
    wire N__47002;
    wire N__46999;
    wire N__46996;
    wire N__46993;
    wire N__46992;
    wire N__46989;
    wire N__46988;
    wire N__46987;
    wire N__46986;
    wire N__46985;
    wire N__46984;
    wire N__46983;
    wire N__46982;
    wire N__46981;
    wire N__46980;
    wire N__46977;
    wire N__46976;
    wire N__46975;
    wire N__46974;
    wire N__46973;
    wire N__46972;
    wire N__46971;
    wire N__46970;
    wire N__46969;
    wire N__46968;
    wire N__46967;
    wire N__46966;
    wire N__46965;
    wire N__46964;
    wire N__46963;
    wire N__46962;
    wire N__46961;
    wire N__46960;
    wire N__46959;
    wire N__46958;
    wire N__46957;
    wire N__46954;
    wire N__46951;
    wire N__46948;
    wire N__46943;
    wire N__46934;
    wire N__46927;
    wire N__46926;
    wire N__46923;
    wire N__46922;
    wire N__46919;
    wire N__46918;
    wire N__46917;
    wire N__46916;
    wire N__46915;
    wire N__46914;
    wire N__46913;
    wire N__46912;
    wire N__46911;
    wire N__46908;
    wire N__46899;
    wire N__46892;
    wire N__46887;
    wire N__46886;
    wire N__46885;
    wire N__46884;
    wire N__46883;
    wire N__46882;
    wire N__46881;
    wire N__46880;
    wire N__46879;
    wire N__46878;
    wire N__46877;
    wire N__46876;
    wire N__46875;
    wire N__46874;
    wire N__46873;
    wire N__46872;
    wire N__46871;
    wire N__46868;
    wire N__46867;
    wire N__46864;
    wire N__46863;
    wire N__46860;
    wire N__46859;
    wire N__46856;
    wire N__46855;
    wire N__46852;
    wire N__46851;
    wire N__46848;
    wire N__46847;
    wire N__46844;
    wire N__46843;
    wire N__46840;
    wire N__46839;
    wire N__46836;
    wire N__46835;
    wire N__46832;
    wire N__46831;
    wire N__46828;
    wire N__46827;
    wire N__46826;
    wire N__46825;
    wire N__46824;
    wire N__46819;
    wire N__46816;
    wire N__46813;
    wire N__46808;
    wire N__46807;
    wire N__46806;
    wire N__46805;
    wire N__46804;
    wire N__46803;
    wire N__46802;
    wire N__46801;
    wire N__46800;
    wire N__46789;
    wire N__46788;
    wire N__46785;
    wire N__46784;
    wire N__46781;
    wire N__46780;
    wire N__46777;
    wire N__46776;
    wire N__46773;
    wire N__46772;
    wire N__46769;
    wire N__46768;
    wire N__46765;
    wire N__46764;
    wire N__46761;
    wire N__46760;
    wire N__46759;
    wire N__46758;
    wire N__46757;
    wire N__46756;
    wire N__46751;
    wire N__46748;
    wire N__46745;
    wire N__46742;
    wire N__46725;
    wire N__46714;
    wire N__46697;
    wire N__46680;
    wire N__46663;
    wire N__46660;
    wire N__46659;
    wire N__46656;
    wire N__46655;
    wire N__46652;
    wire N__46651;
    wire N__46650;
    wire N__46649;
    wire N__46648;
    wire N__46645;
    wire N__46642;
    wire N__46637;
    wire N__46634;
    wire N__46633;
    wire N__46632;
    wire N__46629;
    wire N__46628;
    wire N__46625;
    wire N__46622;
    wire N__46619;
    wire N__46618;
    wire N__46617;
    wire N__46614;
    wire N__46613;
    wire N__46610;
    wire N__46607;
    wire N__46606;
    wire N__46605;
    wire N__46602;
    wire N__46587;
    wire N__46570;
    wire N__46567;
    wire N__46566;
    wire N__46563;
    wire N__46562;
    wire N__46559;
    wire N__46558;
    wire N__46555;
    wire N__46554;
    wire N__46543;
    wire N__46534;
    wire N__46521;
    wire N__46518;
    wire N__46517;
    wire N__46514;
    wire N__46513;
    wire N__46510;
    wire N__46509;
    wire N__46504;
    wire N__46501;
    wire N__46490;
    wire N__46483;
    wire N__46474;
    wire N__46469;
    wire N__46464;
    wire N__46457;
    wire N__46440;
    wire N__46433;
    wire N__46420;
    wire N__46397;
    wire N__46394;
    wire N__46393;
    wire N__46390;
    wire N__46389;
    wire N__46386;
    wire N__46383;
    wire N__46380;
    wire N__46377;
    wire N__46374;
    wire N__46371;
    wire N__46364;
    wire N__46361;
    wire N__46358;
    wire N__46355;
    wire N__46352;
    wire N__46351;
    wire N__46350;
    wire N__46347;
    wire N__46344;
    wire N__46341;
    wire N__46338;
    wire N__46335;
    wire N__46332;
    wire N__46329;
    wire N__46326;
    wire N__46323;
    wire N__46320;
    wire N__46317;
    wire N__46314;
    wire N__46311;
    wire N__46308;
    wire N__46305;
    wire N__46302;
    wire N__46299;
    wire N__46296;
    wire N__46293;
    wire N__46286;
    wire N__46285;
    wire N__46282;
    wire N__46279;
    wire N__46274;
    wire N__46273;
    wire N__46272;
    wire N__46269;
    wire N__46264;
    wire N__46261;
    wire N__46256;
    wire N__46253;
    wire N__46250;
    wire N__46247;
    wire N__46244;
    wire N__46243;
    wire N__46240;
    wire N__46237;
    wire N__46234;
    wire N__46233;
    wire N__46230;
    wire N__46229;
    wire N__46228;
    wire N__46225;
    wire N__46222;
    wire N__46221;
    wire N__46218;
    wire N__46215;
    wire N__46212;
    wire N__46207;
    wire N__46204;
    wire N__46201;
    wire N__46196;
    wire N__46193;
    wire N__46190;
    wire N__46187;
    wire N__46182;
    wire N__46175;
    wire N__46172;
    wire N__46169;
    wire N__46168;
    wire N__46165;
    wire N__46162;
    wire N__46159;
    wire N__46156;
    wire N__46153;
    wire N__46152;
    wire N__46151;
    wire N__46148;
    wire N__46145;
    wire N__46140;
    wire N__46133;
    wire N__46130;
    wire N__46129;
    wire N__46126;
    wire N__46123;
    wire N__46118;
    wire N__46117;
    wire N__46116;
    wire N__46115;
    wire N__46114;
    wire N__46113;
    wire N__46112;
    wire N__46111;
    wire N__46110;
    wire N__46109;
    wire N__46108;
    wire N__46107;
    wire N__46106;
    wire N__46105;
    wire N__46104;
    wire N__46103;
    wire N__46102;
    wire N__46101;
    wire N__46100;
    wire N__46099;
    wire N__46098;
    wire N__46097;
    wire N__46096;
    wire N__46095;
    wire N__46094;
    wire N__46093;
    wire N__46092;
    wire N__46091;
    wire N__46090;
    wire N__46089;
    wire N__46088;
    wire N__46087;
    wire N__46086;
    wire N__46085;
    wire N__46084;
    wire N__46083;
    wire N__46082;
    wire N__46081;
    wire N__46080;
    wire N__46079;
    wire N__46078;
    wire N__46077;
    wire N__46076;
    wire N__46075;
    wire N__46074;
    wire N__46073;
    wire N__46072;
    wire N__46071;
    wire N__46070;
    wire N__46069;
    wire N__46068;
    wire N__46067;
    wire N__46066;
    wire N__46065;
    wire N__46064;
    wire N__46063;
    wire N__46062;
    wire N__46061;
    wire N__46060;
    wire N__46059;
    wire N__46058;
    wire N__46057;
    wire N__46056;
    wire N__46055;
    wire N__46054;
    wire N__46053;
    wire N__46052;
    wire N__46051;
    wire N__46050;
    wire N__46049;
    wire N__46048;
    wire N__46047;
    wire N__46046;
    wire N__46045;
    wire N__46044;
    wire N__46043;
    wire N__46042;
    wire N__46041;
    wire N__46040;
    wire N__46039;
    wire N__46038;
    wire N__46037;
    wire N__46036;
    wire N__46035;
    wire N__46034;
    wire N__46033;
    wire N__46032;
    wire N__46031;
    wire N__46030;
    wire N__46029;
    wire N__46028;
    wire N__46027;
    wire N__46026;
    wire N__46025;
    wire N__46024;
    wire N__46023;
    wire N__46022;
    wire N__46021;
    wire N__46020;
    wire N__46019;
    wire N__46018;
    wire N__46017;
    wire N__46016;
    wire N__46015;
    wire N__46014;
    wire N__46013;
    wire N__46012;
    wire N__46011;
    wire N__46010;
    wire N__46009;
    wire N__46008;
    wire N__46007;
    wire N__46006;
    wire N__46005;
    wire N__46004;
    wire N__46003;
    wire N__46002;
    wire N__46001;
    wire N__46000;
    wire N__45999;
    wire N__45998;
    wire N__45997;
    wire N__45996;
    wire N__45995;
    wire N__45994;
    wire N__45993;
    wire N__45992;
    wire N__45991;
    wire N__45990;
    wire N__45731;
    wire N__45728;
    wire N__45727;
    wire N__45726;
    wire N__45725;
    wire N__45724;
    wire N__45723;
    wire N__45722;
    wire N__45721;
    wire N__45720;
    wire N__45719;
    wire N__45718;
    wire N__45717;
    wire N__45716;
    wire N__45715;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45705;
    wire N__45702;
    wire N__45699;
    wire N__45694;
    wire N__45691;
    wire N__45686;
    wire N__45683;
    wire N__45678;
    wire N__45675;
    wire N__45672;
    wire N__45669;
    wire N__45666;
    wire N__45663;
    wire N__45662;
    wire N__45659;
    wire N__45658;
    wire N__45657;
    wire N__45656;
    wire N__45655;
    wire N__45654;
    wire N__45653;
    wire N__45652;
    wire N__45651;
    wire N__45650;
    wire N__45649;
    wire N__45646;
    wire N__45643;
    wire N__45642;
    wire N__45641;
    wire N__45640;
    wire N__45639;
    wire N__45638;
    wire N__45637;
    wire N__45636;
    wire N__45635;
    wire N__45634;
    wire N__45633;
    wire N__45632;
    wire N__45631;
    wire N__45630;
    wire N__45627;
    wire N__45626;
    wire N__45625;
    wire N__45624;
    wire N__45623;
    wire N__45622;
    wire N__45621;
    wire N__45620;
    wire N__45619;
    wire N__45616;
    wire N__45613;
    wire N__45612;
    wire N__45611;
    wire N__45610;
    wire N__45609;
    wire N__45608;
    wire N__45607;
    wire N__45606;
    wire N__45605;
    wire N__45604;
    wire N__45603;
    wire N__45602;
    wire N__45601;
    wire N__45600;
    wire N__45599;
    wire N__45598;
    wire N__45597;
    wire N__45596;
    wire N__45595;
    wire N__45594;
    wire N__45593;
    wire N__45592;
    wire N__45591;
    wire N__45590;
    wire N__45589;
    wire N__45588;
    wire N__45587;
    wire N__45586;
    wire N__45585;
    wire N__45584;
    wire N__45583;
    wire N__45582;
    wire N__45581;
    wire N__45580;
    wire N__45579;
    wire N__45578;
    wire N__45577;
    wire N__45576;
    wire N__45575;
    wire N__45574;
    wire N__45573;
    wire N__45572;
    wire N__45571;
    wire N__45570;
    wire N__45569;
    wire N__45568;
    wire N__45567;
    wire N__45566;
    wire N__45565;
    wire N__45564;
    wire N__45563;
    wire N__45562;
    wire N__45561;
    wire N__45560;
    wire N__45559;
    wire N__45558;
    wire N__45557;
    wire N__45556;
    wire N__45555;
    wire N__45554;
    wire N__45553;
    wire N__45552;
    wire N__45551;
    wire N__45550;
    wire N__45549;
    wire N__45548;
    wire N__45547;
    wire N__45546;
    wire N__45545;
    wire N__45544;
    wire N__45543;
    wire N__45542;
    wire N__45541;
    wire N__45540;
    wire N__45539;
    wire N__45538;
    wire N__45537;
    wire N__45536;
    wire N__45535;
    wire N__45534;
    wire N__45533;
    wire N__45532;
    wire N__45531;
    wire N__45530;
    wire N__45529;
    wire N__45528;
    wire N__45527;
    wire N__45526;
    wire N__45523;
    wire N__45520;
    wire N__45519;
    wire N__45516;
    wire N__45515;
    wire N__45514;
    wire N__45245;
    wire N__45242;
    wire N__45239;
    wire N__45238;
    wire N__45235;
    wire N__45232;
    wire N__45229;
    wire N__45228;
    wire N__45225;
    wire N__45224;
    wire N__45221;
    wire N__45218;
    wire N__45215;
    wire N__45212;
    wire N__45209;
    wire N__45206;
    wire N__45201;
    wire N__45196;
    wire N__45191;
    wire N__45190;
    wire N__45187;
    wire N__45184;
    wire N__45183;
    wire N__45180;
    wire N__45177;
    wire N__45174;
    wire N__45167;
    wire N__45164;
    wire N__45161;
    wire N__45158;
    wire N__45155;
    wire N__45154;
    wire N__45151;
    wire N__45148;
    wire N__45145;
    wire N__45142;
    wire N__45141;
    wire N__45138;
    wire N__45135;
    wire N__45132;
    wire N__45131;
    wire N__45126;
    wire N__45123;
    wire N__45120;
    wire N__45113;
    wire N__45112;
    wire N__45109;
    wire N__45106;
    wire N__45105;
    wire N__45102;
    wire N__45099;
    wire N__45096;
    wire N__45089;
    wire N__45086;
    wire N__45083;
    wire N__45080;
    wire N__45079;
    wire N__45076;
    wire N__45075;
    wire N__45072;
    wire N__45069;
    wire N__45066;
    wire N__45061;
    wire N__45060;
    wire N__45057;
    wire N__45054;
    wire N__45051;
    wire N__45048;
    wire N__45041;
    wire N__45038;
    wire N__45037;
    wire N__45036;
    wire N__45033;
    wire N__45030;
    wire N__45027;
    wire N__45024;
    wire N__45021;
    wire N__45018;
    wire N__45015;
    wire N__45012;
    wire N__45005;
    wire N__45002;
    wire N__44999;
    wire N__44996;
    wire N__44993;
    wire N__44990;
    wire N__44987;
    wire N__44986;
    wire N__44983;
    wire N__44980;
    wire N__44979;
    wire N__44978;
    wire N__44975;
    wire N__44972;
    wire N__44969;
    wire N__44966;
    wire N__44957;
    wire N__44954;
    wire N__44953;
    wire N__44952;
    wire N__44949;
    wire N__44946;
    wire N__44943;
    wire N__44938;
    wire N__44935;
    wire N__44932;
    wire N__44927;
    wire N__44924;
    wire N__44921;
    wire N__44918;
    wire N__44917;
    wire N__44916;
    wire N__44915;
    wire N__44912;
    wire N__44905;
    wire N__44902;
    wire N__44899;
    wire N__44896;
    wire N__44893;
    wire N__44888;
    wire N__44885;
    wire N__44882;
    wire N__44879;
    wire N__44878;
    wire N__44877;
    wire N__44874;
    wire N__44869;
    wire N__44864;
    wire N__44861;
    wire N__44858;
    wire N__44857;
    wire N__44854;
    wire N__44851;
    wire N__44848;
    wire N__44845;
    wire N__44842;
    wire N__44841;
    wire N__44840;
    wire N__44837;
    wire N__44834;
    wire N__44831;
    wire N__44828;
    wire N__44819;
    wire N__44818;
    wire N__44815;
    wire N__44812;
    wire N__44811;
    wire N__44808;
    wire N__44805;
    wire N__44802;
    wire N__44797;
    wire N__44792;
    wire N__44789;
    wire N__44786;
    wire N__44783;
    wire N__44780;
    wire N__44777;
    wire N__44776;
    wire N__44775;
    wire N__44772;
    wire N__44769;
    wire N__44766;
    wire N__44763;
    wire N__44760;
    wire N__44757;
    wire N__44756;
    wire N__44753;
    wire N__44750;
    wire N__44747;
    wire N__44744;
    wire N__44735;
    wire N__44734;
    wire N__44733;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44719;
    wire N__44714;
    wire N__44711;
    wire N__44708;
    wire N__44705;
    wire N__44702;
    wire N__44699;
    wire N__44698;
    wire N__44697;
    wire N__44694;
    wire N__44691;
    wire N__44688;
    wire N__44681;
    wire N__44680;
    wire N__44679;
    wire N__44676;
    wire N__44673;
    wire N__44670;
    wire N__44667;
    wire N__44664;
    wire N__44663;
    wire N__44660;
    wire N__44655;
    wire N__44652;
    wire N__44645;
    wire N__44642;
    wire N__44639;
    wire N__44636;
    wire N__44633;
    wire N__44630;
    wire N__44627;
    wire N__44624;
    wire N__44621;
    wire N__44618;
    wire N__44615;
    wire N__44612;
    wire N__44609;
    wire N__44606;
    wire N__44603;
    wire N__44600;
    wire N__44597;
    wire N__44594;
    wire N__44591;
    wire N__44588;
    wire N__44585;
    wire N__44582;
    wire N__44579;
    wire N__44576;
    wire N__44573;
    wire N__44570;
    wire N__44567;
    wire N__44564;
    wire N__44561;
    wire N__44558;
    wire N__44555;
    wire N__44552;
    wire N__44549;
    wire N__44546;
    wire N__44543;
    wire N__44540;
    wire N__44539;
    wire N__44536;
    wire N__44533;
    wire N__44530;
    wire N__44527;
    wire N__44524;
    wire N__44519;
    wire N__44516;
    wire N__44513;
    wire N__44510;
    wire N__44507;
    wire N__44504;
    wire N__44501;
    wire N__44498;
    wire N__44495;
    wire N__44492;
    wire N__44489;
    wire N__44486;
    wire N__44483;
    wire N__44480;
    wire N__44477;
    wire N__44474;
    wire N__44471;
    wire N__44468;
    wire N__44465;
    wire N__44462;
    wire N__44459;
    wire N__44456;
    wire N__44453;
    wire N__44450;
    wire N__44447;
    wire N__44444;
    wire N__44441;
    wire N__44438;
    wire N__44435;
    wire N__44432;
    wire N__44429;
    wire N__44426;
    wire N__44423;
    wire N__44420;
    wire N__44417;
    wire N__44414;
    wire N__44411;
    wire N__44408;
    wire N__44405;
    wire N__44402;
    wire N__44399;
    wire N__44396;
    wire N__44393;
    wire N__44390;
    wire N__44387;
    wire N__44384;
    wire N__44381;
    wire N__44378;
    wire N__44375;
    wire N__44372;
    wire N__44369;
    wire N__44366;
    wire N__44363;
    wire N__44360;
    wire N__44357;
    wire N__44354;
    wire N__44351;
    wire N__44348;
    wire N__44345;
    wire N__44342;
    wire N__44339;
    wire N__44336;
    wire N__44333;
    wire N__44330;
    wire N__44327;
    wire N__44324;
    wire N__44321;
    wire N__44318;
    wire N__44315;
    wire N__44312;
    wire N__44309;
    wire N__44306;
    wire N__44303;
    wire N__44300;
    wire N__44297;
    wire N__44294;
    wire N__44293;
    wire N__44292;
    wire N__44291;
    wire N__44290;
    wire N__44289;
    wire N__44286;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44274;
    wire N__44273;
    wire N__44272;
    wire N__44271;
    wire N__44270;
    wire N__44269;
    wire N__44268;
    wire N__44267;
    wire N__44266;
    wire N__44265;
    wire N__44264;
    wire N__44263;
    wire N__44262;
    wire N__44261;
    wire N__44260;
    wire N__44259;
    wire N__44258;
    wire N__44257;
    wire N__44256;
    wire N__44253;
    wire N__44250;
    wire N__44247;
    wire N__44244;
    wire N__44243;
    wire N__44238;
    wire N__44231;
    wire N__44228;
    wire N__44223;
    wire N__44214;
    wire N__44205;
    wire N__44196;
    wire N__44193;
    wire N__44188;
    wire N__44185;
    wire N__44182;
    wire N__44179;
    wire N__44176;
    wire N__44165;
    wire N__44160;
    wire N__44155;
    wire N__44148;
    wire N__44141;
    wire N__44140;
    wire N__44139;
    wire N__44134;
    wire N__44131;
    wire N__44126;
    wire N__44123;
    wire N__44122;
    wire N__44121;
    wire N__44118;
    wire N__44115;
    wire N__44112;
    wire N__44109;
    wire N__44106;
    wire N__44099;
    wire N__44096;
    wire N__44095;
    wire N__44092;
    wire N__44089;
    wire N__44086;
    wire N__44083;
    wire N__44078;
    wire N__44077;
    wire N__44074;
    wire N__44071;
    wire N__44068;
    wire N__44065;
    wire N__44062;
    wire N__44059;
    wire N__44054;
    wire N__44053;
    wire N__44050;
    wire N__44045;
    wire N__44044;
    wire N__44041;
    wire N__44040;
    wire N__44037;
    wire N__44034;
    wire N__44031;
    wire N__44028;
    wire N__44021;
    wire N__44018;
    wire N__44015;
    wire N__44012;
    wire N__44009;
    wire N__44006;
    wire N__44003;
    wire N__44000;
    wire N__43997;
    wire N__43994;
    wire N__43991;
    wire N__43988;
    wire N__43985;
    wire N__43982;
    wire N__43979;
    wire N__43976;
    wire N__43973;
    wire N__43970;
    wire N__43967;
    wire N__43964;
    wire N__43961;
    wire N__43958;
    wire N__43955;
    wire N__43952;
    wire N__43949;
    wire N__43946;
    wire N__43943;
    wire N__43940;
    wire N__43937;
    wire N__43934;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43926;
    wire N__43925;
    wire N__43922;
    wire N__43919;
    wire N__43916;
    wire N__43913;
    wire N__43908;
    wire N__43901;
    wire N__43898;
    wire N__43897;
    wire N__43896;
    wire N__43895;
    wire N__43892;
    wire N__43889;
    wire N__43884;
    wire N__43881;
    wire N__43878;
    wire N__43877;
    wire N__43874;
    wire N__43869;
    wire N__43866;
    wire N__43863;
    wire N__43860;
    wire N__43855;
    wire N__43850;
    wire N__43847;
    wire N__43846;
    wire N__43845;
    wire N__43842;
    wire N__43839;
    wire N__43836;
    wire N__43835;
    wire N__43832;
    wire N__43829;
    wire N__43826;
    wire N__43825;
    wire N__43822;
    wire N__43817;
    wire N__43814;
    wire N__43811;
    wire N__43808;
    wire N__43805;
    wire N__43800;
    wire N__43793;
    wire N__43792;
    wire N__43789;
    wire N__43786;
    wire N__43783;
    wire N__43782;
    wire N__43777;
    wire N__43774;
    wire N__43769;
    wire N__43766;
    wire N__43763;
    wire N__43762;
    wire N__43759;
    wire N__43756;
    wire N__43753;
    wire N__43748;
    wire N__43745;
    wire N__43742;
    wire N__43741;
    wire N__43740;
    wire N__43737;
    wire N__43734;
    wire N__43731;
    wire N__43728;
    wire N__43725;
    wire N__43722;
    wire N__43719;
    wire N__43716;
    wire N__43713;
    wire N__43710;
    wire N__43707;
    wire N__43700;
    wire N__43697;
    wire N__43694;
    wire N__43691;
    wire N__43688;
    wire N__43685;
    wire N__43682;
    wire N__43679;
    wire N__43678;
    wire N__43677;
    wire N__43674;
    wire N__43671;
    wire N__43668;
    wire N__43665;
    wire N__43664;
    wire N__43663;
    wire N__43660;
    wire N__43657;
    wire N__43654;
    wire N__43651;
    wire N__43650;
    wire N__43647;
    wire N__43644;
    wire N__43641;
    wire N__43636;
    wire N__43633;
    wire N__43628;
    wire N__43623;
    wire N__43616;
    wire N__43613;
    wire N__43612;
    wire N__43609;
    wire N__43608;
    wire N__43605;
    wire N__43602;
    wire N__43599;
    wire N__43592;
    wire N__43589;
    wire N__43586;
    wire N__43583;
    wire N__43580;
    wire N__43577;
    wire N__43574;
    wire N__43573;
    wire N__43572;
    wire N__43569;
    wire N__43566;
    wire N__43565;
    wire N__43562;
    wire N__43561;
    wire N__43558;
    wire N__43555;
    wire N__43552;
    wire N__43547;
    wire N__43538;
    wire N__43537;
    wire N__43532;
    wire N__43529;
    wire N__43526;
    wire N__43525;
    wire N__43524;
    wire N__43523;
    wire N__43520;
    wire N__43513;
    wire N__43508;
    wire N__43505;
    wire N__43502;
    wire N__43499;
    wire N__43498;
    wire N__43497;
    wire N__43496;
    wire N__43493;
    wire N__43488;
    wire N__43485;
    wire N__43478;
    wire N__43475;
    wire N__43474;
    wire N__43471;
    wire N__43468;
    wire N__43463;
    wire N__43460;
    wire N__43457;
    wire N__43454;
    wire N__43453;
    wire N__43450;
    wire N__43447;
    wire N__43442;
    wire N__43439;
    wire N__43438;
    wire N__43433;
    wire N__43430;
    wire N__43429;
    wire N__43428;
    wire N__43427;
    wire N__43426;
    wire N__43423;
    wire N__43420;
    wire N__43417;
    wire N__43414;
    wire N__43411;
    wire N__43408;
    wire N__43405;
    wire N__43398;
    wire N__43393;
    wire N__43390;
    wire N__43385;
    wire N__43382;
    wire N__43379;
    wire N__43378;
    wire N__43377;
    wire N__43374;
    wire N__43369;
    wire N__43366;
    wire N__43361;
    wire N__43358;
    wire N__43355;
    wire N__43352;
    wire N__43351;
    wire N__43348;
    wire N__43345;
    wire N__43340;
    wire N__43337;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43329;
    wire N__43324;
    wire N__43323;
    wire N__43320;
    wire N__43317;
    wire N__43314;
    wire N__43307;
    wire N__43306;
    wire N__43303;
    wire N__43300;
    wire N__43297;
    wire N__43294;
    wire N__43289;
    wire N__43286;
    wire N__43283;
    wire N__43280;
    wire N__43279;
    wire N__43276;
    wire N__43273;
    wire N__43268;
    wire N__43267;
    wire N__43264;
    wire N__43261;
    wire N__43258;
    wire N__43255;
    wire N__43252;
    wire N__43249;
    wire N__43244;
    wire N__43241;
    wire N__43240;
    wire N__43237;
    wire N__43234;
    wire N__43229;
    wire N__43228;
    wire N__43225;
    wire N__43222;
    wire N__43219;
    wire N__43216;
    wire N__43213;
    wire N__43210;
    wire N__43205;
    wire N__43204;
    wire N__43201;
    wire N__43198;
    wire N__43193;
    wire N__43190;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43172;
    wire N__43171;
    wire N__43170;
    wire N__43169;
    wire N__43168;
    wire N__43167;
    wire N__43164;
    wire N__43161;
    wire N__43158;
    wire N__43157;
    wire N__43156;
    wire N__43153;
    wire N__43152;
    wire N__43149;
    wire N__43148;
    wire N__43147;
    wire N__43146;
    wire N__43145;
    wire N__43142;
    wire N__43141;
    wire N__43140;
    wire N__43139;
    wire N__43138;
    wire N__43137;
    wire N__43134;
    wire N__43127;
    wire N__43122;
    wire N__43121;
    wire N__43118;
    wire N__43115;
    wire N__43108;
    wire N__43107;
    wire N__43104;
    wire N__43103;
    wire N__43102;
    wire N__43101;
    wire N__43100;
    wire N__43099;
    wire N__43096;
    wire N__43093;
    wire N__43090;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43074;
    wire N__43073;
    wire N__43072;
    wire N__43071;
    wire N__43070;
    wire N__43069;
    wire N__43066;
    wire N__43059;
    wire N__43052;
    wire N__43049;
    wire N__43042;
    wire N__43031;
    wire N__43026;
    wire N__43013;
    wire N__43008;
    wire N__42995;
    wire N__42994;
    wire N__42993;
    wire N__42992;
    wire N__42991;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42983;
    wire N__42982;
    wire N__42979;
    wire N__42976;
    wire N__42975;
    wire N__42972;
    wire N__42971;
    wire N__42968;
    wire N__42963;
    wire N__42962;
    wire N__42959;
    wire N__42958;
    wire N__42957;
    wire N__42956;
    wire N__42953;
    wire N__42952;
    wire N__42951;
    wire N__42950;
    wire N__42947;
    wire N__42944;
    wire N__42943;
    wire N__42942;
    wire N__42941;
    wire N__42940;
    wire N__42937;
    wire N__42934;
    wire N__42931;
    wire N__42926;
    wire N__42923;
    wire N__42916;
    wire N__42913;
    wire N__42908;
    wire N__42903;
    wire N__42898;
    wire N__42889;
    wire N__42886;
    wire N__42881;
    wire N__42878;
    wire N__42857;
    wire N__42854;
    wire N__42853;
    wire N__42850;
    wire N__42847;
    wire N__42842;
    wire N__42839;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42827;
    wire N__42824;
    wire N__42823;
    wire N__42820;
    wire N__42817;
    wire N__42814;
    wire N__42811;
    wire N__42810;
    wire N__42807;
    wire N__42804;
    wire N__42801;
    wire N__42794;
    wire N__42791;
    wire N__42790;
    wire N__42789;
    wire N__42786;
    wire N__42785;
    wire N__42782;
    wire N__42779;
    wire N__42776;
    wire N__42771;
    wire N__42768;
    wire N__42765;
    wire N__42762;
    wire N__42755;
    wire N__42752;
    wire N__42749;
    wire N__42746;
    wire N__42745;
    wire N__42742;
    wire N__42741;
    wire N__42738;
    wire N__42737;
    wire N__42736;
    wire N__42735;
    wire N__42734;
    wire N__42733;
    wire N__42730;
    wire N__42727;
    wire N__42724;
    wire N__42721;
    wire N__42716;
    wire N__42713;
    wire N__42710;
    wire N__42699;
    wire N__42696;
    wire N__42695;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42674;
    wire N__42671;
    wire N__42670;
    wire N__42667;
    wire N__42664;
    wire N__42659;
    wire N__42656;
    wire N__42653;
    wire N__42650;
    wire N__42647;
    wire N__42644;
    wire N__42643;
    wire N__42640;
    wire N__42637;
    wire N__42632;
    wire N__42631;
    wire N__42630;
    wire N__42627;
    wire N__42622;
    wire N__42617;
    wire N__42614;
    wire N__42613;
    wire N__42612;
    wire N__42609;
    wire N__42604;
    wire N__42599;
    wire N__42596;
    wire N__42595;
    wire N__42592;
    wire N__42589;
    wire N__42586;
    wire N__42581;
    wire N__42580;
    wire N__42575;
    wire N__42572;
    wire N__42571;
    wire N__42568;
    wire N__42565;
    wire N__42560;
    wire N__42557;
    wire N__42554;
    wire N__42551;
    wire N__42548;
    wire N__42545;
    wire N__42544;
    wire N__42541;
    wire N__42538;
    wire N__42533;
    wire N__42530;
    wire N__42529;
    wire N__42526;
    wire N__42523;
    wire N__42518;
    wire N__42517;
    wire N__42514;
    wire N__42511;
    wire N__42508;
    wire N__42505;
    wire N__42502;
    wire N__42499;
    wire N__42494;
    wire N__42491;
    wire N__42488;
    wire N__42487;
    wire N__42486;
    wire N__42483;
    wire N__42480;
    wire N__42477;
    wire N__42474;
    wire N__42471;
    wire N__42468;
    wire N__42467;
    wire N__42464;
    wire N__42461;
    wire N__42458;
    wire N__42455;
    wire N__42446;
    wire N__42445;
    wire N__42442;
    wire N__42441;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42429;
    wire N__42426;
    wire N__42423;
    wire N__42420;
    wire N__42415;
    wire N__42410;
    wire N__42407;
    wire N__42404;
    wire N__42401;
    wire N__42398;
    wire N__42395;
    wire N__42394;
    wire N__42391;
    wire N__42388;
    wire N__42387;
    wire N__42386;
    wire N__42383;
    wire N__42380;
    wire N__42377;
    wire N__42374;
    wire N__42371;
    wire N__42368;
    wire N__42365;
    wire N__42362;
    wire N__42353;
    wire N__42350;
    wire N__42347;
    wire N__42344;
    wire N__42341;
    wire N__42340;
    wire N__42337;
    wire N__42334;
    wire N__42331;
    wire N__42330;
    wire N__42327;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42315;
    wire N__42312;
    wire N__42311;
    wire N__42308;
    wire N__42303;
    wire N__42300;
    wire N__42293;
    wire N__42292;
    wire N__42291;
    wire N__42288;
    wire N__42285;
    wire N__42282;
    wire N__42279;
    wire N__42276;
    wire N__42271;
    wire N__42266;
    wire N__42263;
    wire N__42260;
    wire N__42257;
    wire N__42256;
    wire N__42255;
    wire N__42254;
    wire N__42253;
    wire N__42252;
    wire N__42251;
    wire N__42250;
    wire N__42249;
    wire N__42248;
    wire N__42247;
    wire N__42246;
    wire N__42245;
    wire N__42242;
    wire N__42241;
    wire N__42240;
    wire N__42239;
    wire N__42238;
    wire N__42235;
    wire N__42232;
    wire N__42221;
    wire N__42220;
    wire N__42219;
    wire N__42218;
    wire N__42217;
    wire N__42216;
    wire N__42205;
    wire N__42202;
    wire N__42193;
    wire N__42192;
    wire N__42191;
    wire N__42190;
    wire N__42185;
    wire N__42182;
    wire N__42179;
    wire N__42174;
    wire N__42169;
    wire N__42162;
    wire N__42159;
    wire N__42156;
    wire N__42153;
    wire N__42148;
    wire N__42141;
    wire N__42138;
    wire N__42133;
    wire N__42122;
    wire N__42121;
    wire N__42118;
    wire N__42115;
    wire N__42112;
    wire N__42111;
    wire N__42108;
    wire N__42105;
    wire N__42102;
    wire N__42101;
    wire N__42096;
    wire N__42093;
    wire N__42090;
    wire N__42083;
    wire N__42082;
    wire N__42081;
    wire N__42078;
    wire N__42075;
    wire N__42072;
    wire N__42067;
    wire N__42064;
    wire N__42061;
    wire N__42056;
    wire N__42053;
    wire N__42050;
    wire N__42047;
    wire N__42044;
    wire N__42043;
    wire N__42040;
    wire N__42039;
    wire N__42038;
    wire N__42035;
    wire N__42032;
    wire N__42027;
    wire N__42024;
    wire N__42019;
    wire N__42014;
    wire N__42011;
    wire N__42010;
    wire N__42007;
    wire N__42004;
    wire N__42003;
    wire N__42000;
    wire N__41997;
    wire N__41994;
    wire N__41987;
    wire N__41986;
    wire N__41983;
    wire N__41982;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41972;
    wire N__41969;
    wire N__41966;
    wire N__41963;
    wire N__41962;
    wire N__41959;
    wire N__41956;
    wire N__41953;
    wire N__41950;
    wire N__41947;
    wire N__41946;
    wire N__41943;
    wire N__41938;
    wire N__41935;
    wire N__41932;
    wire N__41929;
    wire N__41926;
    wire N__41923;
    wire N__41918;
    wire N__41909;
    wire N__41906;
    wire N__41903;
    wire N__41900;
    wire N__41899;
    wire N__41896;
    wire N__41893;
    wire N__41888;
    wire N__41887;
    wire N__41884;
    wire N__41881;
    wire N__41880;
    wire N__41879;
    wire N__41876;
    wire N__41873;
    wire N__41868;
    wire N__41865;
    wire N__41858;
    wire N__41857;
    wire N__41854;
    wire N__41851;
    wire N__41850;
    wire N__41847;
    wire N__41846;
    wire N__41843;
    wire N__41840;
    wire N__41837;
    wire N__41834;
    wire N__41831;
    wire N__41830;
    wire N__41827;
    wire N__41822;
    wire N__41819;
    wire N__41816;
    wire N__41813;
    wire N__41804;
    wire N__41801;
    wire N__41798;
    wire N__41797;
    wire N__41794;
    wire N__41791;
    wire N__41786;
    wire N__41785;
    wire N__41782;
    wire N__41779;
    wire N__41778;
    wire N__41775;
    wire N__41772;
    wire N__41769;
    wire N__41768;
    wire N__41765;
    wire N__41760;
    wire N__41757;
    wire N__41750;
    wire N__41749;
    wire N__41746;
    wire N__41743;
    wire N__41740;
    wire N__41737;
    wire N__41734;
    wire N__41733;
    wire N__41730;
    wire N__41727;
    wire N__41724;
    wire N__41717;
    wire N__41716;
    wire N__41715;
    wire N__41712;
    wire N__41711;
    wire N__41710;
    wire N__41705;
    wire N__41704;
    wire N__41703;
    wire N__41702;
    wire N__41701;
    wire N__41700;
    wire N__41699;
    wire N__41698;
    wire N__41697;
    wire N__41696;
    wire N__41695;
    wire N__41694;
    wire N__41693;
    wire N__41692;
    wire N__41691;
    wire N__41690;
    wire N__41689;
    wire N__41688;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41676;
    wire N__41671;
    wire N__41668;
    wire N__41663;
    wire N__41656;
    wire N__41649;
    wire N__41638;
    wire N__41635;
    wire N__41630;
    wire N__41609;
    wire N__41606;
    wire N__41605;
    wire N__41602;
    wire N__41601;
    wire N__41598;
    wire N__41595;
    wire N__41590;
    wire N__41587;
    wire N__41584;
    wire N__41579;
    wire N__41576;
    wire N__41575;
    wire N__41574;
    wire N__41573;
    wire N__41570;
    wire N__41569;
    wire N__41568;
    wire N__41567;
    wire N__41566;
    wire N__41565;
    wire N__41564;
    wire N__41563;
    wire N__41558;
    wire N__41555;
    wire N__41552;
    wire N__41551;
    wire N__41550;
    wire N__41549;
    wire N__41546;
    wire N__41545;
    wire N__41544;
    wire N__41541;
    wire N__41534;
    wire N__41531;
    wire N__41530;
    wire N__41527;
    wire N__41524;
    wire N__41523;
    wire N__41522;
    wire N__41521;
    wire N__41520;
    wire N__41519;
    wire N__41518;
    wire N__41515;
    wire N__41512;
    wire N__41511;
    wire N__41508;
    wire N__41505;
    wire N__41504;
    wire N__41501;
    wire N__41500;
    wire N__41499;
    wire N__41498;
    wire N__41497;
    wire N__41496;
    wire N__41493;
    wire N__41490;
    wire N__41487;
    wire N__41484;
    wire N__41481;
    wire N__41478;
    wire N__41475;
    wire N__41472;
    wire N__41469;
    wire N__41464;
    wire N__41461;
    wire N__41454;
    wire N__41449;
    wire N__41444;
    wire N__41441;
    wire N__41434;
    wire N__41425;
    wire N__41416;
    wire N__41387;
    wire N__41386;
    wire N__41383;
    wire N__41380;
    wire N__41377;
    wire N__41374;
    wire N__41373;
    wire N__41370;
    wire N__41367;
    wire N__41364;
    wire N__41359;
    wire N__41354;
    wire N__41353;
    wire N__41350;
    wire N__41347;
    wire N__41344;
    wire N__41341;
    wire N__41340;
    wire N__41337;
    wire N__41334;
    wire N__41331;
    wire N__41328;
    wire N__41325;
    wire N__41322;
    wire N__41321;
    wire N__41318;
    wire N__41313;
    wire N__41310;
    wire N__41303;
    wire N__41302;
    wire N__41299;
    wire N__41296;
    wire N__41293;
    wire N__41292;
    wire N__41289;
    wire N__41286;
    wire N__41283;
    wire N__41276;
    wire N__41273;
    wire N__41270;
    wire N__41267;
    wire N__41264;
    wire N__41261;
    wire N__41260;
    wire N__41257;
    wire N__41254;
    wire N__41253;
    wire N__41250;
    wire N__41247;
    wire N__41244;
    wire N__41241;
    wire N__41236;
    wire N__41231;
    wire N__41228;
    wire N__41227;
    wire N__41226;
    wire N__41223;
    wire N__41218;
    wire N__41215;
    wire N__41212;
    wire N__41211;
    wire N__41206;
    wire N__41203;
    wire N__41198;
    wire N__41197;
    wire N__41196;
    wire N__41189;
    wire N__41186;
    wire N__41183;
    wire N__41182;
    wire N__41179;
    wire N__41176;
    wire N__41171;
    wire N__41168;
    wire N__41167;
    wire N__41166;
    wire N__41159;
    wire N__41156;
    wire N__41153;
    wire N__41150;
    wire N__41147;
    wire N__41144;
    wire N__41141;
    wire N__41138;
    wire N__41135;
    wire N__41132;
    wire N__41129;
    wire N__41126;
    wire N__41123;
    wire N__41120;
    wire N__41117;
    wire N__41116;
    wire N__41115;
    wire N__41108;
    wire N__41105;
    wire N__41102;
    wire N__41101;
    wire N__41098;
    wire N__41095;
    wire N__41090;
    wire N__41087;
    wire N__41086;
    wire N__41085;
    wire N__41078;
    wire N__41075;
    wire N__41072;
    wire N__41069;
    wire N__41066;
    wire N__41063;
    wire N__41060;
    wire N__41057;
    wire N__41054;
    wire N__41053;
    wire N__41052;
    wire N__41049;
    wire N__41046;
    wire N__41043;
    wire N__41038;
    wire N__41035;
    wire N__41030;
    wire N__41027;
    wire N__41024;
    wire N__41023;
    wire N__41022;
    wire N__41021;
    wire N__41020;
    wire N__41019;
    wire N__41018;
    wire N__41017;
    wire N__41016;
    wire N__40997;
    wire N__40994;
    wire N__40991;
    wire N__40988;
    wire N__40985;
    wire N__40982;
    wire N__40979;
    wire N__40976;
    wire N__40973;
    wire N__40970;
    wire N__40967;
    wire N__40964;
    wire N__40961;
    wire N__40958;
    wire N__40955;
    wire N__40952;
    wire N__40949;
    wire N__40946;
    wire N__40943;
    wire N__40940;
    wire N__40937;
    wire N__40936;
    wire N__40935;
    wire N__40934;
    wire N__40933;
    wire N__40932;
    wire N__40931;
    wire N__40930;
    wire N__40929;
    wire N__40928;
    wire N__40927;
    wire N__40926;
    wire N__40925;
    wire N__40922;
    wire N__40913;
    wire N__40902;
    wire N__40895;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40877;
    wire N__40874;
    wire N__40871;
    wire N__40868;
    wire N__40867;
    wire N__40864;
    wire N__40861;
    wire N__40858;
    wire N__40853;
    wire N__40850;
    wire N__40847;
    wire N__40846;
    wire N__40843;
    wire N__40840;
    wire N__40837;
    wire N__40832;
    wire N__40829;
    wire N__40828;
    wire N__40825;
    wire N__40822;
    wire N__40819;
    wire N__40814;
    wire N__40811;
    wire N__40810;
    wire N__40807;
    wire N__40804;
    wire N__40801;
    wire N__40796;
    wire N__40793;
    wire N__40792;
    wire N__40789;
    wire N__40786;
    wire N__40783;
    wire N__40778;
    wire N__40775;
    wire N__40772;
    wire N__40771;
    wire N__40768;
    wire N__40765;
    wire N__40762;
    wire N__40757;
    wire N__40754;
    wire N__40751;
    wire N__40748;
    wire N__40745;
    wire N__40744;
    wire N__40741;
    wire N__40738;
    wire N__40735;
    wire N__40730;
    wire N__40727;
    wire N__40726;
    wire N__40723;
    wire N__40720;
    wire N__40717;
    wire N__40712;
    wire N__40709;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40699;
    wire N__40694;
    wire N__40691;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40676;
    wire N__40673;
    wire N__40672;
    wire N__40669;
    wire N__40666;
    wire N__40663;
    wire N__40658;
    wire N__40655;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40645;
    wire N__40640;
    wire N__40637;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40627;
    wire N__40622;
    wire N__40619;
    wire N__40618;
    wire N__40615;
    wire N__40612;
    wire N__40609;
    wire N__40604;
    wire N__40601;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40586;
    wire N__40583;
    wire N__40580;
    wire N__40577;
    wire N__40576;
    wire N__40573;
    wire N__40570;
    wire N__40565;
    wire N__40564;
    wire N__40561;
    wire N__40558;
    wire N__40555;
    wire N__40552;
    wire N__40551;
    wire N__40548;
    wire N__40545;
    wire N__40542;
    wire N__40539;
    wire N__40534;
    wire N__40531;
    wire N__40528;
    wire N__40525;
    wire N__40522;
    wire N__40517;
    wire N__40514;
    wire N__40513;
    wire N__40510;
    wire N__40507;
    wire N__40502;
    wire N__40499;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40489;
    wire N__40486;
    wire N__40483;
    wire N__40480;
    wire N__40475;
    wire N__40472;
    wire N__40471;
    wire N__40468;
    wire N__40465;
    wire N__40462;
    wire N__40457;
    wire N__40454;
    wire N__40453;
    wire N__40450;
    wire N__40447;
    wire N__40444;
    wire N__40439;
    wire N__40436;
    wire N__40433;
    wire N__40430;
    wire N__40427;
    wire N__40424;
    wire N__40421;
    wire N__40418;
    wire N__40415;
    wire N__40412;
    wire N__40409;
    wire N__40406;
    wire N__40403;
    wire N__40400;
    wire N__40397;
    wire N__40394;
    wire N__40391;
    wire N__40388;
    wire N__40385;
    wire N__40382;
    wire N__40379;
    wire N__40376;
    wire N__40373;
    wire N__40370;
    wire N__40367;
    wire N__40364;
    wire N__40361;
    wire N__40358;
    wire N__40355;
    wire N__40352;
    wire N__40349;
    wire N__40346;
    wire N__40343;
    wire N__40340;
    wire N__40337;
    wire N__40334;
    wire N__40331;
    wire N__40328;
    wire N__40325;
    wire N__40322;
    wire N__40319;
    wire N__40316;
    wire N__40313;
    wire N__40310;
    wire N__40307;
    wire N__40304;
    wire N__40301;
    wire N__40298;
    wire N__40295;
    wire N__40292;
    wire N__40289;
    wire N__40286;
    wire N__40283;
    wire N__40280;
    wire N__40277;
    wire N__40274;
    wire N__40271;
    wire N__40268;
    wire N__40265;
    wire N__40262;
    wire N__40259;
    wire N__40256;
    wire N__40253;
    wire N__40250;
    wire N__40247;
    wire N__40244;
    wire N__40241;
    wire N__40238;
    wire N__40235;
    wire N__40232;
    wire N__40229;
    wire N__40226;
    wire N__40223;
    wire N__40220;
    wire N__40217;
    wire N__40214;
    wire N__40211;
    wire N__40208;
    wire N__40205;
    wire N__40202;
    wire N__40199;
    wire N__40196;
    wire N__40193;
    wire N__40190;
    wire N__40187;
    wire N__40184;
    wire N__40181;
    wire N__40178;
    wire N__40175;
    wire N__40172;
    wire N__40169;
    wire N__40166;
    wire N__40163;
    wire N__40160;
    wire N__40157;
    wire N__40154;
    wire N__40151;
    wire N__40148;
    wire N__40145;
    wire N__40142;
    wire N__40139;
    wire N__40136;
    wire N__40133;
    wire N__40130;
    wire N__40127;
    wire N__40124;
    wire N__40121;
    wire N__40118;
    wire N__40115;
    wire N__40112;
    wire N__40109;
    wire N__40106;
    wire N__40103;
    wire N__40100;
    wire N__40097;
    wire N__40094;
    wire N__40091;
    wire N__40088;
    wire N__40085;
    wire N__40082;
    wire N__40081;
    wire N__40080;
    wire N__40077;
    wire N__40076;
    wire N__40075;
    wire N__40070;
    wire N__40067;
    wire N__40062;
    wire N__40059;
    wire N__40052;
    wire N__40049;
    wire N__40046;
    wire N__40043;
    wire N__40040;
    wire N__40039;
    wire N__40036;
    wire N__40033;
    wire N__40028;
    wire N__40025;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40017;
    wire N__40014;
    wire N__40011;
    wire N__40008;
    wire N__40001;
    wire N__40000;
    wire N__39999;
    wire N__39998;
    wire N__39997;
    wire N__39994;
    wire N__39993;
    wire N__39992;
    wire N__39991;
    wire N__39990;
    wire N__39989;
    wire N__39988;
    wire N__39985;
    wire N__39982;
    wire N__39977;
    wire N__39974;
    wire N__39971;
    wire N__39964;
    wire N__39955;
    wire N__39950;
    wire N__39941;
    wire N__39938;
    wire N__39935;
    wire N__39932;
    wire N__39929;
    wire N__39926;
    wire N__39923;
    wire N__39920;
    wire N__39919;
    wire N__39918;
    wire N__39917;
    wire N__39914;
    wire N__39911;
    wire N__39906;
    wire N__39899;
    wire N__39898;
    wire N__39897;
    wire N__39896;
    wire N__39895;
    wire N__39894;
    wire N__39893;
    wire N__39892;
    wire N__39891;
    wire N__39890;
    wire N__39889;
    wire N__39888;
    wire N__39887;
    wire N__39886;
    wire N__39885;
    wire N__39884;
    wire N__39883;
    wire N__39882;
    wire N__39881;
    wire N__39880;
    wire N__39879;
    wire N__39878;
    wire N__39877;
    wire N__39876;
    wire N__39875;
    wire N__39874;
    wire N__39873;
    wire N__39866;
    wire N__39865;
    wire N__39864;
    wire N__39863;
    wire N__39862;
    wire N__39861;
    wire N__39860;
    wire N__39859;
    wire N__39858;
    wire N__39853;
    wire N__39844;
    wire N__39841;
    wire N__39836;
    wire N__39829;
    wire N__39822;
    wire N__39807;
    wire N__39802;
    wire N__39799;
    wire N__39788;
    wire N__39781;
    wire N__39772;
    wire N__39755;
    wire N__39754;
    wire N__39753;
    wire N__39752;
    wire N__39751;
    wire N__39748;
    wire N__39745;
    wire N__39744;
    wire N__39743;
    wire N__39742;
    wire N__39741;
    wire N__39740;
    wire N__39739;
    wire N__39738;
    wire N__39737;
    wire N__39736;
    wire N__39735;
    wire N__39734;
    wire N__39733;
    wire N__39732;
    wire N__39731;
    wire N__39730;
    wire N__39729;
    wire N__39728;
    wire N__39717;
    wire N__39716;
    wire N__39715;
    wire N__39714;
    wire N__39703;
    wire N__39698;
    wire N__39691;
    wire N__39688;
    wire N__39685;
    wire N__39678;
    wire N__39677;
    wire N__39674;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39660;
    wire N__39653;
    wire N__39646;
    wire N__39643;
    wire N__39636;
    wire N__39633;
    wire N__39628;
    wire N__39623;
    wire N__39620;
    wire N__39611;
    wire N__39608;
    wire N__39605;
    wire N__39602;
    wire N__39599;
    wire N__39598;
    wire N__39597;
    wire N__39594;
    wire N__39591;
    wire N__39590;
    wire N__39589;
    wire N__39588;
    wire N__39587;
    wire N__39586;
    wire N__39585;
    wire N__39582;
    wire N__39581;
    wire N__39580;
    wire N__39579;
    wire N__39578;
    wire N__39575;
    wire N__39572;
    wire N__39563;
    wire N__39560;
    wire N__39557;
    wire N__39554;
    wire N__39553;
    wire N__39552;
    wire N__39551;
    wire N__39550;
    wire N__39549;
    wire N__39548;
    wire N__39547;
    wire N__39546;
    wire N__39545;
    wire N__39544;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39524;
    wire N__39519;
    wire N__39512;
    wire N__39509;
    wire N__39504;
    wire N__39495;
    wire N__39490;
    wire N__39485;
    wire N__39482;
    wire N__39467;
    wire N__39464;
    wire N__39461;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39437;
    wire N__39434;
    wire N__39431;
    wire N__39428;
    wire N__39425;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39404;
    wire N__39401;
    wire N__39398;
    wire N__39397;
    wire N__39394;
    wire N__39391;
    wire N__39386;
    wire N__39383;
    wire N__39382;
    wire N__39379;
    wire N__39376;
    wire N__39371;
    wire N__39370;
    wire N__39367;
    wire N__39364;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39356;
    wire N__39353;
    wire N__39348;
    wire N__39345;
    wire N__39342;
    wire N__39337;
    wire N__39332;
    wire N__39331;
    wire N__39328;
    wire N__39325;
    wire N__39322;
    wire N__39317;
    wire N__39316;
    wire N__39311;
    wire N__39308;
    wire N__39305;
    wire N__39304;
    wire N__39301;
    wire N__39298;
    wire N__39293;
    wire N__39290;
    wire N__39287;
    wire N__39286;
    wire N__39283;
    wire N__39280;
    wire N__39275;
    wire N__39274;
    wire N__39269;
    wire N__39266;
    wire N__39263;
    wire N__39262;
    wire N__39259;
    wire N__39256;
    wire N__39253;
    wire N__39252;
    wire N__39247;
    wire N__39244;
    wire N__39239;
    wire N__39236;
    wire N__39233;
    wire N__39232;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39217;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39207;
    wire N__39200;
    wire N__39199;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39181;
    wire N__39178;
    wire N__39173;
    wire N__39170;
    wire N__39169;
    wire N__39164;
    wire N__39161;
    wire N__39158;
    wire N__39155;
    wire N__39152;
    wire N__39149;
    wire N__39146;
    wire N__39143;
    wire N__39140;
    wire N__39139;
    wire N__39138;
    wire N__39137;
    wire N__39136;
    wire N__39135;
    wire N__39134;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39113;
    wire N__39110;
    wire N__39109;
    wire N__39104;
    wire N__39099;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39082;
    wire N__39079;
    wire N__39068;
    wire N__39065;
    wire N__39064;
    wire N__39063;
    wire N__39062;
    wire N__39059;
    wire N__39056;
    wire N__39051;
    wire N__39044;
    wire N__39041;
    wire N__39040;
    wire N__39037;
    wire N__39034;
    wire N__39033;
    wire N__39030;
    wire N__39025;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39013;
    wire N__39012;
    wire N__39011;
    wire N__39008;
    wire N__39005;
    wire N__39000;
    wire N__38993;
    wire N__38992;
    wire N__38991;
    wire N__38984;
    wire N__38981;
    wire N__38978;
    wire N__38977;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38966;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38939;
    wire N__38936;
    wire N__38933;
    wire N__38930;
    wire N__38929;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38915;
    wire N__38912;
    wire N__38911;
    wire N__38910;
    wire N__38909;
    wire N__38908;
    wire N__38907;
    wire N__38906;
    wire N__38905;
    wire N__38904;
    wire N__38903;
    wire N__38902;
    wire N__38901;
    wire N__38900;
    wire N__38899;
    wire N__38898;
    wire N__38897;
    wire N__38888;
    wire N__38879;
    wire N__38878;
    wire N__38877;
    wire N__38876;
    wire N__38875;
    wire N__38874;
    wire N__38873;
    wire N__38872;
    wire N__38871;
    wire N__38870;
    wire N__38869;
    wire N__38868;
    wire N__38867;
    wire N__38866;
    wire N__38865;
    wire N__38856;
    wire N__38847;
    wire N__38844;
    wire N__38841;
    wire N__38836;
    wire N__38827;
    wire N__38818;
    wire N__38809;
    wire N__38804;
    wire N__38799;
    wire N__38786;
    wire N__38783;
    wire N__38782;
    wire N__38779;
    wire N__38776;
    wire N__38773;
    wire N__38768;
    wire N__38767;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38750;
    wire N__38747;
    wire N__38742;
    wire N__38739;
    wire N__38732;
    wire N__38729;
    wire N__38726;
    wire N__38725;
    wire N__38722;
    wire N__38719;
    wire N__38716;
    wire N__38715;
    wire N__38710;
    wire N__38707;
    wire N__38704;
    wire N__38699;
    wire N__38698;
    wire N__38697;
    wire N__38696;
    wire N__38695;
    wire N__38694;
    wire N__38681;
    wire N__38678;
    wire N__38675;
    wire N__38674;
    wire N__38671;
    wire N__38670;
    wire N__38665;
    wire N__38662;
    wire N__38657;
    wire N__38654;
    wire N__38653;
    wire N__38650;
    wire N__38647;
    wire N__38644;
    wire N__38641;
    wire N__38636;
    wire N__38635;
    wire N__38632;
    wire N__38629;
    wire N__38624;
    wire N__38623;
    wire N__38620;
    wire N__38619;
    wire N__38616;
    wire N__38611;
    wire N__38606;
    wire N__38603;
    wire N__38600;
    wire N__38599;
    wire N__38596;
    wire N__38593;
    wire N__38592;
    wire N__38591;
    wire N__38590;
    wire N__38585;
    wire N__38580;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38564;
    wire N__38561;
    wire N__38558;
    wire N__38557;
    wire N__38554;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38544;
    wire N__38539;
    wire N__38534;
    wire N__38531;
    wire N__38528;
    wire N__38527;
    wire N__38526;
    wire N__38523;
    wire N__38520;
    wire N__38517;
    wire N__38512;
    wire N__38507;
    wire N__38504;
    wire N__38503;
    wire N__38500;
    wire N__38497;
    wire N__38496;
    wire N__38491;
    wire N__38488;
    wire N__38485;
    wire N__38480;
    wire N__38477;
    wire N__38476;
    wire N__38475;
    wire N__38470;
    wire N__38467;
    wire N__38464;
    wire N__38459;
    wire N__38456;
    wire N__38453;
    wire N__38452;
    wire N__38451;
    wire N__38448;
    wire N__38445;
    wire N__38442;
    wire N__38437;
    wire N__38432;
    wire N__38429;
    wire N__38428;
    wire N__38425;
    wire N__38422;
    wire N__38421;
    wire N__38418;
    wire N__38415;
    wire N__38412;
    wire N__38407;
    wire N__38402;
    wire N__38399;
    wire N__38398;
    wire N__38397;
    wire N__38392;
    wire N__38389;
    wire N__38386;
    wire N__38381;
    wire N__38378;
    wire N__38375;
    wire N__38374;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38364;
    wire N__38359;
    wire N__38354;
    wire N__38351;
    wire N__38348;
    wire N__38347;
    wire N__38346;
    wire N__38343;
    wire N__38340;
    wire N__38337;
    wire N__38332;
    wire N__38327;
    wire N__38324;
    wire N__38323;
    wire N__38320;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38310;
    wire N__38305;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38293;
    wire N__38292;
    wire N__38289;
    wire N__38286;
    wire N__38283;
    wire N__38278;
    wire N__38273;
    wire N__38270;
    wire N__38269;
    wire N__38266;
    wire N__38263;
    wire N__38262;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38246;
    wire N__38243;
    wire N__38242;
    wire N__38241;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38225;
    wire N__38222;
    wire N__38219;
    wire N__38218;
    wire N__38217;
    wire N__38214;
    wire N__38211;
    wire N__38208;
    wire N__38203;
    wire N__38198;
    wire N__38195;
    wire N__38194;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38184;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38170;
    wire N__38165;
    wire N__38162;
    wire N__38161;
    wire N__38160;
    wire N__38155;
    wire N__38152;
    wire N__38149;
    wire N__38144;
    wire N__38141;
    wire N__38138;
    wire N__38137;
    wire N__38136;
    wire N__38133;
    wire N__38130;
    wire N__38127;
    wire N__38122;
    wire N__38117;
    wire N__38114;
    wire N__38113;
    wire N__38112;
    wire N__38109;
    wire N__38106;
    wire N__38103;
    wire N__38098;
    wire N__38093;
    wire N__38090;
    wire N__38089;
    wire N__38088;
    wire N__38083;
    wire N__38080;
    wire N__38077;
    wire N__38072;
    wire N__38069;
    wire N__38066;
    wire N__38065;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38050;
    wire N__38045;
    wire N__38042;
    wire N__38041;
    wire N__38038;
    wire N__38035;
    wire N__38034;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38018;
    wire N__38015;
    wire N__38014;
    wire N__38013;
    wire N__38008;
    wire N__38005;
    wire N__38002;
    wire N__37997;
    wire N__37994;
    wire N__37991;
    wire N__37990;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37975;
    wire N__37970;
    wire N__37967;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37959;
    wire N__37956;
    wire N__37953;
    wire N__37950;
    wire N__37945;
    wire N__37940;
    wire N__37937;
    wire N__37936;
    wire N__37935;
    wire N__37930;
    wire N__37927;
    wire N__37924;
    wire N__37919;
    wire N__37916;
    wire N__37915;
    wire N__37914;
    wire N__37913;
    wire N__37912;
    wire N__37911;
    wire N__37908;
    wire N__37907;
    wire N__37904;
    wire N__37903;
    wire N__37900;
    wire N__37899;
    wire N__37898;
    wire N__37897;
    wire N__37896;
    wire N__37895;
    wire N__37892;
    wire N__37891;
    wire N__37888;
    wire N__37887;
    wire N__37886;
    wire N__37885;
    wire N__37884;
    wire N__37883;
    wire N__37882;
    wire N__37881;
    wire N__37880;
    wire N__37879;
    wire N__37864;
    wire N__37859;
    wire N__37846;
    wire N__37843;
    wire N__37842;
    wire N__37839;
    wire N__37838;
    wire N__37835;
    wire N__37834;
    wire N__37831;
    wire N__37830;
    wire N__37829;
    wire N__37826;
    wire N__37825;
    wire N__37822;
    wire N__37821;
    wire N__37818;
    wire N__37817;
    wire N__37814;
    wire N__37813;
    wire N__37812;
    wire N__37811;
    wire N__37810;
    wire N__37809;
    wire N__37808;
    wire N__37807;
    wire N__37806;
    wire N__37805;
    wire N__37804;
    wire N__37803;
    wire N__37796;
    wire N__37779;
    wire N__37764;
    wire N__37763;
    wire N__37762;
    wire N__37759;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37747;
    wire N__37740;
    wire N__37731;
    wire N__37730;
    wire N__37729;
    wire N__37728;
    wire N__37727;
    wire N__37726;
    wire N__37725;
    wire N__37724;
    wire N__37723;
    wire N__37722;
    wire N__37715;
    wire N__37710;
    wire N__37707;
    wire N__37700;
    wire N__37693;
    wire N__37690;
    wire N__37683;
    wire N__37674;
    wire N__37673;
    wire N__37670;
    wire N__37669;
    wire N__37664;
    wire N__37661;
    wire N__37650;
    wire N__37643;
    wire N__37640;
    wire N__37637;
    wire N__37632;
    wire N__37629;
    wire N__37622;
    wire N__37619;
    wire N__37616;
    wire N__37613;
    wire N__37610;
    wire N__37607;
    wire N__37604;
    wire N__37601;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37580;
    wire N__37577;
    wire N__37574;
    wire N__37571;
    wire N__37568;
    wire N__37565;
    wire N__37562;
    wire N__37559;
    wire N__37558;
    wire N__37555;
    wire N__37554;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37542;
    wire N__37535;
    wire N__37532;
    wire N__37529;
    wire N__37528;
    wire N__37525;
    wire N__37522;
    wire N__37519;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37499;
    wire N__37496;
    wire N__37495;
    wire N__37492;
    wire N__37489;
    wire N__37484;
    wire N__37483;
    wire N__37480;
    wire N__37477;
    wire N__37474;
    wire N__37469;
    wire N__37466;
    wire N__37463;
    wire N__37460;
    wire N__37457;
    wire N__37454;
    wire N__37451;
    wire N__37448;
    wire N__37445;
    wire N__37442;
    wire N__37439;
    wire N__37436;
    wire N__37433;
    wire N__37430;
    wire N__37427;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37415;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37397;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37364;
    wire N__37361;
    wire N__37358;
    wire N__37355;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37319;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37295;
    wire N__37292;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37271;
    wire N__37268;
    wire N__37265;
    wire N__37262;
    wire N__37259;
    wire N__37256;
    wire N__37253;
    wire N__37250;
    wire N__37247;
    wire N__37244;
    wire N__37241;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37228;
    wire N__37223;
    wire N__37220;
    wire N__37217;
    wire N__37216;
    wire N__37215;
    wire N__37212;
    wire N__37207;
    wire N__37202;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37094;
    wire N__37091;
    wire N__37088;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37046;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37033;
    wire N__37030;
    wire N__37027;
    wire N__37024;
    wire N__37021;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36985;
    wire N__36982;
    wire N__36981;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36969;
    wire N__36966;
    wire N__36963;
    wire N__36960;
    wire N__36955;
    wire N__36950;
    wire N__36947;
    wire N__36944;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36934;
    wire N__36931;
    wire N__36928;
    wire N__36925;
    wire N__36922;
    wire N__36917;
    wire N__36916;
    wire N__36913;
    wire N__36910;
    wire N__36905;
    wire N__36902;
    wire N__36899;
    wire N__36896;
    wire N__36893;
    wire N__36890;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36875;
    wire N__36872;
    wire N__36869;
    wire N__36866;
    wire N__36863;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36844;
    wire N__36839;
    wire N__36836;
    wire N__36835;
    wire N__36834;
    wire N__36831;
    wire N__36828;
    wire N__36825;
    wire N__36820;
    wire N__36815;
    wire N__36812;
    wire N__36809;
    wire N__36806;
    wire N__36803;
    wire N__36802;
    wire N__36799;
    wire N__36796;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36779;
    wire N__36776;
    wire N__36773;
    wire N__36772;
    wire N__36769;
    wire N__36768;
    wire N__36765;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36751;
    wire N__36750;
    wire N__36747;
    wire N__36744;
    wire N__36741;
    wire N__36734;
    wire N__36731;
    wire N__36728;
    wire N__36727;
    wire N__36726;
    wire N__36723;
    wire N__36718;
    wire N__36713;
    wire N__36712;
    wire N__36711;
    wire N__36706;
    wire N__36703;
    wire N__36700;
    wire N__36695;
    wire N__36692;
    wire N__36691;
    wire N__36690;
    wire N__36685;
    wire N__36682;
    wire N__36679;
    wire N__36674;
    wire N__36671;
    wire N__36670;
    wire N__36667;
    wire N__36666;
    wire N__36663;
    wire N__36660;
    wire N__36657;
    wire N__36652;
    wire N__36647;
    wire N__36644;
    wire N__36643;
    wire N__36640;
    wire N__36639;
    wire N__36636;
    wire N__36633;
    wire N__36630;
    wire N__36625;
    wire N__36620;
    wire N__36617;
    wire N__36616;
    wire N__36613;
    wire N__36610;
    wire N__36609;
    wire N__36604;
    wire N__36601;
    wire N__36598;
    wire N__36593;
    wire N__36590;
    wire N__36589;
    wire N__36586;
    wire N__36583;
    wire N__36582;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36566;
    wire N__36563;
    wire N__36560;
    wire N__36557;
    wire N__36556;
    wire N__36555;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36540;
    wire N__36533;
    wire N__36530;
    wire N__36527;
    wire N__36524;
    wire N__36523;
    wire N__36522;
    wire N__36519;
    wire N__36516;
    wire N__36513;
    wire N__36508;
    wire N__36503;
    wire N__36500;
    wire N__36499;
    wire N__36498;
    wire N__36493;
    wire N__36490;
    wire N__36487;
    wire N__36482;
    wire N__36479;
    wire N__36476;
    wire N__36475;
    wire N__36472;
    wire N__36469;
    wire N__36466;
    wire N__36461;
    wire N__36458;
    wire N__36457;
    wire N__36456;
    wire N__36451;
    wire N__36448;
    wire N__36445;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36433;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36418;
    wire N__36413;
    wire N__36410;
    wire N__36409;
    wire N__36406;
    wire N__36405;
    wire N__36402;
    wire N__36399;
    wire N__36396;
    wire N__36391;
    wire N__36386;
    wire N__36383;
    wire N__36382;
    wire N__36381;
    wire N__36376;
    wire N__36373;
    wire N__36370;
    wire N__36365;
    wire N__36364;
    wire N__36363;
    wire N__36360;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36344;
    wire N__36341;
    wire N__36340;
    wire N__36337;
    wire N__36334;
    wire N__36333;
    wire N__36328;
    wire N__36325;
    wire N__36322;
    wire N__36317;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36309;
    wire N__36306;
    wire N__36303;
    wire N__36300;
    wire N__36297;
    wire N__36292;
    wire N__36287;
    wire N__36284;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36272;
    wire N__36271;
    wire N__36268;
    wire N__36265;
    wire N__36262;
    wire N__36257;
    wire N__36254;
    wire N__36253;
    wire N__36252;
    wire N__36249;
    wire N__36244;
    wire N__36239;
    wire N__36236;
    wire N__36233;
    wire N__36230;
    wire N__36227;
    wire N__36226;
    wire N__36225;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36211;
    wire N__36206;
    wire N__36203;
    wire N__36200;
    wire N__36199;
    wire N__36198;
    wire N__36195;
    wire N__36190;
    wire N__36187;
    wire N__36184;
    wire N__36179;
    wire N__36176;
    wire N__36173;
    wire N__36170;
    wire N__36169;
    wire N__36168;
    wire N__36165;
    wire N__36162;
    wire N__36159;
    wire N__36154;
    wire N__36149;
    wire N__36146;
    wire N__36145;
    wire N__36144;
    wire N__36139;
    wire N__36136;
    wire N__36133;
    wire N__36128;
    wire N__36125;
    wire N__36124;
    wire N__36123;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36107;
    wire N__36104;
    wire N__36103;
    wire N__36100;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36090;
    wire N__36085;
    wire N__36080;
    wire N__36077;
    wire N__36076;
    wire N__36073;
    wire N__36072;
    wire N__36069;
    wire N__36066;
    wire N__36063;
    wire N__36058;
    wire N__36053;
    wire N__36050;
    wire N__36049;
    wire N__36046;
    wire N__36043;
    wire N__36042;
    wire N__36037;
    wire N__36034;
    wire N__36031;
    wire N__36026;
    wire N__36023;
    wire N__36022;
    wire N__36019;
    wire N__36016;
    wire N__36015;
    wire N__36010;
    wire N__36007;
    wire N__36004;
    wire N__35999;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35989;
    wire N__35988;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35956;
    wire N__35955;
    wire N__35952;
    wire N__35949;
    wire N__35946;
    wire N__35941;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35927;
    wire N__35924;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35913;
    wire N__35910;
    wire N__35907;
    wire N__35904;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35890;
    wire N__35887;
    wire N__35886;
    wire N__35883;
    wire N__35880;
    wire N__35877;
    wire N__35872;
    wire N__35867;
    wire N__35864;
    wire N__35861;
    wire N__35860;
    wire N__35857;
    wire N__35854;
    wire N__35849;
    wire N__35846;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35828;
    wire N__35825;
    wire N__35822;
    wire N__35819;
    wire N__35818;
    wire N__35817;
    wire N__35814;
    wire N__35811;
    wire N__35810;
    wire N__35807;
    wire N__35804;
    wire N__35801;
    wire N__35798;
    wire N__35791;
    wire N__35786;
    wire N__35785;
    wire N__35784;
    wire N__35781;
    wire N__35778;
    wire N__35777;
    wire N__35774;
    wire N__35771;
    wire N__35768;
    wire N__35765;
    wire N__35762;
    wire N__35757;
    wire N__35754;
    wire N__35747;
    wire N__35744;
    wire N__35743;
    wire N__35742;
    wire N__35741;
    wire N__35738;
    wire N__35733;
    wire N__35730;
    wire N__35723;
    wire N__35722;
    wire N__35721;
    wire N__35720;
    wire N__35719;
    wire N__35718;
    wire N__35717;
    wire N__35716;
    wire N__35715;
    wire N__35714;
    wire N__35709;
    wire N__35700;
    wire N__35699;
    wire N__35698;
    wire N__35697;
    wire N__35696;
    wire N__35687;
    wire N__35686;
    wire N__35685;
    wire N__35684;
    wire N__35683;
    wire N__35682;
    wire N__35681;
    wire N__35680;
    wire N__35679;
    wire N__35678;
    wire N__35677;
    wire N__35676;
    wire N__35675;
    wire N__35674;
    wire N__35673;
    wire N__35672;
    wire N__35671;
    wire N__35666;
    wire N__35657;
    wire N__35654;
    wire N__35645;
    wire N__35636;
    wire N__35627;
    wire N__35618;
    wire N__35615;
    wire N__35600;
    wire N__35597;
    wire N__35594;
    wire N__35591;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35572;
    wire N__35569;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35559;
    wire N__35556;
    wire N__35551;
    wire N__35550;
    wire N__35547;
    wire N__35544;
    wire N__35541;
    wire N__35534;
    wire N__35531;
    wire N__35528;
    wire N__35525;
    wire N__35522;
    wire N__35519;
    wire N__35516;
    wire N__35515;
    wire N__35512;
    wire N__35509;
    wire N__35508;
    wire N__35503;
    wire N__35500;
    wire N__35499;
    wire N__35496;
    wire N__35493;
    wire N__35490;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35474;
    wire N__35473;
    wire N__35472;
    wire N__35467;
    wire N__35464;
    wire N__35461;
    wire N__35458;
    wire N__35457;
    wire N__35452;
    wire N__35449;
    wire N__35444;
    wire N__35441;
    wire N__35438;
    wire N__35437;
    wire N__35436;
    wire N__35431;
    wire N__35428;
    wire N__35427;
    wire N__35424;
    wire N__35421;
    wire N__35418;
    wire N__35415;
    wire N__35412;
    wire N__35409;
    wire N__35402;
    wire N__35399;
    wire N__35396;
    wire N__35395;
    wire N__35392;
    wire N__35389;
    wire N__35386;
    wire N__35383;
    wire N__35382;
    wire N__35381;
    wire N__35376;
    wire N__35373;
    wire N__35370;
    wire N__35365;
    wire N__35362;
    wire N__35359;
    wire N__35356;
    wire N__35351;
    wire N__35348;
    wire N__35345;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35337;
    wire N__35336;
    wire N__35333;
    wire N__35328;
    wire N__35325;
    wire N__35320;
    wire N__35317;
    wire N__35314;
    wire N__35311;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35294;
    wire N__35293;
    wire N__35290;
    wire N__35287;
    wire N__35284;
    wire N__35279;
    wire N__35278;
    wire N__35275;
    wire N__35274;
    wire N__35271;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35255;
    wire N__35252;
    wire N__35249;
    wire N__35246;
    wire N__35245;
    wire N__35244;
    wire N__35241;
    wire N__35238;
    wire N__35235;
    wire N__35232;
    wire N__35229;
    wire N__35226;
    wire N__35219;
    wire N__35216;
    wire N__35213;
    wire N__35210;
    wire N__35207;
    wire N__35204;
    wire N__35201;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35193;
    wire N__35188;
    wire N__35185;
    wire N__35180;
    wire N__35177;
    wire N__35174;
    wire N__35171;
    wire N__35168;
    wire N__35165;
    wire N__35162;
    wire N__35159;
    wire N__35156;
    wire N__35153;
    wire N__35150;
    wire N__35147;
    wire N__35144;
    wire N__35141;
    wire N__35138;
    wire N__35135;
    wire N__35134;
    wire N__35131;
    wire N__35128;
    wire N__35127;
    wire N__35122;
    wire N__35119;
    wire N__35114;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35106;
    wire N__35103;
    wire N__35100;
    wire N__35097;
    wire N__35090;
    wire N__35087;
    wire N__35084;
    wire N__35081;
    wire N__35078;
    wire N__35075;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35042;
    wire N__35039;
    wire N__35036;
    wire N__35033;
    wire N__35030;
    wire N__35027;
    wire N__35024;
    wire N__35021;
    wire N__35018;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35006;
    wire N__35003;
    wire N__35000;
    wire N__34997;
    wire N__34994;
    wire N__34991;
    wire N__34988;
    wire N__34985;
    wire N__34982;
    wire N__34979;
    wire N__34976;
    wire N__34973;
    wire N__34970;
    wire N__34967;
    wire N__34964;
    wire N__34961;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34946;
    wire N__34943;
    wire N__34940;
    wire N__34937;
    wire N__34934;
    wire N__34931;
    wire N__34928;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34907;
    wire N__34904;
    wire N__34901;
    wire N__34898;
    wire N__34895;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34880;
    wire N__34877;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34865;
    wire N__34862;
    wire N__34859;
    wire N__34856;
    wire N__34855;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34841;
    wire N__34838;
    wire N__34835;
    wire N__34832;
    wire N__34829;
    wire N__34826;
    wire N__34823;
    wire N__34820;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34805;
    wire N__34802;
    wire N__34799;
    wire N__34798;
    wire N__34795;
    wire N__34792;
    wire N__34789;
    wire N__34784;
    wire N__34781;
    wire N__34778;
    wire N__34775;
    wire N__34772;
    wire N__34771;
    wire N__34768;
    wire N__34767;
    wire N__34764;
    wire N__34761;
    wire N__34758;
    wire N__34751;
    wire N__34748;
    wire N__34745;
    wire N__34742;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34724;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34708;
    wire N__34705;
    wire N__34702;
    wire N__34699;
    wire N__34694;
    wire N__34691;
    wire N__34688;
    wire N__34685;
    wire N__34682;
    wire N__34679;
    wire N__34676;
    wire N__34675;
    wire N__34672;
    wire N__34669;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34622;
    wire N__34619;
    wire N__34616;
    wire N__34613;
    wire N__34612;
    wire N__34609;
    wire N__34606;
    wire N__34603;
    wire N__34598;
    wire N__34595;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34585;
    wire N__34582;
    wire N__34579;
    wire N__34576;
    wire N__34571;
    wire N__34568;
    wire N__34565;
    wire N__34562;
    wire N__34559;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34549;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34532;
    wire N__34529;
    wire N__34526;
    wire N__34523;
    wire N__34522;
    wire N__34519;
    wire N__34516;
    wire N__34513;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34499;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34481;
    wire N__34478;
    wire N__34475;
    wire N__34472;
    wire N__34469;
    wire N__34466;
    wire N__34463;
    wire N__34462;
    wire N__34459;
    wire N__34456;
    wire N__34451;
    wire N__34448;
    wire N__34445;
    wire N__34442;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34430;
    wire N__34427;
    wire N__34426;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34412;
    wire N__34409;
    wire N__34406;
    wire N__34403;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34391;
    wire N__34388;
    wire N__34385;
    wire N__34382;
    wire N__34379;
    wire N__34376;
    wire N__34373;
    wire N__34370;
    wire N__34367;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34357;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34343;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34331;
    wire N__34328;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34318;
    wire N__34315;
    wire N__34312;
    wire N__34309;
    wire N__34304;
    wire N__34301;
    wire N__34298;
    wire N__34295;
    wire N__34294;
    wire N__34291;
    wire N__34288;
    wire N__34283;
    wire N__34280;
    wire N__34277;
    wire N__34274;
    wire N__34271;
    wire N__34268;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34256;
    wire N__34253;
    wire N__34250;
    wire N__34249;
    wire N__34246;
    wire N__34243;
    wire N__34240;
    wire N__34235;
    wire N__34232;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34222;
    wire N__34221;
    wire N__34220;
    wire N__34217;
    wire N__34214;
    wire N__34211;
    wire N__34208;
    wire N__34199;
    wire N__34196;
    wire N__34193;
    wire N__34192;
    wire N__34191;
    wire N__34190;
    wire N__34187;
    wire N__34184;
    wire N__34181;
    wire N__34178;
    wire N__34177;
    wire N__34174;
    wire N__34171;
    wire N__34170;
    wire N__34169;
    wire N__34166;
    wire N__34163;
    wire N__34160;
    wire N__34157;
    wire N__34154;
    wire N__34149;
    wire N__34136;
    wire N__34133;
    wire N__34130;
    wire N__34127;
    wire N__34124;
    wire N__34121;
    wire N__34120;
    wire N__34117;
    wire N__34114;
    wire N__34111;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34101;
    wire N__34094;
    wire N__34091;
    wire N__34088;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34063;
    wire N__34058;
    wire N__34055;
    wire N__34052;
    wire N__34051;
    wire N__34050;
    wire N__34049;
    wire N__34046;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34028;
    wire N__34027;
    wire N__34026;
    wire N__34025;
    wire N__34022;
    wire N__34019;
    wire N__34014;
    wire N__34007;
    wire N__34004;
    wire N__34003;
    wire N__34002;
    wire N__34001;
    wire N__34000;
    wire N__33999;
    wire N__33998;
    wire N__33997;
    wire N__33996;
    wire N__33995;
    wire N__33994;
    wire N__33993;
    wire N__33992;
    wire N__33991;
    wire N__33988;
    wire N__33983;
    wire N__33980;
    wire N__33973;
    wire N__33966;
    wire N__33957;
    wire N__33954;
    wire N__33941;
    wire N__33938;
    wire N__33935;
    wire N__33932;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33887;
    wire N__33884;
    wire N__33881;
    wire N__33878;
    wire N__33875;
    wire N__33872;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33851;
    wire N__33848;
    wire N__33845;
    wire N__33842;
    wire N__33839;
    wire N__33836;
    wire N__33833;
    wire N__33830;
    wire N__33827;
    wire N__33824;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33816;
    wire N__33813;
    wire N__33810;
    wire N__33807;
    wire N__33800;
    wire N__33797;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33773;
    wire N__33772;
    wire N__33771;
    wire N__33770;
    wire N__33769;
    wire N__33768;
    wire N__33755;
    wire N__33752;
    wire N__33749;
    wire N__33748;
    wire N__33747;
    wire N__33746;
    wire N__33743;
    wire N__33740;
    wire N__33735;
    wire N__33732;
    wire N__33727;
    wire N__33722;
    wire N__33719;
    wire N__33716;
    wire N__33715;
    wire N__33714;
    wire N__33711;
    wire N__33708;
    wire N__33705;
    wire N__33702;
    wire N__33699;
    wire N__33696;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33635;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33620;
    wire N__33617;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33587;
    wire N__33584;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33572;
    wire N__33569;
    wire N__33566;
    wire N__33563;
    wire N__33560;
    wire N__33557;
    wire N__33554;
    wire N__33553;
    wire N__33548;
    wire N__33545;
    wire N__33542;
    wire N__33539;
    wire N__33536;
    wire N__33533;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33521;
    wire N__33518;
    wire N__33515;
    wire N__33512;
    wire N__33509;
    wire N__33506;
    wire N__33503;
    wire N__33500;
    wire N__33497;
    wire N__33494;
    wire N__33491;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33467;
    wire N__33464;
    wire N__33461;
    wire N__33458;
    wire N__33455;
    wire N__33452;
    wire N__33449;
    wire N__33446;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33434;
    wire N__33431;
    wire N__33428;
    wire N__33425;
    wire N__33422;
    wire N__33421;
    wire N__33418;
    wire N__33417;
    wire N__33414;
    wire N__33411;
    wire N__33410;
    wire N__33407;
    wire N__33404;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33386;
    wire N__33385;
    wire N__33384;
    wire N__33377;
    wire N__33374;
    wire N__33373;
    wire N__33368;
    wire N__33367;
    wire N__33364;
    wire N__33361;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33341;
    wire N__33340;
    wire N__33339;
    wire N__33336;
    wire N__33333;
    wire N__33330;
    wire N__33323;
    wire N__33320;
    wire N__33317;
    wire N__33314;
    wire N__33311;
    wire N__33310;
    wire N__33309;
    wire N__33306;
    wire N__33301;
    wire N__33296;
    wire N__33293;
    wire N__33290;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33278;
    wire N__33277;
    wire N__33276;
    wire N__33273;
    wire N__33270;
    wire N__33267;
    wire N__33264;
    wire N__33263;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33245;
    wire N__33244;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33234;
    wire N__33233;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33219;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33203;
    wire N__33200;
    wire N__33199;
    wire N__33198;
    wire N__33197;
    wire N__33194;
    wire N__33191;
    wire N__33186;
    wire N__33179;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33167;
    wire N__33164;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33152;
    wire N__33149;
    wire N__33146;
    wire N__33143;
    wire N__33140;
    wire N__33137;
    wire N__33136;
    wire N__33135;
    wire N__33134;
    wire N__33133;
    wire N__33132;
    wire N__33131;
    wire N__33130;
    wire N__33129;
    wire N__33128;
    wire N__33127;
    wire N__33126;
    wire N__33125;
    wire N__33122;
    wire N__33117;
    wire N__33116;
    wire N__33113;
    wire N__33112;
    wire N__33111;
    wire N__33110;
    wire N__33109;
    wire N__33106;
    wire N__33105;
    wire N__33104;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33090;
    wire N__33089;
    wire N__33088;
    wire N__33085;
    wire N__33084;
    wire N__33081;
    wire N__33080;
    wire N__33077;
    wire N__33076;
    wire N__33075;
    wire N__33074;
    wire N__33073;
    wire N__33070;
    wire N__33069;
    wire N__33068;
    wire N__33067;
    wire N__33066;
    wire N__33065;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33050;
    wire N__33049;
    wire N__33048;
    wire N__33047;
    wire N__33046;
    wire N__33043;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33011;
    wire N__33008;
    wire N__32993;
    wire N__32986;
    wire N__32983;
    wire N__32982;
    wire N__32979;
    wire N__32978;
    wire N__32975;
    wire N__32974;
    wire N__32965;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32950;
    wire N__32949;
    wire N__32948;
    wire N__32947;
    wire N__32946;
    wire N__32945;
    wire N__32944;
    wire N__32943;
    wire N__32938;
    wire N__32927;
    wire N__32924;
    wire N__32911;
    wire N__32904;
    wire N__32899;
    wire N__32882;
    wire N__32877;
    wire N__32872;
    wire N__32869;
    wire N__32858;
    wire N__32857;
    wire N__32854;
    wire N__32853;
    wire N__32850;
    wire N__32843;
    wire N__32840;
    wire N__32837;
    wire N__32834;
    wire N__32831;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32823;
    wire N__32822;
    wire N__32817;
    wire N__32814;
    wire N__32811;
    wire N__32808;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32794;
    wire N__32791;
    wire N__32788;
    wire N__32785;
    wire N__32782;
    wire N__32779;
    wire N__32774;
    wire N__32771;
    wire N__32768;
    wire N__32765;
    wire N__32764;
    wire N__32763;
    wire N__32760;
    wire N__32755;
    wire N__32754;
    wire N__32753;
    wire N__32748;
    wire N__32743;
    wire N__32738;
    wire N__32735;
    wire N__32734;
    wire N__32731;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32721;
    wire N__32720;
    wire N__32717;
    wire N__32712;
    wire N__32709;
    wire N__32706;
    wire N__32699;
    wire N__32696;
    wire N__32695;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32674;
    wire N__32671;
    wire N__32670;
    wire N__32669;
    wire N__32668;
    wire N__32665;
    wire N__32662;
    wire N__32655;
    wire N__32648;
    wire N__32645;
    wire N__32642;
    wire N__32639;
    wire N__32636;
    wire N__32633;
    wire N__32630;
    wire N__32627;
    wire N__32624;
    wire N__32621;
    wire N__32618;
    wire N__32615;
    wire N__32612;
    wire N__32611;
    wire N__32610;
    wire N__32605;
    wire N__32602;
    wire N__32597;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32587;
    wire N__32582;
    wire N__32579;
    wire N__32578;
    wire N__32577;
    wire N__32576;
    wire N__32575;
    wire N__32574;
    wire N__32571;
    wire N__32568;
    wire N__32567;
    wire N__32564;
    wire N__32561;
    wire N__32560;
    wire N__32559;
    wire N__32558;
    wire N__32555;
    wire N__32552;
    wire N__32551;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32534;
    wire N__32523;
    wire N__32518;
    wire N__32507;
    wire N__32506;
    wire N__32505;
    wire N__32498;
    wire N__32495;
    wire N__32494;
    wire N__32491;
    wire N__32488;
    wire N__32485;
    wire N__32484;
    wire N__32479;
    wire N__32476;
    wire N__32471;
    wire N__32470;
    wire N__32469;
    wire N__32466;
    wire N__32463;
    wire N__32462;
    wire N__32459;
    wire N__32454;
    wire N__32451;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32428;
    wire N__32425;
    wire N__32424;
    wire N__32423;
    wire N__32420;
    wire N__32417;
    wire N__32412;
    wire N__32407;
    wire N__32402;
    wire N__32399;
    wire N__32396;
    wire N__32393;
    wire N__32390;
    wire N__32387;
    wire N__32386;
    wire N__32383;
    wire N__32382;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32363;
    wire N__32362;
    wire N__32359;
    wire N__32356;
    wire N__32351;
    wire N__32348;
    wire N__32347;
    wire N__32346;
    wire N__32343;
    wire N__32340;
    wire N__32337;
    wire N__32330;
    wire N__32327;
    wire N__32326;
    wire N__32325;
    wire N__32322;
    wire N__32317;
    wire N__32312;
    wire N__32309;
    wire N__32308;
    wire N__32307;
    wire N__32304;
    wire N__32299;
    wire N__32294;
    wire N__32291;
    wire N__32290;
    wire N__32287;
    wire N__32284;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32274;
    wire N__32271;
    wire N__32264;
    wire N__32261;
    wire N__32260;
    wire N__32257;
    wire N__32254;
    wire N__32253;
    wire N__32250;
    wire N__32247;
    wire N__32244;
    wire N__32241;
    wire N__32234;
    wire N__32231;
    wire N__32228;
    wire N__32227;
    wire N__32226;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32210;
    wire N__32207;
    wire N__32204;
    wire N__32203;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32193;
    wire N__32186;
    wire N__32183;
    wire N__32182;
    wire N__32179;
    wire N__32176;
    wire N__32171;
    wire N__32168;
    wire N__32167;
    wire N__32166;
    wire N__32165;
    wire N__32164;
    wire N__32163;
    wire N__32162;
    wire N__32161;
    wire N__32160;
    wire N__32159;
    wire N__32158;
    wire N__32157;
    wire N__32156;
    wire N__32155;
    wire N__32154;
    wire N__32153;
    wire N__32152;
    wire N__32151;
    wire N__32150;
    wire N__32149;
    wire N__32148;
    wire N__32147;
    wire N__32146;
    wire N__32145;
    wire N__32144;
    wire N__32143;
    wire N__32142;
    wire N__32141;
    wire N__32140;
    wire N__32139;
    wire N__32130;
    wire N__32125;
    wire N__32116;
    wire N__32107;
    wire N__32098;
    wire N__32089;
    wire N__32080;
    wire N__32071;
    wire N__32068;
    wire N__32057;
    wire N__32052;
    wire N__32047;
    wire N__32044;
    wire N__32039;
    wire N__32036;
    wire N__32035;
    wire N__32032;
    wire N__32029;
    wire N__32024;
    wire N__32021;
    wire N__32020;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32003;
    wire N__32000;
    wire N__31999;
    wire N__31998;
    wire N__31995;
    wire N__31990;
    wire N__31985;
    wire N__31982;
    wire N__31981;
    wire N__31980;
    wire N__31977;
    wire N__31972;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31934;
    wire N__31931;
    wire N__31930;
    wire N__31927;
    wire N__31924;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31904;
    wire N__31901;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31884;
    wire N__31881;
    wire N__31874;
    wire N__31871;
    wire N__31868;
    wire N__31867;
    wire N__31866;
    wire N__31863;
    wire N__31860;
    wire N__31857;
    wire N__31850;
    wire N__31847;
    wire N__31844;
    wire N__31843;
    wire N__31842;
    wire N__31839;
    wire N__31836;
    wire N__31833;
    wire N__31826;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31816;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31799;
    wire N__31796;
    wire N__31795;
    wire N__31794;
    wire N__31791;
    wire N__31786;
    wire N__31781;
    wire N__31778;
    wire N__31777;
    wire N__31776;
    wire N__31773;
    wire N__31768;
    wire N__31763;
    wire N__31760;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31733;
    wire N__31730;
    wire N__31729;
    wire N__31726;
    wire N__31723;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31696;
    wire N__31695;
    wire N__31692;
    wire N__31689;
    wire N__31686;
    wire N__31679;
    wire N__31676;
    wire N__31673;
    wire N__31672;
    wire N__31671;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31648;
    wire N__31647;
    wire N__31644;
    wire N__31641;
    wire N__31638;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31596;
    wire N__31593;
    wire N__31590;
    wire N__31587;
    wire N__31580;
    wire N__31577;
    wire N__31574;
    wire N__31573;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31549;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31532;
    wire N__31529;
    wire N__31526;
    wire N__31525;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31508;
    wire N__31507;
    wire N__31504;
    wire N__31503;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31489;
    wire N__31486;
    wire N__31481;
    wire N__31480;
    wire N__31477;
    wire N__31476;
    wire N__31475;
    wire N__31466;
    wire N__31463;
    wire N__31460;
    wire N__31459;
    wire N__31456;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31448;
    wire N__31445;
    wire N__31442;
    wire N__31439;
    wire N__31436;
    wire N__31431;
    wire N__31428;
    wire N__31423;
    wire N__31418;
    wire N__31415;
    wire N__31412;
    wire N__31409;
    wire N__31408;
    wire N__31405;
    wire N__31402;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31391;
    wire N__31390;
    wire N__31387;
    wire N__31384;
    wire N__31381;
    wire N__31376;
    wire N__31369;
    wire N__31366;
    wire N__31361;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31338;
    wire N__31335;
    wire N__31334;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31315;
    wire N__31312;
    wire N__31307;
    wire N__31304;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31294;
    wire N__31291;
    wire N__31288;
    wire N__31287;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31271;
    wire N__31270;
    wire N__31269;
    wire N__31262;
    wire N__31259;
    wire N__31256;
    wire N__31255;
    wire N__31254;
    wire N__31253;
    wire N__31252;
    wire N__31249;
    wire N__31242;
    wire N__31239;
    wire N__31238;
    wire N__31235;
    wire N__31232;
    wire N__31229;
    wire N__31226;
    wire N__31221;
    wire N__31216;
    wire N__31211;
    wire N__31208;
    wire N__31205;
    wire N__31202;
    wire N__31199;
    wire N__31196;
    wire N__31195;
    wire N__31194;
    wire N__31191;
    wire N__31186;
    wire N__31181;
    wire N__31178;
    wire N__31175;
    wire N__31172;
    wire N__31169;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31142;
    wire N__31139;
    wire N__31136;
    wire N__31133;
    wire N__31130;
    wire N__31127;
    wire N__31126;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31114;
    wire N__31109;
    wire N__31106;
    wire N__31103;
    wire N__31102;
    wire N__31101;
    wire N__31094;
    wire N__31091;
    wire N__31088;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31078;
    wire N__31075;
    wire N__31074;
    wire N__31073;
    wire N__31070;
    wire N__31067;
    wire N__31064;
    wire N__31061;
    wire N__31056;
    wire N__31053;
    wire N__31046;
    wire N__31043;
    wire N__31040;
    wire N__31037;
    wire N__31034;
    wire N__31031;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31019;
    wire N__31016;
    wire N__31015;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31003;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30986;
    wire N__30985;
    wire N__30982;
    wire N__30979;
    wire N__30974;
    wire N__30971;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30961;
    wire N__30958;
    wire N__30955;
    wire N__30950;
    wire N__30947;
    wire N__30944;
    wire N__30941;
    wire N__30940;
    wire N__30937;
    wire N__30934;
    wire N__30929;
    wire N__30926;
    wire N__30923;
    wire N__30920;
    wire N__30919;
    wire N__30916;
    wire N__30913;
    wire N__30908;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30895;
    wire N__30892;
    wire N__30889;
    wire N__30884;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30874;
    wire N__30871;
    wire N__30868;
    wire N__30863;
    wire N__30860;
    wire N__30857;
    wire N__30856;
    wire N__30855;
    wire N__30854;
    wire N__30851;
    wire N__30850;
    wire N__30845;
    wire N__30842;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30830;
    wire N__30827;
    wire N__30824;
    wire N__30821;
    wire N__30816;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30800;
    wire N__30799;
    wire N__30796;
    wire N__30795;
    wire N__30792;
    wire N__30791;
    wire N__30790;
    wire N__30787;
    wire N__30782;
    wire N__30777;
    wire N__30774;
    wire N__30767;
    wire N__30764;
    wire N__30763;
    wire N__30760;
    wire N__30757;
    wire N__30754;
    wire N__30751;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30727;
    wire N__30724;
    wire N__30721;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30711;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30695;
    wire N__30692;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30684;
    wire N__30681;
    wire N__30678;
    wire N__30675;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30661;
    wire N__30658;
    wire N__30657;
    wire N__30654;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30637;
    wire N__30632;
    wire N__30629;
    wire N__30626;
    wire N__30623;
    wire N__30622;
    wire N__30619;
    wire N__30616;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30598;
    wire N__30595;
    wire N__30592;
    wire N__30587;
    wire N__30584;
    wire N__30581;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30569;
    wire N__30566;
    wire N__30563;
    wire N__30560;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30550;
    wire N__30547;
    wire N__30542;
    wire N__30539;
    wire N__30536;
    wire N__30533;
    wire N__30530;
    wire N__30529;
    wire N__30528;
    wire N__30525;
    wire N__30520;
    wire N__30515;
    wire N__30512;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30502;
    wire N__30501;
    wire N__30498;
    wire N__30493;
    wire N__30488;
    wire N__30485;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30473;
    wire N__30472;
    wire N__30471;
    wire N__30470;
    wire N__30467;
    wire N__30464;
    wire N__30461;
    wire N__30458;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30430;
    wire N__30427;
    wire N__30422;
    wire N__30419;
    wire N__30416;
    wire N__30413;
    wire N__30410;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30398;
    wire N__30395;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30385;
    wire N__30382;
    wire N__30379;
    wire N__30374;
    wire N__30371;
    wire N__30368;
    wire N__30365;
    wire N__30362;
    wire N__30361;
    wire N__30358;
    wire N__30355;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30340;
    wire N__30337;
    wire N__30336;
    wire N__30335;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30320;
    wire N__30315;
    wire N__30308;
    wire N__30305;
    wire N__30302;
    wire N__30301;
    wire N__30300;
    wire N__30297;
    wire N__30294;
    wire N__30291;
    wire N__30284;
    wire N__30281;
    wire N__30280;
    wire N__30277;
    wire N__30274;
    wire N__30271;
    wire N__30270;
    wire N__30267;
    wire N__30266;
    wire N__30265;
    wire N__30264;
    wire N__30263;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30247;
    wire N__30244;
    wire N__30233;
    wire N__30232;
    wire N__30231;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30206;
    wire N__30205;
    wire N__30204;
    wire N__30203;
    wire N__30202;
    wire N__30201;
    wire N__30200;
    wire N__30197;
    wire N__30194;
    wire N__30187;
    wire N__30186;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30174;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30157;
    wire N__30146;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30130;
    wire N__30125;
    wire N__30122;
    wire N__30121;
    wire N__30120;
    wire N__30117;
    wire N__30112;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30098;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30074;
    wire N__30073;
    wire N__30070;
    wire N__30067;
    wire N__30062;
    wire N__30059;
    wire N__30058;
    wire N__30057;
    wire N__30052;
    wire N__30049;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30028;
    wire N__30025;
    wire N__30022;
    wire N__30019;
    wire N__30014;
    wire N__30011;
    wire N__30008;
    wire N__30005;
    wire N__30002;
    wire N__29999;
    wire N__29996;
    wire N__29993;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29966;
    wire N__29963;
    wire N__29960;
    wire N__29957;
    wire N__29956;
    wire N__29953;
    wire N__29950;
    wire N__29947;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29933;
    wire N__29930;
    wire N__29929;
    wire N__29926;
    wire N__29925;
    wire N__29922;
    wire N__29919;
    wire N__29916;
    wire N__29913;
    wire N__29910;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29896;
    wire N__29893;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29879;
    wire N__29876;
    wire N__29875;
    wire N__29874;
    wire N__29871;
    wire N__29870;
    wire N__29865;
    wire N__29862;
    wire N__29859;
    wire N__29856;
    wire N__29853;
    wire N__29846;
    wire N__29843;
    wire N__29840;
    wire N__29837;
    wire N__29834;
    wire N__29833;
    wire N__29830;
    wire N__29827;
    wire N__29824;
    wire N__29819;
    wire N__29816;
    wire N__29813;
    wire N__29810;
    wire N__29807;
    wire N__29804;
    wire N__29801;
    wire N__29798;
    wire N__29795;
    wire N__29794;
    wire N__29791;
    wire N__29788;
    wire N__29785;
    wire N__29780;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29765;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29734;
    wire N__29731;
    wire N__29728;
    wire N__29725;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29690;
    wire N__29687;
    wire N__29684;
    wire N__29681;
    wire N__29678;
    wire N__29675;
    wire N__29672;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29657;
    wire N__29654;
    wire N__29651;
    wire N__29648;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29638;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29602;
    wire N__29599;
    wire N__29596;
    wire N__29593;
    wire N__29588;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29566;
    wire N__29563;
    wire N__29560;
    wire N__29557;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29540;
    wire N__29537;
    wire N__29536;
    wire N__29533;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29495;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29480;
    wire N__29477;
    wire N__29474;
    wire N__29471;
    wire N__29468;
    wire N__29467;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29444;
    wire N__29441;
    wire N__29438;
    wire N__29435;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29408;
    wire N__29407;
    wire N__29404;
    wire N__29401;
    wire N__29398;
    wire N__29393;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29359;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29339;
    wire N__29336;
    wire N__29333;
    wire N__29330;
    wire N__29327;
    wire N__29324;
    wire N__29321;
    wire N__29320;
    wire N__29317;
    wire N__29314;
    wire N__29309;
    wire N__29308;
    wire N__29305;
    wire N__29304;
    wire N__29301;
    wire N__29300;
    wire N__29299;
    wire N__29298;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29287;
    wire N__29286;
    wire N__29285;
    wire N__29284;
    wire N__29283;
    wire N__29282;
    wire N__29281;
    wire N__29280;
    wire N__29279;
    wire N__29278;
    wire N__29277;
    wire N__29276;
    wire N__29275;
    wire N__29274;
    wire N__29273;
    wire N__29268;
    wire N__29263;
    wire N__29258;
    wire N__29255;
    wire N__29246;
    wire N__29237;
    wire N__29230;
    wire N__29221;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29199;
    wire N__29196;
    wire N__29191;
    wire N__29188;
    wire N__29183;
    wire N__29180;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29160;
    wire N__29157;
    wire N__29154;
    wire N__29151;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29135;
    wire N__29132;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29120;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29108;
    wire N__29105;
    wire N__29104;
    wire N__29101;
    wire N__29098;
    wire N__29097;
    wire N__29092;
    wire N__29089;
    wire N__29084;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29072;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29064;
    wire N__29059;
    wire N__29056;
    wire N__29051;
    wire N__29050;
    wire N__29045;
    wire N__29042;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29024;
    wire N__29021;
    wire N__29018;
    wire N__29015;
    wire N__29012;
    wire N__29009;
    wire N__29006;
    wire N__29003;
    wire N__29000;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28984;
    wire N__28983;
    wire N__28978;
    wire N__28975;
    wire N__28970;
    wire N__28969;
    wire N__28966;
    wire N__28965;
    wire N__28964;
    wire N__28959;
    wire N__28956;
    wire N__28953;
    wire N__28946;
    wire N__28943;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28931;
    wire N__28928;
    wire N__28927;
    wire N__28926;
    wire N__28921;
    wire N__28918;
    wire N__28913;
    wire N__28912;
    wire N__28909;
    wire N__28906;
    wire N__28901;
    wire N__28898;
    wire N__28897;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28874;
    wire N__28873;
    wire N__28872;
    wire N__28871;
    wire N__28870;
    wire N__28869;
    wire N__28868;
    wire N__28867;
    wire N__28866;
    wire N__28863;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28830;
    wire N__28829;
    wire N__28828;
    wire N__28825;
    wire N__28824;
    wire N__28823;
    wire N__28822;
    wire N__28821;
    wire N__28820;
    wire N__28819;
    wire N__28818;
    wire N__28817;
    wire N__28816;
    wire N__28815;
    wire N__28814;
    wire N__28813;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28794;
    wire N__28791;
    wire N__28784;
    wire N__28781;
    wire N__28772;
    wire N__28763;
    wire N__28758;
    wire N__28753;
    wire N__28748;
    wire N__28733;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28721;
    wire N__28720;
    wire N__28717;
    wire N__28714;
    wire N__28713;
    wire N__28712;
    wire N__28711;
    wire N__28708;
    wire N__28703;
    wire N__28698;
    wire N__28691;
    wire N__28690;
    wire N__28689;
    wire N__28686;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28645;
    wire N__28644;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28634;
    wire N__28631;
    wire N__28628;
    wire N__28623;
    wire N__28616;
    wire N__28613;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28603;
    wire N__28598;
    wire N__28595;
    wire N__28594;
    wire N__28591;
    wire N__28588;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28571;
    wire N__28568;
    wire N__28565;
    wire N__28564;
    wire N__28561;
    wire N__28558;
    wire N__28553;
    wire N__28552;
    wire N__28549;
    wire N__28546;
    wire N__28543;
    wire N__28538;
    wire N__28535;
    wire N__28532;
    wire N__28529;
    wire N__28526;
    wire N__28523;
    wire N__28520;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28508;
    wire N__28507;
    wire N__28504;
    wire N__28501;
    wire N__28496;
    wire N__28495;
    wire N__28494;
    wire N__28491;
    wire N__28490;
    wire N__28489;
    wire N__28486;
    wire N__28485;
    wire N__28482;
    wire N__28481;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28447;
    wire N__28444;
    wire N__28439;
    wire N__28436;
    wire N__28433;
    wire N__28426;
    wire N__28421;
    wire N__28412;
    wire N__28411;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28394;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28382;
    wire N__28379;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28367;
    wire N__28364;
    wire N__28361;
    wire N__28358;
    wire N__28355;
    wire N__28354;
    wire N__28351;
    wire N__28348;
    wire N__28343;
    wire N__28340;
    wire N__28339;
    wire N__28338;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28320;
    wire N__28313;
    wire N__28312;
    wire N__28311;
    wire N__28310;
    wire N__28309;
    wire N__28308;
    wire N__28307;
    wire N__28306;
    wire N__28299;
    wire N__28298;
    wire N__28295;
    wire N__28294;
    wire N__28293;
    wire N__28292;
    wire N__28291;
    wire N__28290;
    wire N__28281;
    wire N__28278;
    wire N__28273;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28247;
    wire N__28246;
    wire N__28245;
    wire N__28244;
    wire N__28243;
    wire N__28242;
    wire N__28241;
    wire N__28240;
    wire N__28239;
    wire N__28238;
    wire N__28237;
    wire N__28236;
    wire N__28235;
    wire N__28234;
    wire N__28233;
    wire N__28232;
    wire N__28231;
    wire N__28230;
    wire N__28229;
    wire N__28228;
    wire N__28227;
    wire N__28226;
    wire N__28215;
    wire N__28212;
    wire N__28201;
    wire N__28186;
    wire N__28177;
    wire N__28176;
    wire N__28175;
    wire N__28174;
    wire N__28173;
    wire N__28172;
    wire N__28171;
    wire N__28170;
    wire N__28169;
    wire N__28168;
    wire N__28167;
    wire N__28166;
    wire N__28165;
    wire N__28164;
    wire N__28163;
    wire N__28160;
    wire N__28157;
    wire N__28150;
    wire N__28147;
    wire N__28140;
    wire N__28127;
    wire N__28118;
    wire N__28115;
    wire N__28106;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28090;
    wire N__28087;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28070;
    wire N__28069;
    wire N__28068;
    wire N__28067;
    wire N__28066;
    wire N__28065;
    wire N__28064;
    wire N__28063;
    wire N__28062;
    wire N__28061;
    wire N__28060;
    wire N__28057;
    wire N__28056;
    wire N__28049;
    wire N__28046;
    wire N__28039;
    wire N__28028;
    wire N__28019;
    wire N__28018;
    wire N__28015;
    wire N__28012;
    wire N__28007;
    wire N__28006;
    wire N__28003;
    wire N__28000;
    wire N__27995;
    wire N__27992;
    wire N__27991;
    wire N__27988;
    wire N__27985;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27965;
    wire N__27964;
    wire N__27961;
    wire N__27960;
    wire N__27959;
    wire N__27958;
    wire N__27957;
    wire N__27954;
    wire N__27947;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27939;
    wire N__27936;
    wire N__27933;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27917;
    wire N__27908;
    wire N__27907;
    wire N__27904;
    wire N__27901;
    wire N__27898;
    wire N__27897;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27885;
    wire N__27878;
    wire N__27875;
    wire N__27874;
    wire N__27873;
    wire N__27872;
    wire N__27871;
    wire N__27870;
    wire N__27869;
    wire N__27868;
    wire N__27867;
    wire N__27866;
    wire N__27865;
    wire N__27864;
    wire N__27863;
    wire N__27862;
    wire N__27861;
    wire N__27858;
    wire N__27857;
    wire N__27856;
    wire N__27855;
    wire N__27854;
    wire N__27853;
    wire N__27852;
    wire N__27851;
    wire N__27850;
    wire N__27841;
    wire N__27830;
    wire N__27819;
    wire N__27816;
    wire N__27815;
    wire N__27812;
    wire N__27811;
    wire N__27810;
    wire N__27807;
    wire N__27794;
    wire N__27791;
    wire N__27784;
    wire N__27777;
    wire N__27774;
    wire N__27761;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27753;
    wire N__27752;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27723;
    wire N__27718;
    wire N__27707;
    wire N__27706;
    wire N__27703;
    wire N__27702;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27692;
    wire N__27689;
    wire N__27680;
    wire N__27679;
    wire N__27678;
    wire N__27677;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27650;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27632;
    wire N__27629;
    wire N__27628;
    wire N__27623;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27598;
    wire N__27595;
    wire N__27592;
    wire N__27587;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27579;
    wire N__27576;
    wire N__27573;
    wire N__27570;
    wire N__27563;
    wire N__27560;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27548;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27529;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27511;
    wire N__27510;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27488;
    wire N__27479;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27467;
    wire N__27464;
    wire N__27461;
    wire N__27460;
    wire N__27459;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27449;
    wire N__27446;
    wire N__27443;
    wire N__27440;
    wire N__27435;
    wire N__27432;
    wire N__27429;
    wire N__27426;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27407;
    wire N__27404;
    wire N__27403;
    wire N__27402;
    wire N__27401;
    wire N__27400;
    wire N__27399;
    wire N__27398;
    wire N__27397;
    wire N__27396;
    wire N__27395;
    wire N__27392;
    wire N__27391;
    wire N__27390;
    wire N__27389;
    wire N__27388;
    wire N__27387;
    wire N__27380;
    wire N__27379;
    wire N__27378;
    wire N__27377;
    wire N__27376;
    wire N__27375;
    wire N__27374;
    wire N__27373;
    wire N__27372;
    wire N__27371;
    wire N__27370;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27342;
    wire N__27339;
    wire N__27328;
    wire N__27327;
    wire N__27326;
    wire N__27325;
    wire N__27324;
    wire N__27323;
    wire N__27322;
    wire N__27311;
    wire N__27310;
    wire N__27305;
    wire N__27302;
    wire N__27295;
    wire N__27282;
    wire N__27279;
    wire N__27276;
    wire N__27273;
    wire N__27268;
    wire N__27257;
    wire N__27256;
    wire N__27255;
    wire N__27254;
    wire N__27253;
    wire N__27252;
    wire N__27251;
    wire N__27250;
    wire N__27249;
    wire N__27248;
    wire N__27247;
    wire N__27244;
    wire N__27241;
    wire N__27240;
    wire N__27239;
    wire N__27238;
    wire N__27225;
    wire N__27224;
    wire N__27223;
    wire N__27222;
    wire N__27221;
    wire N__27210;
    wire N__27203;
    wire N__27202;
    wire N__27201;
    wire N__27200;
    wire N__27199;
    wire N__27198;
    wire N__27197;
    wire N__27196;
    wire N__27195;
    wire N__27194;
    wire N__27193;
    wire N__27190;
    wire N__27181;
    wire N__27178;
    wire N__27175;
    wire N__27164;
    wire N__27153;
    wire N__27150;
    wire N__27143;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27122;
    wire N__27119;
    wire N__27118;
    wire N__27117;
    wire N__27116;
    wire N__27115;
    wire N__27114;
    wire N__27113;
    wire N__27112;
    wire N__27111;
    wire N__27110;
    wire N__27109;
    wire N__27106;
    wire N__27103;
    wire N__27100;
    wire N__27099;
    wire N__27098;
    wire N__27095;
    wire N__27094;
    wire N__27093;
    wire N__27092;
    wire N__27091;
    wire N__27090;
    wire N__27089;
    wire N__27088;
    wire N__27085;
    wire N__27084;
    wire N__27083;
    wire N__27082;
    wire N__27081;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27070;
    wire N__27069;
    wire N__27056;
    wire N__27049;
    wire N__27048;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27037;
    wire N__27036;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27024;
    wire N__27021;
    wire N__27010;
    wire N__27003;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26981;
    wire N__26970;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26942;
    wire N__26939;
    wire N__26938;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26930;
    wire N__26927;
    wire N__26924;
    wire N__26921;
    wire N__26918;
    wire N__26915;
    wire N__26910;
    wire N__26903;
    wire N__26902;
    wire N__26899;
    wire N__26896;
    wire N__26891;
    wire N__26890;
    wire N__26887;
    wire N__26884;
    wire N__26883;
    wire N__26882;
    wire N__26879;
    wire N__26876;
    wire N__26871;
    wire N__26864;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26851;
    wire N__26848;
    wire N__26847;
    wire N__26842;
    wire N__26839;
    wire N__26834;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26822;
    wire N__26819;
    wire N__26816;
    wire N__26815;
    wire N__26812;
    wire N__26811;
    wire N__26808;
    wire N__26805;
    wire N__26804;
    wire N__26803;
    wire N__26800;
    wire N__26797;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26785;
    wire N__26778;
    wire N__26775;
    wire N__26768;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26758;
    wire N__26755;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26729;
    wire N__26726;
    wire N__26723;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26711;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26703;
    wire N__26698;
    wire N__26695;
    wire N__26692;
    wire N__26687;
    wire N__26684;
    wire N__26681;
    wire N__26680;
    wire N__26679;
    wire N__26678;
    wire N__26675;
    wire N__26672;
    wire N__26669;
    wire N__26668;
    wire N__26665;
    wire N__26658;
    wire N__26655;
    wire N__26650;
    wire N__26645;
    wire N__26642;
    wire N__26639;
    wire N__26638;
    wire N__26637;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26615;
    wire N__26612;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26597;
    wire N__26594;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26586;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26571;
    wire N__26564;
    wire N__26563;
    wire N__26560;
    wire N__26559;
    wire N__26556;
    wire N__26553;
    wire N__26550;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26534;
    wire N__26533;
    wire N__26528;
    wire N__26523;
    wire N__26520;
    wire N__26517;
    wire N__26510;
    wire N__26507;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26462;
    wire N__26461;
    wire N__26460;
    wire N__26457;
    wire N__26454;
    wire N__26451;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26433;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26410;
    wire N__26407;
    wire N__26404;
    wire N__26401;
    wire N__26400;
    wire N__26397;
    wire N__26394;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26353;
    wire N__26350;
    wire N__26347;
    wire N__26342;
    wire N__26339;
    wire N__26338;
    wire N__26335;
    wire N__26332;
    wire N__26331;
    wire N__26328;
    wire N__26327;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26312;
    wire N__26309;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26287;
    wire N__26284;
    wire N__26283;
    wire N__26280;
    wire N__26277;
    wire N__26274;
    wire N__26273;
    wire N__26272;
    wire N__26269;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26253;
    wire N__26250;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26212;
    wire N__26209;
    wire N__26206;
    wire N__26203;
    wire N__26202;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26186;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26171;
    wire N__26168;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26150;
    wire N__26149;
    wire N__26146;
    wire N__26143;
    wire N__26142;
    wire N__26139;
    wire N__26138;
    wire N__26135;
    wire N__26134;
    wire N__26131;
    wire N__26128;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26116;
    wire N__26111;
    wire N__26108;
    wire N__26101;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26074;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26064;
    wire N__26061;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26047;
    wire N__26044;
    wire N__26043;
    wire N__26040;
    wire N__26037;
    wire N__26034;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26020;
    wire N__26019;
    wire N__26016;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26000;
    wire N__25997;
    wire N__25996;
    wire N__25995;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25983;
    wire N__25976;
    wire N__25973;
    wire N__25972;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25959;
    wire N__25952;
    wire N__25949;
    wire N__25948;
    wire N__25945;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25935;
    wire N__25930;
    wire N__25925;
    wire N__25922;
    wire N__25921;
    wire N__25920;
    wire N__25917;
    wire N__25914;
    wire N__25911;
    wire N__25908;
    wire N__25901;
    wire N__25898;
    wire N__25897;
    wire N__25894;
    wire N__25893;
    wire N__25890;
    wire N__25887;
    wire N__25884;
    wire N__25877;
    wire N__25874;
    wire N__25873;
    wire N__25872;
    wire N__25871;
    wire N__25870;
    wire N__25869;
    wire N__25868;
    wire N__25867;
    wire N__25866;
    wire N__25865;
    wire N__25856;
    wire N__25851;
    wire N__25842;
    wire N__25835;
    wire N__25832;
    wire N__25831;
    wire N__25828;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25811;
    wire N__25810;
    wire N__25807;
    wire N__25804;
    wire N__25801;
    wire N__25796;
    wire N__25793;
    wire N__25792;
    wire N__25789;
    wire N__25786;
    wire N__25783;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25757;
    wire N__25754;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25739;
    wire N__25736;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25721;
    wire N__25718;
    wire N__25717;
    wire N__25714;
    wire N__25711;
    wire N__25708;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25682;
    wire N__25681;
    wire N__25678;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25661;
    wire N__25658;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25643;
    wire N__25640;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25625;
    wire N__25622;
    wire N__25621;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25607;
    wire N__25604;
    wire N__25603;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25589;
    wire N__25586;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25576;
    wire N__25571;
    wire N__25568;
    wire N__25567;
    wire N__25564;
    wire N__25561;
    wire N__25558;
    wire N__25553;
    wire N__25550;
    wire N__25549;
    wire N__25546;
    wire N__25543;
    wire N__25540;
    wire N__25535;
    wire N__25532;
    wire N__25531;
    wire N__25528;
    wire N__25525;
    wire N__25522;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25487;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25460;
    wire N__25459;
    wire N__25456;
    wire N__25453;
    wire N__25450;
    wire N__25445;
    wire N__25442;
    wire N__25441;
    wire N__25438;
    wire N__25435;
    wire N__25432;
    wire N__25427;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25415;
    wire N__25412;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25117;
    wire N__25112;
    wire N__25109;
    wire N__25108;
    wire N__25105;
    wire N__25102;
    wire N__25097;
    wire N__25094;
    wire N__25093;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25042;
    wire N__25039;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25031;
    wire N__25028;
    wire N__25023;
    wire N__25020;
    wire N__25013;
    wire N__25010;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__25000;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24976;
    wire N__24975;
    wire N__24972;
    wire N__24969;
    wire N__24966;
    wire N__24959;
    wire N__24958;
    wire N__24957;
    wire N__24954;
    wire N__24949;
    wire N__24944;
    wire N__24943;
    wire N__24940;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24914;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24890;
    wire N__24887;
    wire N__24884;
    wire N__24883;
    wire N__24882;
    wire N__24881;
    wire N__24880;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24855;
    wire N__24852;
    wire N__24847;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24826;
    wire N__24823;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24813;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24755;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24662;
    wire N__24659;
    wire N__24656;
    wire N__24653;
    wire N__24650;
    wire N__24647;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24593;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24572;
    wire N__24569;
    wire N__24566;
    wire N__24563;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24476;
    wire N__24473;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24368;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24296;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24281;
    wire N__24278;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24224;
    wire N__24221;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24180;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24168;
    wire N__24167;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24149;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24139;
    wire N__24134;
    wire N__24131;
    wire N__24128;
    wire N__24125;
    wire N__24124;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24112;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24094;
    wire N__24089;
    wire N__24086;
    wire N__24083;
    wire N__24080;
    wire N__24077;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24049;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24039;
    wire N__24038;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24017;
    wire N__24010;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23993;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23980;
    wire N__23977;
    wire N__23974;
    wire N__23973;
    wire N__23970;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23959;
    wire N__23956;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23938;
    wire N__23935;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23878;
    wire N__23875;
    wire N__23872;
    wire N__23869;
    wire N__23868;
    wire N__23867;
    wire N__23866;
    wire N__23861;
    wire N__23856;
    wire N__23853;
    wire N__23846;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23834;
    wire N__23833;
    wire N__23830;
    wire N__23829;
    wire N__23828;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23814;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23777;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23769;
    wire N__23764;
    wire N__23763;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23751;
    wire N__23744;
    wire N__23743;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23732;
    wire N__23727;
    wire N__23724;
    wire N__23721;
    wire N__23714;
    wire N__23713;
    wire N__23712;
    wire N__23709;
    wire N__23708;
    wire N__23707;
    wire N__23704;
    wire N__23701;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23685;
    wire N__23678;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23666;
    wire N__23665;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23655;
    wire N__23652;
    wire N__23645;
    wire N__23644;
    wire N__23641;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23605;
    wire N__23602;
    wire N__23601;
    wire N__23600;
    wire N__23599;
    wire N__23596;
    wire N__23593;
    wire N__23590;
    wire N__23585;
    wire N__23576;
    wire N__23573;
    wire N__23572;
    wire N__23569;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23555;
    wire N__23554;
    wire N__23551;
    wire N__23550;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23538;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23512;
    wire N__23511;
    wire N__23508;
    wire N__23505;
    wire N__23502;
    wire N__23501;
    wire N__23500;
    wire N__23495;
    wire N__23492;
    wire N__23487;
    wire N__23480;
    wire N__23479;
    wire N__23476;
    wire N__23475;
    wire N__23472;
    wire N__23469;
    wire N__23466;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23452;
    wire N__23449;
    wire N__23446;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23428;
    wire N__23427;
    wire N__23424;
    wire N__23421;
    wire N__23418;
    wire N__23417;
    wire N__23416;
    wire N__23413;
    wire N__23410;
    wire N__23407;
    wire N__23402;
    wire N__23397;
    wire N__23392;
    wire N__23387;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23375;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23362;
    wire N__23361;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23347;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23314;
    wire N__23311;
    wire N__23310;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23294;
    wire N__23291;
    wire N__23290;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23266;
    wire N__23263;
    wire N__23256;
    wire N__23253;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23223;
    wire N__23222;
    wire N__23221;
    wire N__23218;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23195;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23187;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23143;
    wire N__23140;
    wire N__23139;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23092;
    wire N__23089;
    wire N__23088;
    wire N__23085;
    wire N__23082;
    wire N__23079;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23065;
    wire N__23062;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23032;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23017;
    wire N__23012;
    wire N__23011;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22994;
    wire N__22991;
    wire N__22990;
    wire N__22989;
    wire N__22986;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22943;
    wire N__22940;
    wire N__22939;
    wire N__22936;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22896;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22862;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22816;
    wire N__22813;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22771;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22755;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22731;
    wire N__22730;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22715;
    wire N__22706;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22695;
    wire N__22690;
    wire N__22687;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22672;
    wire N__22669;
    wire N__22666;
    wire N__22661;
    wire N__22660;
    wire N__22657;
    wire N__22654;
    wire N__22651;
    wire N__22650;
    wire N__22649;
    wire N__22648;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22638;
    wire N__22633;
    wire N__22626;
    wire N__22623;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22558;
    wire N__22555;
    wire N__22554;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22525;
    wire N__22522;
    wire N__22521;
    wire N__22518;
    wire N__22515;
    wire N__22512;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22498;
    wire N__22497;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22475;
    wire N__22472;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22444;
    wire N__22441;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22318;
    wire N__22315;
    wire N__22312;
    wire N__22309;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22298;
    wire N__22297;
    wire N__22294;
    wire N__22289;
    wire N__22284;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21913;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21814;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21799;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21634;
    wire N__21629;
    wire N__21626;
    wire N__21625;
    wire N__21620;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21526;
    wire N__21525;
    wire N__21524;
    wire N__21523;
    wire N__21522;
    wire N__21521;
    wire N__21520;
    wire N__21519;
    wire N__21516;
    wire N__21515;
    wire N__21512;
    wire N__21511;
    wire N__21508;
    wire N__21507;
    wire N__21504;
    wire N__21503;
    wire N__21500;
    wire N__21499;
    wire N__21496;
    wire N__21495;
    wire N__21492;
    wire N__21491;
    wire N__21490;
    wire N__21489;
    wire N__21472;
    wire N__21455;
    wire N__21452;
    wire N__21451;
    wire N__21448;
    wire N__21447;
    wire N__21442;
    wire N__21433;
    wire N__21428;
    wire N__21425;
    wire N__21422;
    wire N__21419;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21385;
    wire N__21380;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21323;
    wire N__21320;
    wire N__21317;
    wire N__21314;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21299;
    wire N__21296;
    wire N__21293;
    wire N__21292;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21278;
    wire N__21277;
    wire N__21274;
    wire N__21273;
    wire N__21272;
    wire N__21271;
    wire N__21270;
    wire N__21269;
    wire N__21266;
    wire N__21265;
    wire N__21264;
    wire N__21261;
    wire N__21254;
    wire N__21253;
    wire N__21248;
    wire N__21245;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21226;
    wire N__21223;
    wire N__21216;
    wire N__21213;
    wire N__21206;
    wire N__21203;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21191;
    wire N__21188;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21169;
    wire N__21166;
    wire N__21163;
    wire N__21158;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21143;
    wire N__21140;
    wire N__21139;
    wire N__21136;
    wire N__21133;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21071;
    wire N__21068;
    wire N__21065;
    wire N__21064;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21047;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21025;
    wire N__21022;
    wire N__21019;
    wire N__21014;
    wire N__21011;
    wire N__21010;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20998;
    wire N__20993;
    wire N__20990;
    wire N__20987;
    wire N__20986;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20974;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20962;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20938;
    wire N__20935;
    wire N__20932;
    wire N__20929;
    wire N__20924;
    wire N__20921;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20908;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20887;
    wire N__20884;
    wire N__20881;
    wire N__20878;
    wire N__20873;
    wire N__20870;
    wire N__20869;
    wire N__20864;
    wire N__20863;
    wire N__20860;
    wire N__20857;
    wire N__20852;
    wire N__20849;
    wire N__20848;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20835;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20823;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20803;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20779;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20752;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20735;
    wire N__20732;
    wire N__20731;
    wire N__20728;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20718;
    wire N__20715;
    wire N__20708;
    wire N__20705;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20697;
    wire N__20692;
    wire N__20689;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20668;
    wire N__20667;
    wire N__20666;
    wire N__20665;
    wire N__20664;
    wire N__20663;
    wire N__20662;
    wire N__20661;
    wire N__20658;
    wire N__20653;
    wire N__20646;
    wire N__20643;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20625;
    wire N__20622;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20543;
    wire N__20540;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20521;
    wire N__20520;
    wire N__20517;
    wire N__20516;
    wire N__20515;
    wire N__20512;
    wire N__20507;
    wire N__20506;
    wire N__20499;
    wire N__20496;
    wire N__20495;
    wire N__20492;
    wire N__20487;
    wire N__20484;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20452;
    wire N__20451;
    wire N__20448;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20432;
    wire N__20429;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20417;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20405;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20397;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20378;
    wire N__20375;
    wire N__20374;
    wire N__20373;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20354;
    wire N__20351;
    wire N__20350;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20330;
    wire N__20329;
    wire N__20328;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20296;
    wire N__20293;
    wire N__20290;
    wire N__20285;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20273;
    wire N__20272;
    wire N__20271;
    wire N__20270;
    wire N__20269;
    wire N__20268;
    wire N__20267;
    wire N__20266;
    wire N__20265;
    wire N__20264;
    wire N__20251;
    wire N__20242;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20206;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20196;
    wire N__20191;
    wire N__20188;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20125;
    wire N__20124;
    wire N__20123;
    wire N__20122;
    wire N__20121;
    wire N__20120;
    wire N__20119;
    wire N__20118;
    wire N__20117;
    wire N__20104;
    wire N__20095;
    wire N__20092;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20077;
    wire N__20076;
    wire N__20075;
    wire N__20074;
    wire N__20073;
    wire N__20070;
    wire N__20069;
    wire N__20068;
    wire N__20067;
    wire N__20066;
    wire N__20065;
    wire N__20064;
    wire N__20063;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20047;
    wire N__20046;
    wire N__20045;
    wire N__20042;
    wire N__20035;
    wire N__20022;
    wire N__20019;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20004;
    wire N__20003;
    wire N__20002;
    wire N__20001;
    wire N__20000;
    wire N__19999;
    wire N__19998;
    wire N__19997;
    wire N__19996;
    wire N__19995;
    wire N__19994;
    wire N__19993;
    wire N__19992;
    wire N__19991;
    wire N__19990;
    wire N__19989;
    wire N__19984;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19956;
    wire N__19941;
    wire N__19936;
    wire N__19925;
    wire N__19922;
    wire N__19921;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19909;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19895;
    wire N__19894;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19855;
    wire N__19854;
    wire N__19853;
    wire N__19850;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19840;
    wire N__19835;
    wire N__19828;
    wire N__19823;
    wire N__19822;
    wire N__19821;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19759;
    wire N__19758;
    wire N__19755;
    wire N__19754;
    wire N__19753;
    wire N__19750;
    wire N__19749;
    wire N__19748;
    wire N__19745;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19727;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19719;
    wire N__19718;
    wire N__19717;
    wire N__19714;
    wire N__19711;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19689;
    wire N__19680;
    wire N__19677;
    wire N__19672;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19447;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19423;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19345;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19270;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19253;
    wire N__19252;
    wire N__19249;
    wire N__19246;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19231;
    wire N__19228;
    wire N__19225;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19204;
    wire N__19203;
    wire N__19198;
    wire N__19195;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19183;
    wire N__19182;
    wire N__19179;
    wire N__19174;
    wire N__19169;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19138;
    wire N__19135;
    wire N__19132;
    wire N__19127;
    wire N__19126;
    wire N__19125;
    wire N__19124;
    wire N__19121;
    wire N__19120;
    wire N__19117;
    wire N__19116;
    wire N__19113;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19105;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19045;
    wire N__19044;
    wire N__19039;
    wire N__19036;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19013;
    wire N__19012;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18982;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18972;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_0 ;
    wire bfn_1_7_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_8 ;
    wire bfn_1_8_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15 ;
    wire bfn_1_9_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_15 ;
    wire bfn_1_10_0_;
    wire \pwm_generator_inst.un2_threshold_acc_2_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_18 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_20 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_21 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_22 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_23 ;
    wire bfn_1_11_0_;
    wire \pwm_generator_inst.un2_threshold_acc_2_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_24 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ;
    wire bfn_1_12_0_;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_25 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ;
    wire rgb_drv_RNOZ0;
    wire N_38_i_i;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_ ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_13_cascade_ ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17 ;
    wire \pwm_generator_inst.un3_threshold_acc ;
    wire bfn_2_10_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ;
    wire bfn_2_11_0_;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ;
    wire bfn_2_12_0_;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ;
    wire bfn_3_8_0_;
    wire \pwm_generator_inst.un19_threshold_acc_axb_1 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_2 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_3 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_5 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_6 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_7 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_7 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_8 ;
    wire bfn_3_9_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un1_duty_inputlt3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3_cascade_ ;
    wire pwm_duty_input_0;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire pwm_duty_input_2;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire pwm_duty_input_1;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.N_153 ;
    wire \current_shift_inst.PI_CTRL.N_154 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_2 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_3 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_7 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_8 ;
    wire \pwm_generator_inst.N_16 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ;
    wire N_19_1;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire pwm_duty_input_9;
    wire pwm_duty_input_7;
    wire pwm_duty_input_6;
    wire pwm_duty_input_8;
    wire pwm_duty_input_3;
    wire pwm_duty_input_4;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ;
    wire pwm_duty_input_5;
    wire \pwm_generator_inst.N_17 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.N_155 ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.N_149 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_53 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_1 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire bfn_5_10_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire bfn_5_11_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire bfn_5_12_0_;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire bfn_5_13_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire delay_hc_input_c_g;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire \pwm_generator_inst.threshold_ACCZ0Z_6 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_4 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_74_16_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_74_16 ;
    wire \current_shift_inst.PI_CTRL.N_74_21 ;
    wire \current_shift_inst.PI_CTRL.N_72 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_1_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_7_15_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire bfn_7_16_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.N_432_i ;
    wire il_max_comp1_c;
    wire il_max_comp2_c;
    wire il_min_comp2_c;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_75 ;
    wire \current_shift_inst.PI_CTRL.N_62 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ;
    wire bfn_8_15_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ;
    wire bfn_8_16_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ;
    wire bfn_8_17_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ;
    wire bfn_8_18_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_31 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_ ;
    wire elapsed_time_ns_1_RNI3VBED1_0_16_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2 ;
    wire elapsed_time_ns_1_RNI40CED1_0_17_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_cascade_ ;
    wire \pwm_generator_inst.thresholdZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_9_6_0_;
    wire \pwm_generator_inst.thresholdZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.thresholdZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.thresholdZ0Z_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.thresholdZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.thresholdZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.thresholdZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.thresholdZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.thresholdZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_9_7_0_;
    wire \pwm_generator_inst.thresholdZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire il_min_comp1_c;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_6 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.N_275_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_325_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1_cascade_ ;
    wire elapsed_time_ns_1_RNIB4DJ11_0_5_cascade_;
    wire elapsed_time_ns_1_RNIL13KD1_0_9;
    wire \phase_controller_inst1.stoper_hc.N_266_iZ0Z_1 ;
    wire elapsed_time_ns_1_RNI3VBED1_0_16;
    wire \phase_controller_inst1.stoper_hc.N_287 ;
    wire elapsed_time_ns_1_RNI1TBED1_0_14;
    wire elapsed_time_ns_1_RNI51CED1_0_18;
    wire elapsed_time_ns_1_RNI40CED1_0_17;
    wire elapsed_time_ns_1_RNI62CED1_0_19;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire s3_phy_c;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire il_max_comp2_D1;
    wire il_min_comp1_D1;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire bfn_10_13_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire bfn_10_14_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire bfn_10_15_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire bfn_10_16_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_29 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_30 ;
    wire bfn_10_17_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_23 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_ ;
    wire elapsed_time_ns_1_RNIP1MD11_0_12_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.N_337 ;
    wire elapsed_time_ns_1_RNINVLD11_0_10;
    wire elapsed_time_ns_1_RNIP2ND11_0_21;
    wire elapsed_time_ns_1_RNIP2ND11_0_21_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15_cascade_ ;
    wire elapsed_time_ns_1_RNIU7ND11_0_26;
    wire elapsed_time_ns_1_RNIR4ND11_0_23;
    wire elapsed_time_ns_1_RNIR4ND11_0_23_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15 ;
    wire elapsed_time_ns_1_RNI0AND11_0_28;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15 ;
    wire elapsed_time_ns_1_RNI1BND11_0_29;
    wire elapsed_time_ns_1_RNIO1ND11_0_20;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15_cascade_ ;
    wire elapsed_time_ns_1_RNIV8ND11_0_27;
    wire \phase_controller_inst2.stoper_hc.un6_running_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_10_21_0_;
    wire \phase_controller_inst2.stoper_hc.un6_running_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_10_22_0_;
    wire \phase_controller_inst2.stoper_hc.un6_running_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_16 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_17 ;
    wire bfn_10_23_0_;
    wire \phase_controller_inst2.stoper_hc.un6_running_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ;
    wire bfn_10_24_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJBZ0Z21 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_10_25_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire bfn_10_26_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire bfn_11_6_0_;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire bfn_11_7_0_;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_21 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_20 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.N_103 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire elapsed_time_ns_1_RNIO0MD11_0_11;
    wire elapsed_time_ns_1_RNIP1MD11_0_12;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2Z0Z_10 ;
    wire elapsed_time_ns_1_RNIQ2MD11_0_13;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ;
    wire elapsed_time_ns_1_RNID6DJ11_0_7;
    wire elapsed_time_ns_1_RNIE7DJ11_0_8;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ;
    wire elapsed_time_ns_1_RNIDP2KD1_0_1;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ;
    wire elapsed_time_ns_1_RNIDP2KD1_0_1_cascade_;
    wire \phase_controller_inst1.stoper_hc.N_307 ;
    wire elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ;
    wire elapsed_time_ns_1_RNIA3DJ11_0_4;
    wire \phase_controller_inst1.stoper_hc.N_325 ;
    wire elapsed_time_ns_1_RNIQ4OD11_0_31;
    wire elapsed_time_ns_1_RNIB4DJ11_0_5;
    wire \phase_controller_inst1.stoper_hc.N_327 ;
    wire elapsed_time_ns_1_RNIP3OD11_0_30;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.N_382_i_cascade_ ;
    wire elapsed_time_ns_1_RNIS5ND11_0_24;
    wire elapsed_time_ns_1_RNIT6ND11_0_25;
    wire elapsed_time_ns_1_RNIS4MD11_0_15;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16 ;
    wire elapsed_time_ns_1_RNIQ3ND11_0_22;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_ ;
    wire elapsed_time_ns_1_RNIQURR91_0_3;
    wire elapsed_time_ns_1_RNIQURR91_0_3_cascade_;
    wire \phase_controller_inst1.stoper_hc.N_283 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire s4_phy_c;
    wire il_max_comp1_D1;
    wire il_min_comp2_D1;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst1.N_55 ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst1.start_timer_tr_0_sqmuxa ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire il_max_comp1_D2;
    wire \phase_controller_inst1.N_56 ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ;
    wire bfn_12_13_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNII3DZ0Z41 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire bfn_12_14_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_12_15_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_12_16_0_;
    wire \phase_controller_inst1.stoper_hc.un6_running_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_12_17_0_;
    wire \phase_controller_inst1.stoper_hc.un6_running_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_17 ;
    wire bfn_12_18_0_;
    wire \phase_controller_inst1.stoper_hc.un6_running_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ;
    wire elapsed_time_ns_1_RNIIU2KD1_0_6;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5 ;
    wire elapsed_time_ns_1_RNIIU2KD1_0_6_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire bfn_12_20_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lto6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire bfn_12_21_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lto14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc5lto15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire bfn_12_22_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire bfn_12_23_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire \pll_inst.red_c_i ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6_cascade_ ;
    wire elapsed_time_ns_1_RNIUKL2M1_0_6_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19_cascade_ ;
    wire elapsed_time_ns_1_RNIIJ4DM1_0_19_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ;
    wire bfn_13_11_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire bfn_13_12_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_13_13_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.time_passed_RNI9M3O_cascade_ ;
    wire state_3;
    wire s1_phy_c;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_28 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire bfn_13_21_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_13_22_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_13_23_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_13_24_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.N_433_i ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.N_166_i ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_ ;
    wire elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_;
    wire elapsed_time_ns_1_RNIUKL2M1_0_6;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ;
    wire elapsed_time_ns_1_RNIUCHF91_0_15_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9 ;
    wire elapsed_time_ns_1_RNI1OL2M1_0_9_cascade_;
    wire \phase_controller_inst1.stoper_tr.N_211_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1 ;
    wire elapsed_time_ns_1_RNIPFL2M1_0_1;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2 ;
    wire elapsed_time_ns_1_RNICG2591_0_4;
    wire elapsed_time_ns_1_RNICG2591_0_4_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16_cascade_ ;
    wire elapsed_time_ns_1_RNIFG4DM1_0_16;
    wire elapsed_time_ns_1_RNIGH4DM1_0_17_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18_cascade_ ;
    wire elapsed_time_ns_1_RNIHI4DM1_0_18_cascade_;
    wire elapsed_time_ns_1_RNIGH4DM1_0_17;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.N_251 ;
    wire elapsed_time_ns_1_RNISCJF91_0_31_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9 ;
    wire elapsed_time_ns_1_RNI1OL2M1_0_9;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_ ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIP6NZ0Z32 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_0_12 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire bfn_14_17_0_;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire bfn_14_18_0_;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire bfn_14_19_0_;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire bfn_14_20_0_;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.N_432_i_g ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire il_max_comp2_D2;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa ;
    wire \delay_measurement_inst.delay_tr_timer.N_434_i ;
    wire bfn_15_5_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_15_6_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_15_7_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_15_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire elapsed_time_ns_1_RNIGK2591_0_8;
    wire elapsed_time_ns_1_RNIHI4DM1_0_18;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.N_214 ;
    wire elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_;
    wire elapsed_time_ns_1_RNIUCHF91_0_15;
    wire \phase_controller_inst1.stoper_tr.N_241_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un6_running_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_15_11_0_;
    wire \phase_controller_inst1.stoper_tr.un6_running_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_15_12_0_;
    wire \phase_controller_inst1.stoper_tr.un6_running_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_17 ;
    wire bfn_15_13_0_;
    wire \phase_controller_inst1.stoper_tr.un6_running_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire bfn_15_14_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ;
    wire bfn_15_15_0_;
    wire \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ;
    wire bfn_15_16_0_;
    wire \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire bfn_15_17_0_;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire bfn_15_20_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire bfn_15_21_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire bfn_15_22_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire bfn_15_23_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \phase_controller_inst2.start_timer_hc_RNOZ0Z_0 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_435_i ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ;
    wire elapsed_time_ns_1_RNIAE2591_0_2;
    wire bfn_16_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_16_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire bfn_16_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_16_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire T45_c;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.control_input_1_axb_0 ;
    wire \current_shift_inst.N_1572_i ;
    wire \current_shift_inst.control_inputZ0Z_0 ;
    wire bfn_16_15_0_;
    wire \current_shift_inst.control_inputZ0Z_1 ;
    wire \current_shift_inst.control_input_1_cry_0 ;
    wire \current_shift_inst.control_inputZ0Z_2 ;
    wire \current_shift_inst.control_input_1_cry_1 ;
    wire \current_shift_inst.control_input_1_axb_3 ;
    wire \current_shift_inst.control_inputZ0Z_3 ;
    wire \current_shift_inst.control_input_1_cry_2 ;
    wire \current_shift_inst.control_input_1_axb_4 ;
    wire \current_shift_inst.control_inputZ0Z_4 ;
    wire \current_shift_inst.control_input_1_cry_3 ;
    wire \current_shift_inst.control_input_1_axb_5 ;
    wire \current_shift_inst.control_inputZ0Z_5 ;
    wire \current_shift_inst.control_input_1_cry_4 ;
    wire \current_shift_inst.control_inputZ0Z_6 ;
    wire \current_shift_inst.control_input_1_cry_5 ;
    wire \current_shift_inst.control_inputZ0Z_7 ;
    wire \current_shift_inst.control_input_1_cry_6 ;
    wire \current_shift_inst.control_input_1_cry_7 ;
    wire \current_shift_inst.control_inputZ0Z_8 ;
    wire bfn_16_16_0_;
    wire \current_shift_inst.control_input_1_cry_8 ;
    wire \current_shift_inst.control_inputZ0Z_10 ;
    wire \current_shift_inst.control_input_1_cry_9 ;
    wire \current_shift_inst.control_input_1_axb_11 ;
    wire \current_shift_inst.control_input_1_cry_10 ;
    wire \current_shift_inst.control_inputZ0Z_11 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.control_input_1_axb_1 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.control_input_1_axb_7 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.control_input_1_axb_10 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.control_input_1_axb_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire bfn_16_17_0_;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire bfn_16_18_0_;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire bfn_16_19_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_16_20_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_16_22_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_16_23_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_16_24_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_16_25_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_167_i ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_434_i_g ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.delay_tr_timer.N_341 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ;
    wire elapsed_time_ns_1_RNIRHL2M1_0_3;
    wire \delay_measurement_inst.delay_tr_timer.N_381_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_358_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_381 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.N_348_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire elapsed_time_ns_1_RNIFJ2591_0_7;
    wire elapsed_time_ns_1_RNITCIF91_0_23;
    wire elapsed_time_ns_1_RNITCIF91_0_23_cascade_;
    wire elapsed_time_ns_1_RNIRAIF91_0_21;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire elapsed_time_ns_1_RNIDH2591_0_5;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.N_347 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire elapsed_time_ns_1_RNIQ8HF91_0_11;
    wire elapsed_time_ns_1_RNIQ8HF91_0_11_cascade_;
    wire elapsed_time_ns_1_RNIR9HF91_0_12;
    wire \phase_controller_inst1.stoper_tr.N_244 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire elapsed_time_ns_1_RNI3JIF91_0_29;
    wire elapsed_time_ns_1_RNI3JIF91_0_29_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15 ;
    wire elapsed_time_ns_1_RNIDE4DM1_0_14;
    wire \phase_controller_inst1.stoper_tr.un6_running_14 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire elapsed_time_ns_1_RNISAHF91_0_13;
    wire \phase_controller_inst1.stoper_tr.N_241 ;
    wire elapsed_time_ns_1_RNISAHF91_0_13_cascade_;
    wire \phase_controller_inst1.stoper_tr.un6_running_13 ;
    wire elapsed_time_ns_1_RNIIJ4DM1_0_19;
    wire elapsed_time_ns_1_RNISCJF91_0_31;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_19 ;
    wire \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_17_11_0_;
    wire \phase_controller_inst2.stoper_tr.un6_running_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_17_12_0_;
    wire \phase_controller_inst2.stoper_tr.un6_running_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_17 ;
    wire bfn_17_13_0_;
    wire \phase_controller_inst2.stoper_tr.un6_running_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_19 ;
    wire start_stop_c;
    wire state_ns_i_a3_1;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ;
    wire bfn_17_14_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_17_15_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire bfn_17_16_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.timer_s1.N_166_i_g ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.control_input_1_axb_6 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.control_input_1_axb_8 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.control_input_1_axb_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.N_382_i ;
    wire elapsed_time_ns_1_RNI81DJ11_0_2;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire T01_c;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire T12_c;
    wire \delay_measurement_inst.delay_tr_timer.N_367 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ;
    wire \delay_measurement_inst.delay_tr_timer.N_349 ;
    wire \delay_measurement_inst.delay_tr_timer.N_363_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9 ;
    wire \delay_measurement_inst.delay_tr_timer.N_380 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7 ;
    wire \delay_measurement_inst.delay_tr_timer.N_365 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_345 ;
    wire \delay_measurement_inst.delay_tr_timer.N_359_1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire elapsed_time_ns_1_RNIUDIF91_0_24;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire elapsed_time_ns_1_RNIVEIF91_0_25;
    wire elapsed_time_ns_1_RNIVEIF91_0_25_cascade_;
    wire elapsed_time_ns_1_RNI0GIF91_0_26;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire elapsed_time_ns_1_RNI2IIF91_0_28;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.delay_tr_timer.N_378 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_ ;
    wire elapsed_time_ns_1_RNIP7HF91_0_10;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire elapsed_time_ns_1_RNI1HIF91_0_27;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire elapsed_time_ns_1_RNISBIF91_0_22;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire elapsed_time_ns_1_RNIQ9IF91_0_20;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ;
    wire elapsed_time_ns_1_RNIRBJF91_0_30;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire il_min_comp2_D2;
    wire \phase_controller_inst2.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_inst2.time_passed_RNI9M3O ;
    wire phase_controller_inst1_state_4;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIUMLHZ0Z1 ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire bfn_18_14_0_;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ;
    wire bfn_18_15_0_;
    wire \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire bfn_18_16_0_;
    wire \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire bfn_18_17_0_;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un4_control_input_0_31 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ;
    wire \current_shift_inst.control_inputZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire delay_tr_input_c_g;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire T23_c;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__21362),
            .RESETB(N__31034),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__37810),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__37803),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({dangling_wire_16,N__20002,N__19995,N__20000,N__19994,N__20001,N__19993,N__20003,N__19990,N__19996,N__19989,N__19997,N__19991,N__19998,N__19992,N__19999}),
            .C({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32}),
            .B({dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__37809,N__37806,dangling_wire_40,dangling_wire_41,dangling_wire_42,N__37804,N__37808,N__37805,N__37807}),
            .OHOLDTOP(),
            .O({dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,\pwm_generator_inst.un2_threshold_acc_2_1_16 ,\pwm_generator_inst.un2_threshold_acc_2_1_15 ,\pwm_generator_inst.un2_threshold_acc_2_14 ,\pwm_generator_inst.un2_threshold_acc_2_13 ,\pwm_generator_inst.un2_threshold_acc_2_12 ,\pwm_generator_inst.un2_threshold_acc_2_11 ,\pwm_generator_inst.un2_threshold_acc_2_10 ,\pwm_generator_inst.un2_threshold_acc_2_9 ,\pwm_generator_inst.un2_threshold_acc_2_8 ,\pwm_generator_inst.un2_threshold_acc_2_7 ,\pwm_generator_inst.un2_threshold_acc_2_6 ,\pwm_generator_inst.un2_threshold_acc_2_5 ,\pwm_generator_inst.un2_threshold_acc_2_4 ,\pwm_generator_inst.un2_threshold_acc_2_3 ,\pwm_generator_inst.un2_threshold_acc_2_2 ,\pwm_generator_inst.un2_threshold_acc_2_1 ,\pwm_generator_inst.un2_threshold_acc_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__37730),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__37723),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .ADDSUBBOT(),
            .A({dangling_wire_74,N__20066,N__20045,N__20067,N__20046,N__20068,N__20456,N__20378,N__20416,N__20405,N__20284,N__20328,N__20354,N__19913,N__19886,N__19658}),
            .C({dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90}),
            .B({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,N__37729,N__37726,dangling_wire_98,dangling_wire_99,dangling_wire_100,N__37724,N__37728,N__37725,N__37727}),
            .OHOLDTOP(),
            .O({dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\pwm_generator_inst.un2_threshold_acc_1_25 ,\pwm_generator_inst.un2_threshold_acc_1_24 ,\pwm_generator_inst.un2_threshold_acc_1_23 ,\pwm_generator_inst.un2_threshold_acc_1_22 ,\pwm_generator_inst.un2_threshold_acc_1_21 ,\pwm_generator_inst.un2_threshold_acc_1_20 ,\pwm_generator_inst.un2_threshold_acc_1_19 ,\pwm_generator_inst.un2_threshold_acc_1_18 ,\pwm_generator_inst.un2_threshold_acc_1_17 ,\pwm_generator_inst.un2_threshold_acc_1_16 ,\pwm_generator_inst.un2_threshold_acc_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold_acc ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__47637),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__47639),
            .DIN(N__47638),
            .DOUT(N__47637),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__47639),
            .PADOUT(N__47638),
            .PADIN(N__47637),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T01_obuf_iopad (
            .OE(N__47628),
            .DIN(N__47627),
            .DOUT(N__47626),
            .PACKAGEPIN(T01));
    defparam T01_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T01_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T01_obuf_preio (
            .PADOEN(N__47628),
            .PADOUT(N__47627),
            .PADIN(N__47626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__41909),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__47619),
            .DIN(N__47618),
            .DOUT(N__47617),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__47619),
            .PADOUT(N__47618),
            .PADIN(N__47617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__47610),
            .DIN(N__47609),
            .DOUT(N__47608),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__47610),
            .PADOUT(N__47609),
            .PADIN(N__47608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T23_obuf_iopad (
            .OE(N__47601),
            .DIN(N__47600),
            .DOUT(N__47599),
            .PACKAGEPIN(T23));
    defparam T23_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T23_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T23_obuf_preio (
            .PADOEN(N__47601),
            .PADOUT(N__47600),
            .PADIN(N__47599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__46133),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__47592),
            .DIN(N__47591),
            .DOUT(N__47590),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__47592),
            .PADOUT(N__47591),
            .PADIN(N__47590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22349),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__47583),
            .DIN(N__47582),
            .DOUT(N__47581),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__47583),
            .PADOUT(N__47582),
            .PADIN(N__47581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__47574),
            .DIN(N__47573),
            .DOUT(N__47572),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__47574),
            .PADOUT(N__47573),
            .PADIN(N__47572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31046),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T12_obuf_iopad (
            .OE(N__47565),
            .DIN(N__47564),
            .DOUT(N__47563),
            .PACKAGEPIN(T12));
    defparam T12_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T12_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T12_obuf_preio (
            .PADOEN(N__47565),
            .PADOUT(N__47564),
            .PADIN(N__47563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__41804),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__47556),
            .DIN(N__47555),
            .DOUT(N__47554),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__47556),
            .PADOUT(N__47555),
            .PADIN(N__47554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__47547),
            .DIN(N__47546),
            .DOUT(N__47545),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__47547),
            .PADOUT(N__47546),
            .PADIN(N__47545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31211),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__47538),
            .DIN(N__47537),
            .DOUT(N__47536),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__47538),
            .PADOUT(N__47537),
            .PADIN(N__47536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28664),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__47529),
            .DIN(N__47528),
            .DOUT(N__47527),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__47529),
            .PADOUT(N__47528),
            .PADIN(N__47527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__47520),
            .DIN(N__47519),
            .DOUT(N__47518),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__47520),
            .PADOUT(N__47519),
            .PADIN(N__47518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23615),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T45_obuf_iopad (
            .OE(N__47511),
            .DIN(N__47510),
            .DOUT(N__47509),
            .PACKAGEPIN(T45));
    defparam T45_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T45_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T45_obuf_preio (
            .PADOEN(N__47511),
            .PADOUT(N__47510),
            .PADIN(N__47509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36809),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__47502),
            .DIN(N__47501),
            .DOUT(N__47500),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__47502),
            .PADOUT(N__47501),
            .PADIN(N__47500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__47493),
            .DIN(N__47492),
            .DOUT(N__47491),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__47493),
            .PADOUT(N__47492),
            .PADIN(N__47491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__11239 (
            .O(N__47474),
            .I(N__47471));
    InMux I__11238 (
            .O(N__47471),
            .I(N__47467));
    InMux I__11237 (
            .O(N__47470),
            .I(N__47463));
    LocalMux I__11236 (
            .O(N__47467),
            .I(N__47460));
    InMux I__11235 (
            .O(N__47466),
            .I(N__47457));
    LocalMux I__11234 (
            .O(N__47463),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv12 I__11233 (
            .O(N__47460),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__11232 (
            .O(N__47457),
            .I(\current_shift_inst.un4_control_input1_20 ));
    CascadeMux I__11231 (
            .O(N__47450),
            .I(N__47446));
    InMux I__11230 (
            .O(N__47449),
            .I(N__47443));
    InMux I__11229 (
            .O(N__47446),
            .I(N__47440));
    LocalMux I__11228 (
            .O(N__47443),
            .I(N__47436));
    LocalMux I__11227 (
            .O(N__47440),
            .I(N__47433));
    InMux I__11226 (
            .O(N__47439),
            .I(N__47430));
    Span4Mux_h I__11225 (
            .O(N__47436),
            .I(N__47424));
    Span4Mux_h I__11224 (
            .O(N__47433),
            .I(N__47424));
    LocalMux I__11223 (
            .O(N__47430),
            .I(N__47421));
    InMux I__11222 (
            .O(N__47429),
            .I(N__47418));
    Odrv4 I__11221 (
            .O(N__47424),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__11220 (
            .O(N__47421),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    LocalMux I__11219 (
            .O(N__47418),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__11218 (
            .O(N__47411),
            .I(N__47408));
    LocalMux I__11217 (
            .O(N__47408),
            .I(N__47405));
    Span4Mux_h I__11216 (
            .O(N__47405),
            .I(N__47402));
    Odrv4 I__11215 (
            .O(N__47402),
            .I(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ));
    InMux I__11214 (
            .O(N__47399),
            .I(N__47396));
    LocalMux I__11213 (
            .O(N__47396),
            .I(N__47393));
    Span4Mux_v I__11212 (
            .O(N__47393),
            .I(N__47390));
    Odrv4 I__11211 (
            .O(N__47390),
            .I(\current_shift_inst.control_inputZ0Z_9 ));
    InMux I__11210 (
            .O(N__47387),
            .I(N__47384));
    LocalMux I__11209 (
            .O(N__47384),
            .I(N__47381));
    Span4Mux_h I__11208 (
            .O(N__47381),
            .I(N__47378));
    Span4Mux_h I__11207 (
            .O(N__47378),
            .I(N__47375));
    Span4Mux_h I__11206 (
            .O(N__47375),
            .I(N__47372));
    Odrv4 I__11205 (
            .O(N__47372),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__11204 (
            .O(N__47369),
            .I(N__47347));
    InMux I__11203 (
            .O(N__47368),
            .I(N__47329));
    InMux I__11202 (
            .O(N__47367),
            .I(N__47322));
    InMux I__11201 (
            .O(N__47366),
            .I(N__47311));
    InMux I__11200 (
            .O(N__47365),
            .I(N__47311));
    InMux I__11199 (
            .O(N__47364),
            .I(N__47311));
    InMux I__11198 (
            .O(N__47363),
            .I(N__47311));
    InMux I__11197 (
            .O(N__47362),
            .I(N__47311));
    InMux I__11196 (
            .O(N__47361),
            .I(N__47308));
    InMux I__11195 (
            .O(N__47360),
            .I(N__47299));
    InMux I__11194 (
            .O(N__47359),
            .I(N__47299));
    InMux I__11193 (
            .O(N__47358),
            .I(N__47299));
    InMux I__11192 (
            .O(N__47357),
            .I(N__47299));
    InMux I__11191 (
            .O(N__47356),
            .I(N__47292));
    InMux I__11190 (
            .O(N__47355),
            .I(N__47292));
    InMux I__11189 (
            .O(N__47354),
            .I(N__47292));
    InMux I__11188 (
            .O(N__47353),
            .I(N__47289));
    InMux I__11187 (
            .O(N__47352),
            .I(N__47286));
    InMux I__11186 (
            .O(N__47351),
            .I(N__47281));
    InMux I__11185 (
            .O(N__47350),
            .I(N__47281));
    LocalMux I__11184 (
            .O(N__47347),
            .I(N__47278));
    InMux I__11183 (
            .O(N__47346),
            .I(N__47265));
    InMux I__11182 (
            .O(N__47345),
            .I(N__47265));
    InMux I__11181 (
            .O(N__47344),
            .I(N__47265));
    InMux I__11180 (
            .O(N__47343),
            .I(N__47265));
    InMux I__11179 (
            .O(N__47342),
            .I(N__47265));
    InMux I__11178 (
            .O(N__47341),
            .I(N__47265));
    InMux I__11177 (
            .O(N__47340),
            .I(N__47258));
    InMux I__11176 (
            .O(N__47339),
            .I(N__47258));
    InMux I__11175 (
            .O(N__47338),
            .I(N__47258));
    InMux I__11174 (
            .O(N__47337),
            .I(N__47253));
    InMux I__11173 (
            .O(N__47336),
            .I(N__47250));
    InMux I__11172 (
            .O(N__47335),
            .I(N__47241));
    InMux I__11171 (
            .O(N__47334),
            .I(N__47241));
    InMux I__11170 (
            .O(N__47333),
            .I(N__47241));
    InMux I__11169 (
            .O(N__47332),
            .I(N__47241));
    LocalMux I__11168 (
            .O(N__47329),
            .I(N__47238));
    InMux I__11167 (
            .O(N__47328),
            .I(N__47229));
    InMux I__11166 (
            .O(N__47327),
            .I(N__47229));
    InMux I__11165 (
            .O(N__47326),
            .I(N__47229));
    InMux I__11164 (
            .O(N__47325),
            .I(N__47229));
    LocalMux I__11163 (
            .O(N__47322),
            .I(N__47218));
    LocalMux I__11162 (
            .O(N__47311),
            .I(N__47215));
    LocalMux I__11161 (
            .O(N__47308),
            .I(N__47206));
    LocalMux I__11160 (
            .O(N__47299),
            .I(N__47206));
    LocalMux I__11159 (
            .O(N__47292),
            .I(N__47206));
    LocalMux I__11158 (
            .O(N__47289),
            .I(N__47206));
    LocalMux I__11157 (
            .O(N__47286),
            .I(N__47188));
    LocalMux I__11156 (
            .O(N__47281),
            .I(N__47188));
    Span4Mux_v I__11155 (
            .O(N__47278),
            .I(N__47181));
    LocalMux I__11154 (
            .O(N__47265),
            .I(N__47181));
    LocalMux I__11153 (
            .O(N__47258),
            .I(N__47181));
    InMux I__11152 (
            .O(N__47257),
            .I(N__47172));
    InMux I__11151 (
            .O(N__47256),
            .I(N__47172));
    LocalMux I__11150 (
            .O(N__47253),
            .I(N__47169));
    LocalMux I__11149 (
            .O(N__47250),
            .I(N__47160));
    LocalMux I__11148 (
            .O(N__47241),
            .I(N__47160));
    Span4Mux_h I__11147 (
            .O(N__47238),
            .I(N__47160));
    LocalMux I__11146 (
            .O(N__47229),
            .I(N__47160));
    InMux I__11145 (
            .O(N__47228),
            .I(N__47143));
    InMux I__11144 (
            .O(N__47227),
            .I(N__47143));
    InMux I__11143 (
            .O(N__47226),
            .I(N__47143));
    InMux I__11142 (
            .O(N__47225),
            .I(N__47143));
    InMux I__11141 (
            .O(N__47224),
            .I(N__47143));
    InMux I__11140 (
            .O(N__47223),
            .I(N__47143));
    InMux I__11139 (
            .O(N__47222),
            .I(N__47143));
    InMux I__11138 (
            .O(N__47221),
            .I(N__47143));
    Span4Mux_h I__11137 (
            .O(N__47218),
            .I(N__47136));
    Span4Mux_v I__11136 (
            .O(N__47215),
            .I(N__47136));
    Span4Mux_v I__11135 (
            .O(N__47206),
            .I(N__47136));
    InMux I__11134 (
            .O(N__47205),
            .I(N__47119));
    InMux I__11133 (
            .O(N__47204),
            .I(N__47119));
    InMux I__11132 (
            .O(N__47203),
            .I(N__47119));
    InMux I__11131 (
            .O(N__47202),
            .I(N__47119));
    InMux I__11130 (
            .O(N__47201),
            .I(N__47119));
    InMux I__11129 (
            .O(N__47200),
            .I(N__47119));
    InMux I__11128 (
            .O(N__47199),
            .I(N__47119));
    InMux I__11127 (
            .O(N__47198),
            .I(N__47119));
    InMux I__11126 (
            .O(N__47197),
            .I(N__47110));
    InMux I__11125 (
            .O(N__47196),
            .I(N__47110));
    InMux I__11124 (
            .O(N__47195),
            .I(N__47110));
    InMux I__11123 (
            .O(N__47194),
            .I(N__47110));
    CascadeMux I__11122 (
            .O(N__47193),
            .I(N__47106));
    Span4Mux_v I__11121 (
            .O(N__47188),
            .I(N__47100));
    Span4Mux_v I__11120 (
            .O(N__47181),
            .I(N__47097));
    InMux I__11119 (
            .O(N__47180),
            .I(N__47088));
    InMux I__11118 (
            .O(N__47179),
            .I(N__47088));
    InMux I__11117 (
            .O(N__47178),
            .I(N__47088));
    InMux I__11116 (
            .O(N__47177),
            .I(N__47088));
    LocalMux I__11115 (
            .O(N__47172),
            .I(N__47085));
    Span4Mux_h I__11114 (
            .O(N__47169),
            .I(N__47072));
    Span4Mux_v I__11113 (
            .O(N__47160),
            .I(N__47072));
    LocalMux I__11112 (
            .O(N__47143),
            .I(N__47072));
    Span4Mux_h I__11111 (
            .O(N__47136),
            .I(N__47072));
    LocalMux I__11110 (
            .O(N__47119),
            .I(N__47072));
    LocalMux I__11109 (
            .O(N__47110),
            .I(N__47072));
    InMux I__11108 (
            .O(N__47109),
            .I(N__47061));
    InMux I__11107 (
            .O(N__47106),
            .I(N__47061));
    InMux I__11106 (
            .O(N__47105),
            .I(N__47061));
    InMux I__11105 (
            .O(N__47104),
            .I(N__47061));
    InMux I__11104 (
            .O(N__47103),
            .I(N__47061));
    Odrv4 I__11103 (
            .O(N__47100),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__11102 (
            .O(N__47097),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11101 (
            .O(N__47088),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv12 I__11100 (
            .O(N__47085),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__11099 (
            .O(N__47072),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__11098 (
            .O(N__47061),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    InMux I__11097 (
            .O(N__47048),
            .I(N__47043));
    InMux I__11096 (
            .O(N__47047),
            .I(N__47040));
    InMux I__11095 (
            .O(N__47046),
            .I(N__47037));
    LocalMux I__11094 (
            .O(N__47043),
            .I(N__47034));
    LocalMux I__11093 (
            .O(N__47040),
            .I(N__47031));
    LocalMux I__11092 (
            .O(N__47037),
            .I(N__47028));
    Span12Mux_v I__11091 (
            .O(N__47034),
            .I(N__47024));
    Span4Mux_h I__11090 (
            .O(N__47031),
            .I(N__47021));
    Sp12to4 I__11089 (
            .O(N__47028),
            .I(N__47018));
    InMux I__11088 (
            .O(N__47027),
            .I(N__47015));
    Odrv12 I__11087 (
            .O(N__47024),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv4 I__11086 (
            .O(N__47021),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv12 I__11085 (
            .O(N__47018),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__11084 (
            .O(N__47015),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    CascadeMux I__11083 (
            .O(N__47006),
            .I(N__46999));
    CascadeMux I__11082 (
            .O(N__47005),
            .I(N__46996));
    CascadeMux I__11081 (
            .O(N__47004),
            .I(N__46993));
    CascadeMux I__11080 (
            .O(N__47003),
            .I(N__46989));
    InMux I__11079 (
            .O(N__47002),
            .I(N__46977));
    InMux I__11078 (
            .O(N__46999),
            .I(N__46954));
    InMux I__11077 (
            .O(N__46996),
            .I(N__46951));
    InMux I__11076 (
            .O(N__46993),
            .I(N__46948));
    InMux I__11075 (
            .O(N__46992),
            .I(N__46943));
    InMux I__11074 (
            .O(N__46989),
            .I(N__46943));
    InMux I__11073 (
            .O(N__46988),
            .I(N__46934));
    InMux I__11072 (
            .O(N__46987),
            .I(N__46934));
    InMux I__11071 (
            .O(N__46986),
            .I(N__46934));
    InMux I__11070 (
            .O(N__46985),
            .I(N__46934));
    InMux I__11069 (
            .O(N__46984),
            .I(N__46927));
    InMux I__11068 (
            .O(N__46983),
            .I(N__46927));
    InMux I__11067 (
            .O(N__46982),
            .I(N__46927));
    CascadeMux I__11066 (
            .O(N__46981),
            .I(N__46923));
    CascadeMux I__11065 (
            .O(N__46980),
            .I(N__46919));
    LocalMux I__11064 (
            .O(N__46977),
            .I(N__46908));
    InMux I__11063 (
            .O(N__46976),
            .I(N__46899));
    InMux I__11062 (
            .O(N__46975),
            .I(N__46899));
    InMux I__11061 (
            .O(N__46974),
            .I(N__46899));
    InMux I__11060 (
            .O(N__46973),
            .I(N__46899));
    InMux I__11059 (
            .O(N__46972),
            .I(N__46892));
    InMux I__11058 (
            .O(N__46971),
            .I(N__46892));
    InMux I__11057 (
            .O(N__46970),
            .I(N__46892));
    InMux I__11056 (
            .O(N__46969),
            .I(N__46887));
    InMux I__11055 (
            .O(N__46968),
            .I(N__46887));
    CascadeMux I__11054 (
            .O(N__46967),
            .I(N__46868));
    CascadeMux I__11053 (
            .O(N__46966),
            .I(N__46864));
    CascadeMux I__11052 (
            .O(N__46965),
            .I(N__46860));
    CascadeMux I__11051 (
            .O(N__46964),
            .I(N__46856));
    CascadeMux I__11050 (
            .O(N__46963),
            .I(N__46852));
    CascadeMux I__11049 (
            .O(N__46962),
            .I(N__46848));
    CascadeMux I__11048 (
            .O(N__46961),
            .I(N__46844));
    CascadeMux I__11047 (
            .O(N__46960),
            .I(N__46840));
    CascadeMux I__11046 (
            .O(N__46959),
            .I(N__46836));
    CascadeMux I__11045 (
            .O(N__46958),
            .I(N__46832));
    CascadeMux I__11044 (
            .O(N__46957),
            .I(N__46828));
    LocalMux I__11043 (
            .O(N__46954),
            .I(N__46819));
    LocalMux I__11042 (
            .O(N__46951),
            .I(N__46819));
    LocalMux I__11041 (
            .O(N__46948),
            .I(N__46816));
    LocalMux I__11040 (
            .O(N__46943),
            .I(N__46813));
    LocalMux I__11039 (
            .O(N__46934),
            .I(N__46808));
    LocalMux I__11038 (
            .O(N__46927),
            .I(N__46808));
    InMux I__11037 (
            .O(N__46926),
            .I(N__46789));
    InMux I__11036 (
            .O(N__46923),
            .I(N__46789));
    InMux I__11035 (
            .O(N__46922),
            .I(N__46789));
    InMux I__11034 (
            .O(N__46919),
            .I(N__46789));
    InMux I__11033 (
            .O(N__46918),
            .I(N__46789));
    CascadeMux I__11032 (
            .O(N__46917),
            .I(N__46785));
    CascadeMux I__11031 (
            .O(N__46916),
            .I(N__46781));
    CascadeMux I__11030 (
            .O(N__46915),
            .I(N__46777));
    CascadeMux I__11029 (
            .O(N__46914),
            .I(N__46773));
    CascadeMux I__11028 (
            .O(N__46913),
            .I(N__46769));
    CascadeMux I__11027 (
            .O(N__46912),
            .I(N__46765));
    CascadeMux I__11026 (
            .O(N__46911),
            .I(N__46761));
    Span4Mux_v I__11025 (
            .O(N__46908),
            .I(N__46751));
    LocalMux I__11024 (
            .O(N__46899),
            .I(N__46751));
    LocalMux I__11023 (
            .O(N__46892),
            .I(N__46748));
    LocalMux I__11022 (
            .O(N__46887),
            .I(N__46745));
    InMux I__11021 (
            .O(N__46886),
            .I(N__46742));
    InMux I__11020 (
            .O(N__46885),
            .I(N__46725));
    InMux I__11019 (
            .O(N__46884),
            .I(N__46725));
    InMux I__11018 (
            .O(N__46883),
            .I(N__46725));
    InMux I__11017 (
            .O(N__46882),
            .I(N__46725));
    InMux I__11016 (
            .O(N__46881),
            .I(N__46725));
    InMux I__11015 (
            .O(N__46880),
            .I(N__46725));
    InMux I__11014 (
            .O(N__46879),
            .I(N__46725));
    InMux I__11013 (
            .O(N__46878),
            .I(N__46725));
    InMux I__11012 (
            .O(N__46877),
            .I(N__46714));
    InMux I__11011 (
            .O(N__46876),
            .I(N__46714));
    InMux I__11010 (
            .O(N__46875),
            .I(N__46714));
    InMux I__11009 (
            .O(N__46874),
            .I(N__46714));
    InMux I__11008 (
            .O(N__46873),
            .I(N__46714));
    InMux I__11007 (
            .O(N__46872),
            .I(N__46697));
    InMux I__11006 (
            .O(N__46871),
            .I(N__46697));
    InMux I__11005 (
            .O(N__46868),
            .I(N__46697));
    InMux I__11004 (
            .O(N__46867),
            .I(N__46697));
    InMux I__11003 (
            .O(N__46864),
            .I(N__46697));
    InMux I__11002 (
            .O(N__46863),
            .I(N__46697));
    InMux I__11001 (
            .O(N__46860),
            .I(N__46697));
    InMux I__11000 (
            .O(N__46859),
            .I(N__46697));
    InMux I__10999 (
            .O(N__46856),
            .I(N__46680));
    InMux I__10998 (
            .O(N__46855),
            .I(N__46680));
    InMux I__10997 (
            .O(N__46852),
            .I(N__46680));
    InMux I__10996 (
            .O(N__46851),
            .I(N__46680));
    InMux I__10995 (
            .O(N__46848),
            .I(N__46680));
    InMux I__10994 (
            .O(N__46847),
            .I(N__46680));
    InMux I__10993 (
            .O(N__46844),
            .I(N__46680));
    InMux I__10992 (
            .O(N__46843),
            .I(N__46680));
    InMux I__10991 (
            .O(N__46840),
            .I(N__46663));
    InMux I__10990 (
            .O(N__46839),
            .I(N__46663));
    InMux I__10989 (
            .O(N__46836),
            .I(N__46663));
    InMux I__10988 (
            .O(N__46835),
            .I(N__46663));
    InMux I__10987 (
            .O(N__46832),
            .I(N__46663));
    InMux I__10986 (
            .O(N__46831),
            .I(N__46663));
    InMux I__10985 (
            .O(N__46828),
            .I(N__46663));
    InMux I__10984 (
            .O(N__46827),
            .I(N__46663));
    CascadeMux I__10983 (
            .O(N__46826),
            .I(N__46660));
    CascadeMux I__10982 (
            .O(N__46825),
            .I(N__46656));
    CascadeMux I__10981 (
            .O(N__46824),
            .I(N__46652));
    Span4Mux_v I__10980 (
            .O(N__46819),
            .I(N__46645));
    Span4Mux_v I__10979 (
            .O(N__46816),
            .I(N__46642));
    Span4Mux_h I__10978 (
            .O(N__46813),
            .I(N__46637));
    Span4Mux_h I__10977 (
            .O(N__46808),
            .I(N__46637));
    CascadeMux I__10976 (
            .O(N__46807),
            .I(N__46634));
    CascadeMux I__10975 (
            .O(N__46806),
            .I(N__46629));
    CascadeMux I__10974 (
            .O(N__46805),
            .I(N__46625));
    CascadeMux I__10973 (
            .O(N__46804),
            .I(N__46622));
    CascadeMux I__10972 (
            .O(N__46803),
            .I(N__46619));
    CascadeMux I__10971 (
            .O(N__46802),
            .I(N__46614));
    CascadeMux I__10970 (
            .O(N__46801),
            .I(N__46610));
    CascadeMux I__10969 (
            .O(N__46800),
            .I(N__46607));
    LocalMux I__10968 (
            .O(N__46789),
            .I(N__46602));
    InMux I__10967 (
            .O(N__46788),
            .I(N__46587));
    InMux I__10966 (
            .O(N__46785),
            .I(N__46587));
    InMux I__10965 (
            .O(N__46784),
            .I(N__46587));
    InMux I__10964 (
            .O(N__46781),
            .I(N__46587));
    InMux I__10963 (
            .O(N__46780),
            .I(N__46587));
    InMux I__10962 (
            .O(N__46777),
            .I(N__46587));
    InMux I__10961 (
            .O(N__46776),
            .I(N__46587));
    InMux I__10960 (
            .O(N__46773),
            .I(N__46570));
    InMux I__10959 (
            .O(N__46772),
            .I(N__46570));
    InMux I__10958 (
            .O(N__46769),
            .I(N__46570));
    InMux I__10957 (
            .O(N__46768),
            .I(N__46570));
    InMux I__10956 (
            .O(N__46765),
            .I(N__46570));
    InMux I__10955 (
            .O(N__46764),
            .I(N__46570));
    InMux I__10954 (
            .O(N__46761),
            .I(N__46570));
    InMux I__10953 (
            .O(N__46760),
            .I(N__46570));
    CascadeMux I__10952 (
            .O(N__46759),
            .I(N__46567));
    CascadeMux I__10951 (
            .O(N__46758),
            .I(N__46563));
    CascadeMux I__10950 (
            .O(N__46757),
            .I(N__46559));
    CascadeMux I__10949 (
            .O(N__46756),
            .I(N__46555));
    Span4Mux_h I__10948 (
            .O(N__46751),
            .I(N__46543));
    Span4Mux_h I__10947 (
            .O(N__46748),
            .I(N__46543));
    Span4Mux_v I__10946 (
            .O(N__46745),
            .I(N__46543));
    LocalMux I__10945 (
            .O(N__46742),
            .I(N__46543));
    LocalMux I__10944 (
            .O(N__46725),
            .I(N__46543));
    LocalMux I__10943 (
            .O(N__46714),
            .I(N__46534));
    LocalMux I__10942 (
            .O(N__46697),
            .I(N__46534));
    LocalMux I__10941 (
            .O(N__46680),
            .I(N__46534));
    LocalMux I__10940 (
            .O(N__46663),
            .I(N__46534));
    InMux I__10939 (
            .O(N__46660),
            .I(N__46521));
    InMux I__10938 (
            .O(N__46659),
            .I(N__46521));
    InMux I__10937 (
            .O(N__46656),
            .I(N__46521));
    InMux I__10936 (
            .O(N__46655),
            .I(N__46521));
    InMux I__10935 (
            .O(N__46652),
            .I(N__46521));
    InMux I__10934 (
            .O(N__46651),
            .I(N__46521));
    CascadeMux I__10933 (
            .O(N__46650),
            .I(N__46518));
    CascadeMux I__10932 (
            .O(N__46649),
            .I(N__46514));
    CascadeMux I__10931 (
            .O(N__46648),
            .I(N__46510));
    Span4Mux_v I__10930 (
            .O(N__46645),
            .I(N__46504));
    Span4Mux_v I__10929 (
            .O(N__46642),
            .I(N__46504));
    Span4Mux_v I__10928 (
            .O(N__46637),
            .I(N__46501));
    InMux I__10927 (
            .O(N__46634),
            .I(N__46490));
    InMux I__10926 (
            .O(N__46633),
            .I(N__46490));
    InMux I__10925 (
            .O(N__46632),
            .I(N__46490));
    InMux I__10924 (
            .O(N__46629),
            .I(N__46490));
    InMux I__10923 (
            .O(N__46628),
            .I(N__46490));
    InMux I__10922 (
            .O(N__46625),
            .I(N__46483));
    InMux I__10921 (
            .O(N__46622),
            .I(N__46483));
    InMux I__10920 (
            .O(N__46619),
            .I(N__46483));
    InMux I__10919 (
            .O(N__46618),
            .I(N__46474));
    InMux I__10918 (
            .O(N__46617),
            .I(N__46474));
    InMux I__10917 (
            .O(N__46614),
            .I(N__46474));
    InMux I__10916 (
            .O(N__46613),
            .I(N__46474));
    InMux I__10915 (
            .O(N__46610),
            .I(N__46469));
    InMux I__10914 (
            .O(N__46607),
            .I(N__46469));
    InMux I__10913 (
            .O(N__46606),
            .I(N__46464));
    InMux I__10912 (
            .O(N__46605),
            .I(N__46464));
    Span4Mux_h I__10911 (
            .O(N__46602),
            .I(N__46457));
    LocalMux I__10910 (
            .O(N__46587),
            .I(N__46457));
    LocalMux I__10909 (
            .O(N__46570),
            .I(N__46457));
    InMux I__10908 (
            .O(N__46567),
            .I(N__46440));
    InMux I__10907 (
            .O(N__46566),
            .I(N__46440));
    InMux I__10906 (
            .O(N__46563),
            .I(N__46440));
    InMux I__10905 (
            .O(N__46562),
            .I(N__46440));
    InMux I__10904 (
            .O(N__46559),
            .I(N__46440));
    InMux I__10903 (
            .O(N__46558),
            .I(N__46440));
    InMux I__10902 (
            .O(N__46555),
            .I(N__46440));
    InMux I__10901 (
            .O(N__46554),
            .I(N__46440));
    Span4Mux_v I__10900 (
            .O(N__46543),
            .I(N__46433));
    Span4Mux_v I__10899 (
            .O(N__46534),
            .I(N__46433));
    LocalMux I__10898 (
            .O(N__46521),
            .I(N__46433));
    InMux I__10897 (
            .O(N__46518),
            .I(N__46420));
    InMux I__10896 (
            .O(N__46517),
            .I(N__46420));
    InMux I__10895 (
            .O(N__46514),
            .I(N__46420));
    InMux I__10894 (
            .O(N__46513),
            .I(N__46420));
    InMux I__10893 (
            .O(N__46510),
            .I(N__46420));
    InMux I__10892 (
            .O(N__46509),
            .I(N__46420));
    Odrv4 I__10891 (
            .O(N__46504),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10890 (
            .O(N__46501),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10889 (
            .O(N__46490),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10888 (
            .O(N__46483),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10887 (
            .O(N__46474),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10886 (
            .O(N__46469),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10885 (
            .O(N__46464),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10884 (
            .O(N__46457),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10883 (
            .O(N__46440),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10882 (
            .O(N__46433),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10881 (
            .O(N__46420),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    CascadeMux I__10880 (
            .O(N__46397),
            .I(N__46394));
    InMux I__10879 (
            .O(N__46394),
            .I(N__46390));
    InMux I__10878 (
            .O(N__46393),
            .I(N__46386));
    LocalMux I__10877 (
            .O(N__46390),
            .I(N__46383));
    InMux I__10876 (
            .O(N__46389),
            .I(N__46380));
    LocalMux I__10875 (
            .O(N__46386),
            .I(N__46377));
    Span4Mux_h I__10874 (
            .O(N__46383),
            .I(N__46374));
    LocalMux I__10873 (
            .O(N__46380),
            .I(N__46371));
    Odrv12 I__10872 (
            .O(N__46377),
            .I(\current_shift_inst.un4_control_input1_28 ));
    Odrv4 I__10871 (
            .O(N__46374),
            .I(\current_shift_inst.un4_control_input1_28 ));
    Odrv12 I__10870 (
            .O(N__46371),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__10869 (
            .O(N__46364),
            .I(N__46361));
    LocalMux I__10868 (
            .O(N__46361),
            .I(N__46358));
    Odrv4 I__10867 (
            .O(N__46358),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__10866 (
            .O(N__46355),
            .I(N__46352));
    LocalMux I__10865 (
            .O(N__46352),
            .I(N__46347));
    InMux I__10864 (
            .O(N__46351),
            .I(N__46344));
    InMux I__10863 (
            .O(N__46350),
            .I(N__46341));
    Span4Mux_h I__10862 (
            .O(N__46347),
            .I(N__46338));
    LocalMux I__10861 (
            .O(N__46344),
            .I(N__46335));
    LocalMux I__10860 (
            .O(N__46341),
            .I(N__46332));
    Span4Mux_v I__10859 (
            .O(N__46338),
            .I(N__46329));
    Span4Mux_h I__10858 (
            .O(N__46335),
            .I(N__46326));
    Span4Mux_h I__10857 (
            .O(N__46332),
            .I(N__46323));
    Span4Mux_v I__10856 (
            .O(N__46329),
            .I(N__46320));
    Sp12to4 I__10855 (
            .O(N__46326),
            .I(N__46317));
    Span4Mux_v I__10854 (
            .O(N__46323),
            .I(N__46314));
    Span4Mux_v I__10853 (
            .O(N__46320),
            .I(N__46311));
    Span12Mux_v I__10852 (
            .O(N__46317),
            .I(N__46308));
    Sp12to4 I__10851 (
            .O(N__46314),
            .I(N__46305));
    Span4Mux_v I__10850 (
            .O(N__46311),
            .I(N__46302));
    Span12Mux_v I__10849 (
            .O(N__46308),
            .I(N__46299));
    Span12Mux_v I__10848 (
            .O(N__46305),
            .I(N__46296));
    Span4Mux_v I__10847 (
            .O(N__46302),
            .I(N__46293));
    Odrv12 I__10846 (
            .O(N__46299),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv12 I__10845 (
            .O(N__46296),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__10844 (
            .O(N__46293),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__10843 (
            .O(N__46286),
            .I(N__46282));
    InMux I__10842 (
            .O(N__46285),
            .I(N__46279));
    LocalMux I__10841 (
            .O(N__46282),
            .I(N__46274));
    LocalMux I__10840 (
            .O(N__46279),
            .I(N__46274));
    Span12Mux_v I__10839 (
            .O(N__46274),
            .I(N__46269));
    InMux I__10838 (
            .O(N__46273),
            .I(N__46264));
    InMux I__10837 (
            .O(N__46272),
            .I(N__46264));
    Span12Mux_v I__10836 (
            .O(N__46269),
            .I(N__46261));
    LocalMux I__10835 (
            .O(N__46264),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv12 I__10834 (
            .O(N__46261),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    ClkMux I__10833 (
            .O(N__46256),
            .I(N__46253));
    GlobalMux I__10832 (
            .O(N__46253),
            .I(N__46250));
    gio2CtrlBuf I__10831 (
            .O(N__46250),
            .I(delay_tr_input_c_g));
    CascadeMux I__10830 (
            .O(N__46247),
            .I(N__46244));
    InMux I__10829 (
            .O(N__46244),
            .I(N__46240));
    InMux I__10828 (
            .O(N__46243),
            .I(N__46237));
    LocalMux I__10827 (
            .O(N__46240),
            .I(N__46234));
    LocalMux I__10826 (
            .O(N__46237),
            .I(N__46230));
    Span4Mux_v I__10825 (
            .O(N__46234),
            .I(N__46225));
    InMux I__10824 (
            .O(N__46233),
            .I(N__46222));
    Span4Mux_h I__10823 (
            .O(N__46230),
            .I(N__46218));
    InMux I__10822 (
            .O(N__46229),
            .I(N__46215));
    InMux I__10821 (
            .O(N__46228),
            .I(N__46212));
    Span4Mux_h I__10820 (
            .O(N__46225),
            .I(N__46207));
    LocalMux I__10819 (
            .O(N__46222),
            .I(N__46207));
    CascadeMux I__10818 (
            .O(N__46221),
            .I(N__46204));
    Span4Mux_h I__10817 (
            .O(N__46218),
            .I(N__46201));
    LocalMux I__10816 (
            .O(N__46215),
            .I(N__46196));
    LocalMux I__10815 (
            .O(N__46212),
            .I(N__46196));
    Span4Mux_v I__10814 (
            .O(N__46207),
            .I(N__46193));
    InMux I__10813 (
            .O(N__46204),
            .I(N__46190));
    Span4Mux_v I__10812 (
            .O(N__46201),
            .I(N__46187));
    Span4Mux_v I__10811 (
            .O(N__46196),
            .I(N__46182));
    Span4Mux_v I__10810 (
            .O(N__46193),
            .I(N__46182));
    LocalMux I__10809 (
            .O(N__46190),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__10808 (
            .O(N__46187),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__10807 (
            .O(N__46182),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    InMux I__10806 (
            .O(N__46175),
            .I(N__46172));
    LocalMux I__10805 (
            .O(N__46172),
            .I(N__46169));
    Span4Mux_v I__10804 (
            .O(N__46169),
            .I(N__46165));
    InMux I__10803 (
            .O(N__46168),
            .I(N__46162));
    Span4Mux_h I__10802 (
            .O(N__46165),
            .I(N__46159));
    LocalMux I__10801 (
            .O(N__46162),
            .I(N__46156));
    Span4Mux_v I__10800 (
            .O(N__46159),
            .I(N__46153));
    Span4Mux_h I__10799 (
            .O(N__46156),
            .I(N__46148));
    Span4Mux_v I__10798 (
            .O(N__46153),
            .I(N__46145));
    InMux I__10797 (
            .O(N__46152),
            .I(N__46140));
    InMux I__10796 (
            .O(N__46151),
            .I(N__46140));
    Odrv4 I__10795 (
            .O(N__46148),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    Odrv4 I__10794 (
            .O(N__46145),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__10793 (
            .O(N__46140),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    IoInMux I__10792 (
            .O(N__46133),
            .I(N__46130));
    LocalMux I__10791 (
            .O(N__46130),
            .I(N__46126));
    InMux I__10790 (
            .O(N__46129),
            .I(N__46123));
    Odrv12 I__10789 (
            .O(N__46126),
            .I(T23_c));
    LocalMux I__10788 (
            .O(N__46123),
            .I(T23_c));
    ClkMux I__10787 (
            .O(N__46118),
            .I(N__45731));
    ClkMux I__10786 (
            .O(N__46117),
            .I(N__45731));
    ClkMux I__10785 (
            .O(N__46116),
            .I(N__45731));
    ClkMux I__10784 (
            .O(N__46115),
            .I(N__45731));
    ClkMux I__10783 (
            .O(N__46114),
            .I(N__45731));
    ClkMux I__10782 (
            .O(N__46113),
            .I(N__45731));
    ClkMux I__10781 (
            .O(N__46112),
            .I(N__45731));
    ClkMux I__10780 (
            .O(N__46111),
            .I(N__45731));
    ClkMux I__10779 (
            .O(N__46110),
            .I(N__45731));
    ClkMux I__10778 (
            .O(N__46109),
            .I(N__45731));
    ClkMux I__10777 (
            .O(N__46108),
            .I(N__45731));
    ClkMux I__10776 (
            .O(N__46107),
            .I(N__45731));
    ClkMux I__10775 (
            .O(N__46106),
            .I(N__45731));
    ClkMux I__10774 (
            .O(N__46105),
            .I(N__45731));
    ClkMux I__10773 (
            .O(N__46104),
            .I(N__45731));
    ClkMux I__10772 (
            .O(N__46103),
            .I(N__45731));
    ClkMux I__10771 (
            .O(N__46102),
            .I(N__45731));
    ClkMux I__10770 (
            .O(N__46101),
            .I(N__45731));
    ClkMux I__10769 (
            .O(N__46100),
            .I(N__45731));
    ClkMux I__10768 (
            .O(N__46099),
            .I(N__45731));
    ClkMux I__10767 (
            .O(N__46098),
            .I(N__45731));
    ClkMux I__10766 (
            .O(N__46097),
            .I(N__45731));
    ClkMux I__10765 (
            .O(N__46096),
            .I(N__45731));
    ClkMux I__10764 (
            .O(N__46095),
            .I(N__45731));
    ClkMux I__10763 (
            .O(N__46094),
            .I(N__45731));
    ClkMux I__10762 (
            .O(N__46093),
            .I(N__45731));
    ClkMux I__10761 (
            .O(N__46092),
            .I(N__45731));
    ClkMux I__10760 (
            .O(N__46091),
            .I(N__45731));
    ClkMux I__10759 (
            .O(N__46090),
            .I(N__45731));
    ClkMux I__10758 (
            .O(N__46089),
            .I(N__45731));
    ClkMux I__10757 (
            .O(N__46088),
            .I(N__45731));
    ClkMux I__10756 (
            .O(N__46087),
            .I(N__45731));
    ClkMux I__10755 (
            .O(N__46086),
            .I(N__45731));
    ClkMux I__10754 (
            .O(N__46085),
            .I(N__45731));
    ClkMux I__10753 (
            .O(N__46084),
            .I(N__45731));
    ClkMux I__10752 (
            .O(N__46083),
            .I(N__45731));
    ClkMux I__10751 (
            .O(N__46082),
            .I(N__45731));
    ClkMux I__10750 (
            .O(N__46081),
            .I(N__45731));
    ClkMux I__10749 (
            .O(N__46080),
            .I(N__45731));
    ClkMux I__10748 (
            .O(N__46079),
            .I(N__45731));
    ClkMux I__10747 (
            .O(N__46078),
            .I(N__45731));
    ClkMux I__10746 (
            .O(N__46077),
            .I(N__45731));
    ClkMux I__10745 (
            .O(N__46076),
            .I(N__45731));
    ClkMux I__10744 (
            .O(N__46075),
            .I(N__45731));
    ClkMux I__10743 (
            .O(N__46074),
            .I(N__45731));
    ClkMux I__10742 (
            .O(N__46073),
            .I(N__45731));
    ClkMux I__10741 (
            .O(N__46072),
            .I(N__45731));
    ClkMux I__10740 (
            .O(N__46071),
            .I(N__45731));
    ClkMux I__10739 (
            .O(N__46070),
            .I(N__45731));
    ClkMux I__10738 (
            .O(N__46069),
            .I(N__45731));
    ClkMux I__10737 (
            .O(N__46068),
            .I(N__45731));
    ClkMux I__10736 (
            .O(N__46067),
            .I(N__45731));
    ClkMux I__10735 (
            .O(N__46066),
            .I(N__45731));
    ClkMux I__10734 (
            .O(N__46065),
            .I(N__45731));
    ClkMux I__10733 (
            .O(N__46064),
            .I(N__45731));
    ClkMux I__10732 (
            .O(N__46063),
            .I(N__45731));
    ClkMux I__10731 (
            .O(N__46062),
            .I(N__45731));
    ClkMux I__10730 (
            .O(N__46061),
            .I(N__45731));
    ClkMux I__10729 (
            .O(N__46060),
            .I(N__45731));
    ClkMux I__10728 (
            .O(N__46059),
            .I(N__45731));
    ClkMux I__10727 (
            .O(N__46058),
            .I(N__45731));
    ClkMux I__10726 (
            .O(N__46057),
            .I(N__45731));
    ClkMux I__10725 (
            .O(N__46056),
            .I(N__45731));
    ClkMux I__10724 (
            .O(N__46055),
            .I(N__45731));
    ClkMux I__10723 (
            .O(N__46054),
            .I(N__45731));
    ClkMux I__10722 (
            .O(N__46053),
            .I(N__45731));
    ClkMux I__10721 (
            .O(N__46052),
            .I(N__45731));
    ClkMux I__10720 (
            .O(N__46051),
            .I(N__45731));
    ClkMux I__10719 (
            .O(N__46050),
            .I(N__45731));
    ClkMux I__10718 (
            .O(N__46049),
            .I(N__45731));
    ClkMux I__10717 (
            .O(N__46048),
            .I(N__45731));
    ClkMux I__10716 (
            .O(N__46047),
            .I(N__45731));
    ClkMux I__10715 (
            .O(N__46046),
            .I(N__45731));
    ClkMux I__10714 (
            .O(N__46045),
            .I(N__45731));
    ClkMux I__10713 (
            .O(N__46044),
            .I(N__45731));
    ClkMux I__10712 (
            .O(N__46043),
            .I(N__45731));
    ClkMux I__10711 (
            .O(N__46042),
            .I(N__45731));
    ClkMux I__10710 (
            .O(N__46041),
            .I(N__45731));
    ClkMux I__10709 (
            .O(N__46040),
            .I(N__45731));
    ClkMux I__10708 (
            .O(N__46039),
            .I(N__45731));
    ClkMux I__10707 (
            .O(N__46038),
            .I(N__45731));
    ClkMux I__10706 (
            .O(N__46037),
            .I(N__45731));
    ClkMux I__10705 (
            .O(N__46036),
            .I(N__45731));
    ClkMux I__10704 (
            .O(N__46035),
            .I(N__45731));
    ClkMux I__10703 (
            .O(N__46034),
            .I(N__45731));
    ClkMux I__10702 (
            .O(N__46033),
            .I(N__45731));
    ClkMux I__10701 (
            .O(N__46032),
            .I(N__45731));
    ClkMux I__10700 (
            .O(N__46031),
            .I(N__45731));
    ClkMux I__10699 (
            .O(N__46030),
            .I(N__45731));
    ClkMux I__10698 (
            .O(N__46029),
            .I(N__45731));
    ClkMux I__10697 (
            .O(N__46028),
            .I(N__45731));
    ClkMux I__10696 (
            .O(N__46027),
            .I(N__45731));
    ClkMux I__10695 (
            .O(N__46026),
            .I(N__45731));
    ClkMux I__10694 (
            .O(N__46025),
            .I(N__45731));
    ClkMux I__10693 (
            .O(N__46024),
            .I(N__45731));
    ClkMux I__10692 (
            .O(N__46023),
            .I(N__45731));
    ClkMux I__10691 (
            .O(N__46022),
            .I(N__45731));
    ClkMux I__10690 (
            .O(N__46021),
            .I(N__45731));
    ClkMux I__10689 (
            .O(N__46020),
            .I(N__45731));
    ClkMux I__10688 (
            .O(N__46019),
            .I(N__45731));
    ClkMux I__10687 (
            .O(N__46018),
            .I(N__45731));
    ClkMux I__10686 (
            .O(N__46017),
            .I(N__45731));
    ClkMux I__10685 (
            .O(N__46016),
            .I(N__45731));
    ClkMux I__10684 (
            .O(N__46015),
            .I(N__45731));
    ClkMux I__10683 (
            .O(N__46014),
            .I(N__45731));
    ClkMux I__10682 (
            .O(N__46013),
            .I(N__45731));
    ClkMux I__10681 (
            .O(N__46012),
            .I(N__45731));
    ClkMux I__10680 (
            .O(N__46011),
            .I(N__45731));
    ClkMux I__10679 (
            .O(N__46010),
            .I(N__45731));
    ClkMux I__10678 (
            .O(N__46009),
            .I(N__45731));
    ClkMux I__10677 (
            .O(N__46008),
            .I(N__45731));
    ClkMux I__10676 (
            .O(N__46007),
            .I(N__45731));
    ClkMux I__10675 (
            .O(N__46006),
            .I(N__45731));
    ClkMux I__10674 (
            .O(N__46005),
            .I(N__45731));
    ClkMux I__10673 (
            .O(N__46004),
            .I(N__45731));
    ClkMux I__10672 (
            .O(N__46003),
            .I(N__45731));
    ClkMux I__10671 (
            .O(N__46002),
            .I(N__45731));
    ClkMux I__10670 (
            .O(N__46001),
            .I(N__45731));
    ClkMux I__10669 (
            .O(N__46000),
            .I(N__45731));
    ClkMux I__10668 (
            .O(N__45999),
            .I(N__45731));
    ClkMux I__10667 (
            .O(N__45998),
            .I(N__45731));
    ClkMux I__10666 (
            .O(N__45997),
            .I(N__45731));
    ClkMux I__10665 (
            .O(N__45996),
            .I(N__45731));
    ClkMux I__10664 (
            .O(N__45995),
            .I(N__45731));
    ClkMux I__10663 (
            .O(N__45994),
            .I(N__45731));
    ClkMux I__10662 (
            .O(N__45993),
            .I(N__45731));
    ClkMux I__10661 (
            .O(N__45992),
            .I(N__45731));
    ClkMux I__10660 (
            .O(N__45991),
            .I(N__45731));
    ClkMux I__10659 (
            .O(N__45990),
            .I(N__45731));
    GlobalMux I__10658 (
            .O(N__45731),
            .I(clk_100mhz_0));
    InMux I__10657 (
            .O(N__45728),
            .I(N__45711));
    InMux I__10656 (
            .O(N__45727),
            .I(N__45708));
    InMux I__10655 (
            .O(N__45726),
            .I(N__45705));
    InMux I__10654 (
            .O(N__45725),
            .I(N__45702));
    InMux I__10653 (
            .O(N__45724),
            .I(N__45699));
    InMux I__10652 (
            .O(N__45723),
            .I(N__45694));
    InMux I__10651 (
            .O(N__45722),
            .I(N__45694));
    InMux I__10650 (
            .O(N__45721),
            .I(N__45691));
    InMux I__10649 (
            .O(N__45720),
            .I(N__45686));
    InMux I__10648 (
            .O(N__45719),
            .I(N__45686));
    InMux I__10647 (
            .O(N__45718),
            .I(N__45683));
    InMux I__10646 (
            .O(N__45717),
            .I(N__45678));
    InMux I__10645 (
            .O(N__45716),
            .I(N__45678));
    InMux I__10644 (
            .O(N__45715),
            .I(N__45675));
    InMux I__10643 (
            .O(N__45714),
            .I(N__45672));
    LocalMux I__10642 (
            .O(N__45711),
            .I(N__45669));
    LocalMux I__10641 (
            .O(N__45708),
            .I(N__45666));
    LocalMux I__10640 (
            .O(N__45705),
            .I(N__45663));
    LocalMux I__10639 (
            .O(N__45702),
            .I(N__45659));
    LocalMux I__10638 (
            .O(N__45699),
            .I(N__45646));
    LocalMux I__10637 (
            .O(N__45694),
            .I(N__45643));
    LocalMux I__10636 (
            .O(N__45691),
            .I(N__45627));
    LocalMux I__10635 (
            .O(N__45686),
            .I(N__45616));
    LocalMux I__10634 (
            .O(N__45683),
            .I(N__45613));
    LocalMux I__10633 (
            .O(N__45678),
            .I(N__45523));
    LocalMux I__10632 (
            .O(N__45675),
            .I(N__45520));
    LocalMux I__10631 (
            .O(N__45672),
            .I(N__45516));
    Glb2LocalMux I__10630 (
            .O(N__45669),
            .I(N__45245));
    Glb2LocalMux I__10629 (
            .O(N__45666),
            .I(N__45245));
    Glb2LocalMux I__10628 (
            .O(N__45663),
            .I(N__45245));
    SRMux I__10627 (
            .O(N__45662),
            .I(N__45245));
    Glb2LocalMux I__10626 (
            .O(N__45659),
            .I(N__45245));
    SRMux I__10625 (
            .O(N__45658),
            .I(N__45245));
    SRMux I__10624 (
            .O(N__45657),
            .I(N__45245));
    SRMux I__10623 (
            .O(N__45656),
            .I(N__45245));
    SRMux I__10622 (
            .O(N__45655),
            .I(N__45245));
    SRMux I__10621 (
            .O(N__45654),
            .I(N__45245));
    SRMux I__10620 (
            .O(N__45653),
            .I(N__45245));
    SRMux I__10619 (
            .O(N__45652),
            .I(N__45245));
    SRMux I__10618 (
            .O(N__45651),
            .I(N__45245));
    SRMux I__10617 (
            .O(N__45650),
            .I(N__45245));
    SRMux I__10616 (
            .O(N__45649),
            .I(N__45245));
    Glb2LocalMux I__10615 (
            .O(N__45646),
            .I(N__45245));
    Glb2LocalMux I__10614 (
            .O(N__45643),
            .I(N__45245));
    SRMux I__10613 (
            .O(N__45642),
            .I(N__45245));
    SRMux I__10612 (
            .O(N__45641),
            .I(N__45245));
    SRMux I__10611 (
            .O(N__45640),
            .I(N__45245));
    SRMux I__10610 (
            .O(N__45639),
            .I(N__45245));
    SRMux I__10609 (
            .O(N__45638),
            .I(N__45245));
    SRMux I__10608 (
            .O(N__45637),
            .I(N__45245));
    SRMux I__10607 (
            .O(N__45636),
            .I(N__45245));
    SRMux I__10606 (
            .O(N__45635),
            .I(N__45245));
    SRMux I__10605 (
            .O(N__45634),
            .I(N__45245));
    SRMux I__10604 (
            .O(N__45633),
            .I(N__45245));
    SRMux I__10603 (
            .O(N__45632),
            .I(N__45245));
    SRMux I__10602 (
            .O(N__45631),
            .I(N__45245));
    SRMux I__10601 (
            .O(N__45630),
            .I(N__45245));
    Glb2LocalMux I__10600 (
            .O(N__45627),
            .I(N__45245));
    SRMux I__10599 (
            .O(N__45626),
            .I(N__45245));
    SRMux I__10598 (
            .O(N__45625),
            .I(N__45245));
    SRMux I__10597 (
            .O(N__45624),
            .I(N__45245));
    SRMux I__10596 (
            .O(N__45623),
            .I(N__45245));
    SRMux I__10595 (
            .O(N__45622),
            .I(N__45245));
    SRMux I__10594 (
            .O(N__45621),
            .I(N__45245));
    SRMux I__10593 (
            .O(N__45620),
            .I(N__45245));
    SRMux I__10592 (
            .O(N__45619),
            .I(N__45245));
    Glb2LocalMux I__10591 (
            .O(N__45616),
            .I(N__45245));
    Glb2LocalMux I__10590 (
            .O(N__45613),
            .I(N__45245));
    SRMux I__10589 (
            .O(N__45612),
            .I(N__45245));
    SRMux I__10588 (
            .O(N__45611),
            .I(N__45245));
    SRMux I__10587 (
            .O(N__45610),
            .I(N__45245));
    SRMux I__10586 (
            .O(N__45609),
            .I(N__45245));
    SRMux I__10585 (
            .O(N__45608),
            .I(N__45245));
    SRMux I__10584 (
            .O(N__45607),
            .I(N__45245));
    SRMux I__10583 (
            .O(N__45606),
            .I(N__45245));
    SRMux I__10582 (
            .O(N__45605),
            .I(N__45245));
    SRMux I__10581 (
            .O(N__45604),
            .I(N__45245));
    SRMux I__10580 (
            .O(N__45603),
            .I(N__45245));
    SRMux I__10579 (
            .O(N__45602),
            .I(N__45245));
    SRMux I__10578 (
            .O(N__45601),
            .I(N__45245));
    SRMux I__10577 (
            .O(N__45600),
            .I(N__45245));
    SRMux I__10576 (
            .O(N__45599),
            .I(N__45245));
    SRMux I__10575 (
            .O(N__45598),
            .I(N__45245));
    SRMux I__10574 (
            .O(N__45597),
            .I(N__45245));
    SRMux I__10573 (
            .O(N__45596),
            .I(N__45245));
    SRMux I__10572 (
            .O(N__45595),
            .I(N__45245));
    SRMux I__10571 (
            .O(N__45594),
            .I(N__45245));
    SRMux I__10570 (
            .O(N__45593),
            .I(N__45245));
    SRMux I__10569 (
            .O(N__45592),
            .I(N__45245));
    SRMux I__10568 (
            .O(N__45591),
            .I(N__45245));
    SRMux I__10567 (
            .O(N__45590),
            .I(N__45245));
    SRMux I__10566 (
            .O(N__45589),
            .I(N__45245));
    SRMux I__10565 (
            .O(N__45588),
            .I(N__45245));
    SRMux I__10564 (
            .O(N__45587),
            .I(N__45245));
    SRMux I__10563 (
            .O(N__45586),
            .I(N__45245));
    SRMux I__10562 (
            .O(N__45585),
            .I(N__45245));
    SRMux I__10561 (
            .O(N__45584),
            .I(N__45245));
    SRMux I__10560 (
            .O(N__45583),
            .I(N__45245));
    SRMux I__10559 (
            .O(N__45582),
            .I(N__45245));
    SRMux I__10558 (
            .O(N__45581),
            .I(N__45245));
    SRMux I__10557 (
            .O(N__45580),
            .I(N__45245));
    SRMux I__10556 (
            .O(N__45579),
            .I(N__45245));
    SRMux I__10555 (
            .O(N__45578),
            .I(N__45245));
    SRMux I__10554 (
            .O(N__45577),
            .I(N__45245));
    SRMux I__10553 (
            .O(N__45576),
            .I(N__45245));
    SRMux I__10552 (
            .O(N__45575),
            .I(N__45245));
    SRMux I__10551 (
            .O(N__45574),
            .I(N__45245));
    SRMux I__10550 (
            .O(N__45573),
            .I(N__45245));
    SRMux I__10549 (
            .O(N__45572),
            .I(N__45245));
    SRMux I__10548 (
            .O(N__45571),
            .I(N__45245));
    SRMux I__10547 (
            .O(N__45570),
            .I(N__45245));
    SRMux I__10546 (
            .O(N__45569),
            .I(N__45245));
    SRMux I__10545 (
            .O(N__45568),
            .I(N__45245));
    SRMux I__10544 (
            .O(N__45567),
            .I(N__45245));
    SRMux I__10543 (
            .O(N__45566),
            .I(N__45245));
    SRMux I__10542 (
            .O(N__45565),
            .I(N__45245));
    SRMux I__10541 (
            .O(N__45564),
            .I(N__45245));
    SRMux I__10540 (
            .O(N__45563),
            .I(N__45245));
    SRMux I__10539 (
            .O(N__45562),
            .I(N__45245));
    SRMux I__10538 (
            .O(N__45561),
            .I(N__45245));
    SRMux I__10537 (
            .O(N__45560),
            .I(N__45245));
    SRMux I__10536 (
            .O(N__45559),
            .I(N__45245));
    SRMux I__10535 (
            .O(N__45558),
            .I(N__45245));
    SRMux I__10534 (
            .O(N__45557),
            .I(N__45245));
    SRMux I__10533 (
            .O(N__45556),
            .I(N__45245));
    SRMux I__10532 (
            .O(N__45555),
            .I(N__45245));
    SRMux I__10531 (
            .O(N__45554),
            .I(N__45245));
    SRMux I__10530 (
            .O(N__45553),
            .I(N__45245));
    SRMux I__10529 (
            .O(N__45552),
            .I(N__45245));
    SRMux I__10528 (
            .O(N__45551),
            .I(N__45245));
    SRMux I__10527 (
            .O(N__45550),
            .I(N__45245));
    SRMux I__10526 (
            .O(N__45549),
            .I(N__45245));
    SRMux I__10525 (
            .O(N__45548),
            .I(N__45245));
    SRMux I__10524 (
            .O(N__45547),
            .I(N__45245));
    SRMux I__10523 (
            .O(N__45546),
            .I(N__45245));
    SRMux I__10522 (
            .O(N__45545),
            .I(N__45245));
    SRMux I__10521 (
            .O(N__45544),
            .I(N__45245));
    SRMux I__10520 (
            .O(N__45543),
            .I(N__45245));
    SRMux I__10519 (
            .O(N__45542),
            .I(N__45245));
    SRMux I__10518 (
            .O(N__45541),
            .I(N__45245));
    SRMux I__10517 (
            .O(N__45540),
            .I(N__45245));
    SRMux I__10516 (
            .O(N__45539),
            .I(N__45245));
    SRMux I__10515 (
            .O(N__45538),
            .I(N__45245));
    SRMux I__10514 (
            .O(N__45537),
            .I(N__45245));
    SRMux I__10513 (
            .O(N__45536),
            .I(N__45245));
    SRMux I__10512 (
            .O(N__45535),
            .I(N__45245));
    SRMux I__10511 (
            .O(N__45534),
            .I(N__45245));
    SRMux I__10510 (
            .O(N__45533),
            .I(N__45245));
    SRMux I__10509 (
            .O(N__45532),
            .I(N__45245));
    SRMux I__10508 (
            .O(N__45531),
            .I(N__45245));
    SRMux I__10507 (
            .O(N__45530),
            .I(N__45245));
    SRMux I__10506 (
            .O(N__45529),
            .I(N__45245));
    SRMux I__10505 (
            .O(N__45528),
            .I(N__45245));
    SRMux I__10504 (
            .O(N__45527),
            .I(N__45245));
    SRMux I__10503 (
            .O(N__45526),
            .I(N__45245));
    Glb2LocalMux I__10502 (
            .O(N__45523),
            .I(N__45245));
    Glb2LocalMux I__10501 (
            .O(N__45520),
            .I(N__45245));
    SRMux I__10500 (
            .O(N__45519),
            .I(N__45245));
    Glb2LocalMux I__10499 (
            .O(N__45516),
            .I(N__45245));
    SRMux I__10498 (
            .O(N__45515),
            .I(N__45245));
    SRMux I__10497 (
            .O(N__45514),
            .I(N__45245));
    GlobalMux I__10496 (
            .O(N__45245),
            .I(N__45242));
    gio2CtrlBuf I__10495 (
            .O(N__45242),
            .I(red_c_g));
    CascadeMux I__10494 (
            .O(N__45239),
            .I(N__45235));
    CascadeMux I__10493 (
            .O(N__45238),
            .I(N__45232));
    InMux I__10492 (
            .O(N__45235),
            .I(N__45229));
    InMux I__10491 (
            .O(N__45232),
            .I(N__45225));
    LocalMux I__10490 (
            .O(N__45229),
            .I(N__45221));
    InMux I__10489 (
            .O(N__45228),
            .I(N__45218));
    LocalMux I__10488 (
            .O(N__45225),
            .I(N__45215));
    InMux I__10487 (
            .O(N__45224),
            .I(N__45212));
    Span4Mux_h I__10486 (
            .O(N__45221),
            .I(N__45209));
    LocalMux I__10485 (
            .O(N__45218),
            .I(N__45206));
    Span4Mux_h I__10484 (
            .O(N__45215),
            .I(N__45201));
    LocalMux I__10483 (
            .O(N__45212),
            .I(N__45201));
    Span4Mux_v I__10482 (
            .O(N__45209),
            .I(N__45196));
    Span4Mux_h I__10481 (
            .O(N__45206),
            .I(N__45196));
    Odrv4 I__10480 (
            .O(N__45201),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__10479 (
            .O(N__45196),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__10478 (
            .O(N__45191),
            .I(N__45187));
    InMux I__10477 (
            .O(N__45190),
            .I(N__45184));
    LocalMux I__10476 (
            .O(N__45187),
            .I(N__45180));
    LocalMux I__10475 (
            .O(N__45184),
            .I(N__45177));
    InMux I__10474 (
            .O(N__45183),
            .I(N__45174));
    Odrv12 I__10473 (
            .O(N__45180),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv4 I__10472 (
            .O(N__45177),
            .I(\current_shift_inst.un4_control_input1_17 ));
    LocalMux I__10471 (
            .O(N__45174),
            .I(\current_shift_inst.un4_control_input1_17 ));
    CascadeMux I__10470 (
            .O(N__45167),
            .I(N__45164));
    InMux I__10469 (
            .O(N__45164),
            .I(N__45161));
    LocalMux I__10468 (
            .O(N__45161),
            .I(N__45158));
    Odrv12 I__10467 (
            .O(N__45158),
            .I(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ));
    CascadeMux I__10466 (
            .O(N__45155),
            .I(N__45151));
    CascadeMux I__10465 (
            .O(N__45154),
            .I(N__45148));
    InMux I__10464 (
            .O(N__45151),
            .I(N__45145));
    InMux I__10463 (
            .O(N__45148),
            .I(N__45142));
    LocalMux I__10462 (
            .O(N__45145),
            .I(N__45138));
    LocalMux I__10461 (
            .O(N__45142),
            .I(N__45135));
    InMux I__10460 (
            .O(N__45141),
            .I(N__45132));
    Span4Mux_h I__10459 (
            .O(N__45138),
            .I(N__45126));
    Span4Mux_v I__10458 (
            .O(N__45135),
            .I(N__45126));
    LocalMux I__10457 (
            .O(N__45132),
            .I(N__45123));
    InMux I__10456 (
            .O(N__45131),
            .I(N__45120));
    Odrv4 I__10455 (
            .O(N__45126),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv12 I__10454 (
            .O(N__45123),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__10453 (
            .O(N__45120),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__10452 (
            .O(N__45113),
            .I(N__45109));
    InMux I__10451 (
            .O(N__45112),
            .I(N__45106));
    LocalMux I__10450 (
            .O(N__45109),
            .I(N__45102));
    LocalMux I__10449 (
            .O(N__45106),
            .I(N__45099));
    InMux I__10448 (
            .O(N__45105),
            .I(N__45096));
    Odrv12 I__10447 (
            .O(N__45102),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__10446 (
            .O(N__45099),
            .I(\current_shift_inst.un4_control_input1_12 ));
    LocalMux I__10445 (
            .O(N__45096),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__10444 (
            .O(N__45089),
            .I(N__45086));
    LocalMux I__10443 (
            .O(N__45086),
            .I(N__45083));
    Odrv4 I__10442 (
            .O(N__45083),
            .I(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ));
    InMux I__10441 (
            .O(N__45080),
            .I(N__45076));
    InMux I__10440 (
            .O(N__45079),
            .I(N__45072));
    LocalMux I__10439 (
            .O(N__45076),
            .I(N__45069));
    InMux I__10438 (
            .O(N__45075),
            .I(N__45066));
    LocalMux I__10437 (
            .O(N__45072),
            .I(N__45061));
    Span4Mux_v I__10436 (
            .O(N__45069),
            .I(N__45061));
    LocalMux I__10435 (
            .O(N__45066),
            .I(N__45057));
    Span4Mux_h I__10434 (
            .O(N__45061),
            .I(N__45054));
    InMux I__10433 (
            .O(N__45060),
            .I(N__45051));
    Span4Mux_h I__10432 (
            .O(N__45057),
            .I(N__45048));
    Odrv4 I__10431 (
            .O(N__45054),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    LocalMux I__10430 (
            .O(N__45051),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv4 I__10429 (
            .O(N__45048),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    CascadeMux I__10428 (
            .O(N__45041),
            .I(N__45038));
    InMux I__10427 (
            .O(N__45038),
            .I(N__45033));
    InMux I__10426 (
            .O(N__45037),
            .I(N__45030));
    InMux I__10425 (
            .O(N__45036),
            .I(N__45027));
    LocalMux I__10424 (
            .O(N__45033),
            .I(N__45024));
    LocalMux I__10423 (
            .O(N__45030),
            .I(N__45021));
    LocalMux I__10422 (
            .O(N__45027),
            .I(N__45018));
    Span4Mux_h I__10421 (
            .O(N__45024),
            .I(N__45015));
    Span4Mux_h I__10420 (
            .O(N__45021),
            .I(N__45012));
    Odrv4 I__10419 (
            .O(N__45018),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__10418 (
            .O(N__45015),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__10417 (
            .O(N__45012),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__10416 (
            .O(N__45005),
            .I(N__45002));
    LocalMux I__10415 (
            .O(N__45002),
            .I(N__44999));
    Odrv4 I__10414 (
            .O(N__44999),
            .I(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ));
    CascadeMux I__10413 (
            .O(N__44996),
            .I(N__44993));
    InMux I__10412 (
            .O(N__44993),
            .I(N__44990));
    LocalMux I__10411 (
            .O(N__44990),
            .I(N__44987));
    Span4Mux_h I__10410 (
            .O(N__44987),
            .I(N__44983));
    InMux I__10409 (
            .O(N__44986),
            .I(N__44980));
    Span4Mux_v I__10408 (
            .O(N__44983),
            .I(N__44975));
    LocalMux I__10407 (
            .O(N__44980),
            .I(N__44972));
    InMux I__10406 (
            .O(N__44979),
            .I(N__44969));
    InMux I__10405 (
            .O(N__44978),
            .I(N__44966));
    Odrv4 I__10404 (
            .O(N__44975),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv12 I__10403 (
            .O(N__44972),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__10402 (
            .O(N__44969),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__10401 (
            .O(N__44966),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__10400 (
            .O(N__44957),
            .I(N__44954));
    LocalMux I__10399 (
            .O(N__44954),
            .I(N__44949));
    InMux I__10398 (
            .O(N__44953),
            .I(N__44946));
    CascadeMux I__10397 (
            .O(N__44952),
            .I(N__44943));
    Span4Mux_v I__10396 (
            .O(N__44949),
            .I(N__44938));
    LocalMux I__10395 (
            .O(N__44946),
            .I(N__44938));
    InMux I__10394 (
            .O(N__44943),
            .I(N__44935));
    Span4Mux_h I__10393 (
            .O(N__44938),
            .I(N__44932));
    LocalMux I__10392 (
            .O(N__44935),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv4 I__10391 (
            .O(N__44932),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__10390 (
            .O(N__44927),
            .I(N__44924));
    LocalMux I__10389 (
            .O(N__44924),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    CascadeMux I__10388 (
            .O(N__44921),
            .I(N__44918));
    InMux I__10387 (
            .O(N__44918),
            .I(N__44912));
    InMux I__10386 (
            .O(N__44917),
            .I(N__44905));
    InMux I__10385 (
            .O(N__44916),
            .I(N__44905));
    InMux I__10384 (
            .O(N__44915),
            .I(N__44905));
    LocalMux I__10383 (
            .O(N__44912),
            .I(N__44902));
    LocalMux I__10382 (
            .O(N__44905),
            .I(N__44899));
    Span4Mux_v I__10381 (
            .O(N__44902),
            .I(N__44896));
    Span4Mux_h I__10380 (
            .O(N__44899),
            .I(N__44893));
    Span4Mux_v I__10379 (
            .O(N__44896),
            .I(N__44888));
    Span4Mux_v I__10378 (
            .O(N__44893),
            .I(N__44888));
    Odrv4 I__10377 (
            .O(N__44888),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__10376 (
            .O(N__44885),
            .I(N__44882));
    LocalMux I__10375 (
            .O(N__44882),
            .I(N__44879));
    Span4Mux_h I__10374 (
            .O(N__44879),
            .I(N__44874));
    InMux I__10373 (
            .O(N__44878),
            .I(N__44869));
    InMux I__10372 (
            .O(N__44877),
            .I(N__44869));
    Odrv4 I__10371 (
            .O(N__44874),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__10370 (
            .O(N__44869),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__10369 (
            .O(N__44864),
            .I(N__44861));
    LocalMux I__10368 (
            .O(N__44861),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    CascadeMux I__10367 (
            .O(N__44858),
            .I(N__44854));
    CascadeMux I__10366 (
            .O(N__44857),
            .I(N__44851));
    InMux I__10365 (
            .O(N__44854),
            .I(N__44848));
    InMux I__10364 (
            .O(N__44851),
            .I(N__44845));
    LocalMux I__10363 (
            .O(N__44848),
            .I(N__44842));
    LocalMux I__10362 (
            .O(N__44845),
            .I(N__44837));
    Span4Mux_v I__10361 (
            .O(N__44842),
            .I(N__44834));
    InMux I__10360 (
            .O(N__44841),
            .I(N__44831));
    InMux I__10359 (
            .O(N__44840),
            .I(N__44828));
    Odrv12 I__10358 (
            .O(N__44837),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__10357 (
            .O(N__44834),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__10356 (
            .O(N__44831),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__10355 (
            .O(N__44828),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__10354 (
            .O(N__44819),
            .I(N__44815));
    InMux I__10353 (
            .O(N__44818),
            .I(N__44812));
    LocalMux I__10352 (
            .O(N__44815),
            .I(N__44808));
    LocalMux I__10351 (
            .O(N__44812),
            .I(N__44805));
    InMux I__10350 (
            .O(N__44811),
            .I(N__44802));
    Span4Mux_h I__10349 (
            .O(N__44808),
            .I(N__44797));
    Span4Mux_v I__10348 (
            .O(N__44805),
            .I(N__44797));
    LocalMux I__10347 (
            .O(N__44802),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv4 I__10346 (
            .O(N__44797),
            .I(\current_shift_inst.un4_control_input1_25 ));
    CascadeMux I__10345 (
            .O(N__44792),
            .I(N__44789));
    InMux I__10344 (
            .O(N__44789),
            .I(N__44786));
    LocalMux I__10343 (
            .O(N__44786),
            .I(N__44783));
    Odrv4 I__10342 (
            .O(N__44783),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    CascadeMux I__10341 (
            .O(N__44780),
            .I(N__44777));
    InMux I__10340 (
            .O(N__44777),
            .I(N__44772));
    CascadeMux I__10339 (
            .O(N__44776),
            .I(N__44769));
    InMux I__10338 (
            .O(N__44775),
            .I(N__44766));
    LocalMux I__10337 (
            .O(N__44772),
            .I(N__44763));
    InMux I__10336 (
            .O(N__44769),
            .I(N__44760));
    LocalMux I__10335 (
            .O(N__44766),
            .I(N__44757));
    Span12Mux_v I__10334 (
            .O(N__44763),
            .I(N__44753));
    LocalMux I__10333 (
            .O(N__44760),
            .I(N__44750));
    Span4Mux_v I__10332 (
            .O(N__44757),
            .I(N__44747));
    InMux I__10331 (
            .O(N__44756),
            .I(N__44744));
    Odrv12 I__10330 (
            .O(N__44753),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv12 I__10329 (
            .O(N__44750),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__10328 (
            .O(N__44747),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    LocalMux I__10327 (
            .O(N__44744),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__10326 (
            .O(N__44735),
            .I(N__44730));
    InMux I__10325 (
            .O(N__44734),
            .I(N__44727));
    InMux I__10324 (
            .O(N__44733),
            .I(N__44724));
    LocalMux I__10323 (
            .O(N__44730),
            .I(N__44719));
    LocalMux I__10322 (
            .O(N__44727),
            .I(N__44719));
    LocalMux I__10321 (
            .O(N__44724),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv12 I__10320 (
            .O(N__44719),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__10319 (
            .O(N__44714),
            .I(N__44711));
    LocalMux I__10318 (
            .O(N__44711),
            .I(N__44708));
    Odrv4 I__10317 (
            .O(N__44708),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    CascadeMux I__10316 (
            .O(N__44705),
            .I(N__44702));
    InMux I__10315 (
            .O(N__44702),
            .I(N__44699));
    LocalMux I__10314 (
            .O(N__44699),
            .I(N__44694));
    InMux I__10313 (
            .O(N__44698),
            .I(N__44691));
    InMux I__10312 (
            .O(N__44697),
            .I(N__44688));
    Odrv12 I__10311 (
            .O(N__44694),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__10310 (
            .O(N__44691),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__10309 (
            .O(N__44688),
            .I(\current_shift_inst.un4_control_input1_21 ));
    InMux I__10308 (
            .O(N__44681),
            .I(N__44676));
    InMux I__10307 (
            .O(N__44680),
            .I(N__44673));
    InMux I__10306 (
            .O(N__44679),
            .I(N__44670));
    LocalMux I__10305 (
            .O(N__44676),
            .I(N__44667));
    LocalMux I__10304 (
            .O(N__44673),
            .I(N__44664));
    LocalMux I__10303 (
            .O(N__44670),
            .I(N__44660));
    Span4Mux_v I__10302 (
            .O(N__44667),
            .I(N__44655));
    Span4Mux_v I__10301 (
            .O(N__44664),
            .I(N__44655));
    InMux I__10300 (
            .O(N__44663),
            .I(N__44652));
    Odrv4 I__10299 (
            .O(N__44660),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__10298 (
            .O(N__44655),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    LocalMux I__10297 (
            .O(N__44652),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    CascadeMux I__10296 (
            .O(N__44645),
            .I(N__44642));
    InMux I__10295 (
            .O(N__44642),
            .I(N__44639));
    LocalMux I__10294 (
            .O(N__44639),
            .I(N__44636));
    Span4Mux_h I__10293 (
            .O(N__44636),
            .I(N__44633));
    Odrv4 I__10292 (
            .O(N__44633),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    InMux I__10291 (
            .O(N__44630),
            .I(N__44627));
    LocalMux I__10290 (
            .O(N__44627),
            .I(N__44624));
    Span4Mux_h I__10289 (
            .O(N__44624),
            .I(N__44621));
    Odrv4 I__10288 (
            .O(N__44621),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__10287 (
            .O(N__44618),
            .I(bfn_18_17_0_));
    InMux I__10286 (
            .O(N__44615),
            .I(N__44612));
    LocalMux I__10285 (
            .O(N__44612),
            .I(N__44609));
    Span4Mux_h I__10284 (
            .O(N__44609),
            .I(N__44606));
    Odrv4 I__10283 (
            .O(N__44606),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__10282 (
            .O(N__44603),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    CascadeMux I__10281 (
            .O(N__44600),
            .I(N__44597));
    InMux I__10280 (
            .O(N__44597),
            .I(N__44594));
    LocalMux I__10279 (
            .O(N__44594),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__10278 (
            .O(N__44591),
            .I(N__44588));
    LocalMux I__10277 (
            .O(N__44588),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__10276 (
            .O(N__44585),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__10275 (
            .O(N__44582),
            .I(N__44579));
    LocalMux I__10274 (
            .O(N__44579),
            .I(N__44576));
    Span4Mux_h I__10273 (
            .O(N__44576),
            .I(N__44573));
    Odrv4 I__10272 (
            .O(N__44573),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__10271 (
            .O(N__44570),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    CascadeMux I__10270 (
            .O(N__44567),
            .I(N__44564));
    InMux I__10269 (
            .O(N__44564),
            .I(N__44561));
    LocalMux I__10268 (
            .O(N__44561),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__10267 (
            .O(N__44558),
            .I(N__44555));
    LocalMux I__10266 (
            .O(N__44555),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__10265 (
            .O(N__44552),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__10264 (
            .O(N__44549),
            .I(N__44546));
    LocalMux I__10263 (
            .O(N__44546),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__10262 (
            .O(N__44543),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    CascadeMux I__10261 (
            .O(N__44540),
            .I(N__44536));
    CascadeMux I__10260 (
            .O(N__44539),
            .I(N__44533));
    InMux I__10259 (
            .O(N__44536),
            .I(N__44530));
    InMux I__10258 (
            .O(N__44533),
            .I(N__44527));
    LocalMux I__10257 (
            .O(N__44530),
            .I(N__44524));
    LocalMux I__10256 (
            .O(N__44527),
            .I(N__44519));
    Span4Mux_h I__10255 (
            .O(N__44524),
            .I(N__44519));
    Odrv4 I__10254 (
            .O(N__44519),
            .I(\current_shift_inst.un4_control_input_0_31 ));
    InMux I__10253 (
            .O(N__44516),
            .I(N__44513));
    LocalMux I__10252 (
            .O(N__44513),
            .I(N__44510));
    Span4Mux_h I__10251 (
            .O(N__44510),
            .I(N__44507));
    Odrv4 I__10250 (
            .O(N__44507),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__10249 (
            .O(N__44504),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__10248 (
            .O(N__44501),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    CascadeMux I__10247 (
            .O(N__44498),
            .I(N__44495));
    InMux I__10246 (
            .O(N__44495),
            .I(N__44492));
    LocalMux I__10245 (
            .O(N__44492),
            .I(N__44489));
    Odrv4 I__10244 (
            .O(N__44489),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__10243 (
            .O(N__44486),
            .I(N__44483));
    LocalMux I__10242 (
            .O(N__44483),
            .I(N__44480));
    Odrv4 I__10241 (
            .O(N__44480),
            .I(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ));
    CascadeMux I__10240 (
            .O(N__44477),
            .I(N__44474));
    InMux I__10239 (
            .O(N__44474),
            .I(N__44471));
    LocalMux I__10238 (
            .O(N__44471),
            .I(N__44468));
    Span4Mux_h I__10237 (
            .O(N__44468),
            .I(N__44465));
    Span4Mux_h I__10236 (
            .O(N__44465),
            .I(N__44462));
    Odrv4 I__10235 (
            .O(N__44462),
            .I(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ));
    InMux I__10234 (
            .O(N__44459),
            .I(N__44456));
    LocalMux I__10233 (
            .O(N__44456),
            .I(N__44453));
    Span4Mux_h I__10232 (
            .O(N__44453),
            .I(N__44450));
    Odrv4 I__10231 (
            .O(N__44450),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__10230 (
            .O(N__44447),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__10229 (
            .O(N__44444),
            .I(N__44441));
    LocalMux I__10228 (
            .O(N__44441),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__10227 (
            .O(N__44438),
            .I(N__44435));
    LocalMux I__10226 (
            .O(N__44435),
            .I(N__44432));
    Odrv4 I__10225 (
            .O(N__44432),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__10224 (
            .O(N__44429),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    CascadeMux I__10223 (
            .O(N__44426),
            .I(N__44423));
    InMux I__10222 (
            .O(N__44423),
            .I(N__44420));
    LocalMux I__10221 (
            .O(N__44420),
            .I(N__44417));
    Span4Mux_h I__10220 (
            .O(N__44417),
            .I(N__44414));
    Odrv4 I__10219 (
            .O(N__44414),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__10218 (
            .O(N__44411),
            .I(N__44408));
    LocalMux I__10217 (
            .O(N__44408),
            .I(N__44405));
    Odrv12 I__10216 (
            .O(N__44405),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__10215 (
            .O(N__44402),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__10214 (
            .O(N__44399),
            .I(N__44396));
    LocalMux I__10213 (
            .O(N__44396),
            .I(N__44393));
    Span4Mux_h I__10212 (
            .O(N__44393),
            .I(N__44390));
    Odrv4 I__10211 (
            .O(N__44390),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__10210 (
            .O(N__44387),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__10209 (
            .O(N__44384),
            .I(N__44381));
    LocalMux I__10208 (
            .O(N__44381),
            .I(N__44378));
    Odrv4 I__10207 (
            .O(N__44378),
            .I(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ));
    CascadeMux I__10206 (
            .O(N__44375),
            .I(N__44372));
    InMux I__10205 (
            .O(N__44372),
            .I(N__44369));
    LocalMux I__10204 (
            .O(N__44369),
            .I(N__44366));
    Span4Mux_h I__10203 (
            .O(N__44366),
            .I(N__44363));
    Odrv4 I__10202 (
            .O(N__44363),
            .I(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ));
    InMux I__10201 (
            .O(N__44360),
            .I(N__44357));
    LocalMux I__10200 (
            .O(N__44357),
            .I(N__44354));
    Span4Mux_h I__10199 (
            .O(N__44354),
            .I(N__44351));
    Odrv4 I__10198 (
            .O(N__44351),
            .I(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ));
    CascadeMux I__10197 (
            .O(N__44348),
            .I(N__44345));
    InMux I__10196 (
            .O(N__44345),
            .I(N__44342));
    LocalMux I__10195 (
            .O(N__44342),
            .I(N__44339));
    Odrv12 I__10194 (
            .O(N__44339),
            .I(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ));
    CascadeMux I__10193 (
            .O(N__44336),
            .I(N__44333));
    InMux I__10192 (
            .O(N__44333),
            .I(N__44330));
    LocalMux I__10191 (
            .O(N__44330),
            .I(N__44327));
    Span4Mux_h I__10190 (
            .O(N__44327),
            .I(N__44324));
    Odrv4 I__10189 (
            .O(N__44324),
            .I(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ));
    CascadeMux I__10188 (
            .O(N__44321),
            .I(N__44318));
    InMux I__10187 (
            .O(N__44318),
            .I(N__44315));
    LocalMux I__10186 (
            .O(N__44315),
            .I(N__44312));
    Span4Mux_v I__10185 (
            .O(N__44312),
            .I(N__44309));
    Odrv4 I__10184 (
            .O(N__44309),
            .I(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ));
    InMux I__10183 (
            .O(N__44306),
            .I(N__44303));
    LocalMux I__10182 (
            .O(N__44303),
            .I(N__44300));
    Span4Mux_h I__10181 (
            .O(N__44300),
            .I(N__44297));
    Odrv4 I__10180 (
            .O(N__44297),
            .I(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ));
    CEMux I__10179 (
            .O(N__44294),
            .I(N__44286));
    CEMux I__10178 (
            .O(N__44293),
            .I(N__44283));
    CEMux I__10177 (
            .O(N__44292),
            .I(N__44280));
    CEMux I__10176 (
            .O(N__44291),
            .I(N__44277));
    CEMux I__10175 (
            .O(N__44290),
            .I(N__44274));
    CEMux I__10174 (
            .O(N__44289),
            .I(N__44253));
    LocalMux I__10173 (
            .O(N__44286),
            .I(N__44250));
    LocalMux I__10172 (
            .O(N__44283),
            .I(N__44247));
    LocalMux I__10171 (
            .O(N__44280),
            .I(N__44244));
    LocalMux I__10170 (
            .O(N__44277),
            .I(N__44238));
    LocalMux I__10169 (
            .O(N__44274),
            .I(N__44238));
    InMux I__10168 (
            .O(N__44273),
            .I(N__44231));
    InMux I__10167 (
            .O(N__44272),
            .I(N__44231));
    InMux I__10166 (
            .O(N__44271),
            .I(N__44231));
    InMux I__10165 (
            .O(N__44270),
            .I(N__44228));
    InMux I__10164 (
            .O(N__44269),
            .I(N__44223));
    InMux I__10163 (
            .O(N__44268),
            .I(N__44223));
    InMux I__10162 (
            .O(N__44267),
            .I(N__44214));
    InMux I__10161 (
            .O(N__44266),
            .I(N__44214));
    InMux I__10160 (
            .O(N__44265),
            .I(N__44214));
    InMux I__10159 (
            .O(N__44264),
            .I(N__44214));
    InMux I__10158 (
            .O(N__44263),
            .I(N__44205));
    InMux I__10157 (
            .O(N__44262),
            .I(N__44205));
    InMux I__10156 (
            .O(N__44261),
            .I(N__44205));
    InMux I__10155 (
            .O(N__44260),
            .I(N__44205));
    InMux I__10154 (
            .O(N__44259),
            .I(N__44196));
    InMux I__10153 (
            .O(N__44258),
            .I(N__44196));
    InMux I__10152 (
            .O(N__44257),
            .I(N__44196));
    InMux I__10151 (
            .O(N__44256),
            .I(N__44196));
    LocalMux I__10150 (
            .O(N__44253),
            .I(N__44193));
    Span4Mux_v I__10149 (
            .O(N__44250),
            .I(N__44188));
    Span4Mux_h I__10148 (
            .O(N__44247),
            .I(N__44188));
    Span4Mux_v I__10147 (
            .O(N__44244),
            .I(N__44185));
    InMux I__10146 (
            .O(N__44243),
            .I(N__44182));
    Span4Mux_v I__10145 (
            .O(N__44238),
            .I(N__44179));
    LocalMux I__10144 (
            .O(N__44231),
            .I(N__44176));
    LocalMux I__10143 (
            .O(N__44228),
            .I(N__44165));
    LocalMux I__10142 (
            .O(N__44223),
            .I(N__44165));
    LocalMux I__10141 (
            .O(N__44214),
            .I(N__44165));
    LocalMux I__10140 (
            .O(N__44205),
            .I(N__44165));
    LocalMux I__10139 (
            .O(N__44196),
            .I(N__44165));
    Span4Mux_v I__10138 (
            .O(N__44193),
            .I(N__44160));
    Span4Mux_v I__10137 (
            .O(N__44188),
            .I(N__44160));
    Span4Mux_h I__10136 (
            .O(N__44185),
            .I(N__44155));
    LocalMux I__10135 (
            .O(N__44182),
            .I(N__44155));
    Span4Mux_v I__10134 (
            .O(N__44179),
            .I(N__44148));
    Span4Mux_v I__10133 (
            .O(N__44176),
            .I(N__44148));
    Span4Mux_v I__10132 (
            .O(N__44165),
            .I(N__44148));
    Odrv4 I__10131 (
            .O(N__44160),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__10130 (
            .O(N__44155),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__10129 (
            .O(N__44148),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    InMux I__10128 (
            .O(N__44141),
            .I(N__44134));
    InMux I__10127 (
            .O(N__44140),
            .I(N__44134));
    InMux I__10126 (
            .O(N__44139),
            .I(N__44131));
    LocalMux I__10125 (
            .O(N__44134),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__10124 (
            .O(N__44131),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    CascadeMux I__10123 (
            .O(N__44126),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0_cascade_ ));
    CascadeMux I__10122 (
            .O(N__44123),
            .I(N__44118));
    InMux I__10121 (
            .O(N__44122),
            .I(N__44115));
    InMux I__10120 (
            .O(N__44121),
            .I(N__44112));
    InMux I__10119 (
            .O(N__44118),
            .I(N__44109));
    LocalMux I__10118 (
            .O(N__44115),
            .I(N__44106));
    LocalMux I__10117 (
            .O(N__44112),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__10116 (
            .O(N__44109),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__10115 (
            .O(N__44106),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__10114 (
            .O(N__44099),
            .I(N__44096));
    LocalMux I__10113 (
            .O(N__44096),
            .I(N__44092));
    CascadeMux I__10112 (
            .O(N__44095),
            .I(N__44089));
    Span4Mux_h I__10111 (
            .O(N__44092),
            .I(N__44086));
    InMux I__10110 (
            .O(N__44089),
            .I(N__44083));
    Odrv4 I__10109 (
            .O(N__44086),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    LocalMux I__10108 (
            .O(N__44083),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    InMux I__10107 (
            .O(N__44078),
            .I(N__44074));
    CascadeMux I__10106 (
            .O(N__44077),
            .I(N__44071));
    LocalMux I__10105 (
            .O(N__44074),
            .I(N__44068));
    InMux I__10104 (
            .O(N__44071),
            .I(N__44065));
    Span4Mux_v I__10103 (
            .O(N__44068),
            .I(N__44062));
    LocalMux I__10102 (
            .O(N__44065),
            .I(N__44059));
    Odrv4 I__10101 (
            .O(N__44062),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    Odrv12 I__10100 (
            .O(N__44059),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    CascadeMux I__10099 (
            .O(N__44054),
            .I(N__44050));
    InMux I__10098 (
            .O(N__44053),
            .I(N__44045));
    InMux I__10097 (
            .O(N__44050),
            .I(N__44045));
    LocalMux I__10096 (
            .O(N__44045),
            .I(N__44041));
    InMux I__10095 (
            .O(N__44044),
            .I(N__44037));
    Span4Mux_v I__10094 (
            .O(N__44041),
            .I(N__44034));
    InMux I__10093 (
            .O(N__44040),
            .I(N__44031));
    LocalMux I__10092 (
            .O(N__44037),
            .I(N__44028));
    Odrv4 I__10091 (
            .O(N__44034),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__10090 (
            .O(N__44031),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv12 I__10089 (
            .O(N__44028),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    CascadeMux I__10088 (
            .O(N__44021),
            .I(N__44018));
    InMux I__10087 (
            .O(N__44018),
            .I(N__44015));
    LocalMux I__10086 (
            .O(N__44015),
            .I(N__44012));
    Span4Mux_h I__10085 (
            .O(N__44012),
            .I(N__44009));
    Span4Mux_h I__10084 (
            .O(N__44009),
            .I(N__44006));
    Odrv4 I__10083 (
            .O(N__44006),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    CascadeMux I__10082 (
            .O(N__44003),
            .I(N__44000));
    InMux I__10081 (
            .O(N__44000),
            .I(N__43997));
    LocalMux I__10080 (
            .O(N__43997),
            .I(N__43994));
    Span4Mux_h I__10079 (
            .O(N__43994),
            .I(N__43991));
    Odrv4 I__10078 (
            .O(N__43991),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    InMux I__10077 (
            .O(N__43988),
            .I(N__43985));
    LocalMux I__10076 (
            .O(N__43985),
            .I(N__43982));
    Span4Mux_v I__10075 (
            .O(N__43982),
            .I(N__43979));
    Odrv4 I__10074 (
            .O(N__43979),
            .I(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ));
    CascadeMux I__10073 (
            .O(N__43976),
            .I(N__43973));
    InMux I__10072 (
            .O(N__43973),
            .I(N__43970));
    LocalMux I__10071 (
            .O(N__43970),
            .I(N__43967));
    Span4Mux_h I__10070 (
            .O(N__43967),
            .I(N__43964));
    Odrv4 I__10069 (
            .O(N__43964),
            .I(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ));
    InMux I__10068 (
            .O(N__43961),
            .I(N__43958));
    LocalMux I__10067 (
            .O(N__43958),
            .I(N__43955));
    Span4Mux_h I__10066 (
            .O(N__43955),
            .I(N__43952));
    Span4Mux_h I__10065 (
            .O(N__43952),
            .I(N__43949));
    Odrv4 I__10064 (
            .O(N__43949),
            .I(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ));
    CascadeMux I__10063 (
            .O(N__43946),
            .I(N__43943));
    InMux I__10062 (
            .O(N__43943),
            .I(N__43940));
    LocalMux I__10061 (
            .O(N__43940),
            .I(N__43937));
    Odrv12 I__10060 (
            .O(N__43937),
            .I(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ));
    InMux I__10059 (
            .O(N__43934),
            .I(N__43930));
    InMux I__10058 (
            .O(N__43933),
            .I(N__43927));
    LocalMux I__10057 (
            .O(N__43930),
            .I(N__43922));
    LocalMux I__10056 (
            .O(N__43927),
            .I(N__43919));
    InMux I__10055 (
            .O(N__43926),
            .I(N__43916));
    InMux I__10054 (
            .O(N__43925),
            .I(N__43913));
    Span12Mux_s7_h I__10053 (
            .O(N__43922),
            .I(N__43908));
    Span12Mux_s9_v I__10052 (
            .O(N__43919),
            .I(N__43908));
    LocalMux I__10051 (
            .O(N__43916),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__10050 (
            .O(N__43913),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv12 I__10049 (
            .O(N__43908),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__10048 (
            .O(N__43901),
            .I(N__43898));
    LocalMux I__10047 (
            .O(N__43898),
            .I(N__43892));
    InMux I__10046 (
            .O(N__43897),
            .I(N__43889));
    InMux I__10045 (
            .O(N__43896),
            .I(N__43884));
    InMux I__10044 (
            .O(N__43895),
            .I(N__43884));
    Span4Mux_h I__10043 (
            .O(N__43892),
            .I(N__43881));
    LocalMux I__10042 (
            .O(N__43889),
            .I(N__43878));
    LocalMux I__10041 (
            .O(N__43884),
            .I(N__43874));
    Span4Mux_v I__10040 (
            .O(N__43881),
            .I(N__43869));
    Span4Mux_h I__10039 (
            .O(N__43878),
            .I(N__43869));
    InMux I__10038 (
            .O(N__43877),
            .I(N__43866));
    Span4Mux_h I__10037 (
            .O(N__43874),
            .I(N__43863));
    Span4Mux_h I__10036 (
            .O(N__43869),
            .I(N__43860));
    LocalMux I__10035 (
            .O(N__43866),
            .I(N__43855));
    Span4Mux_h I__10034 (
            .O(N__43863),
            .I(N__43855));
    Odrv4 I__10033 (
            .O(N__43860),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__10032 (
            .O(N__43855),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    CascadeMux I__10031 (
            .O(N__43850),
            .I(N__43847));
    InMux I__10030 (
            .O(N__43847),
            .I(N__43842));
    InMux I__10029 (
            .O(N__43846),
            .I(N__43839));
    InMux I__10028 (
            .O(N__43845),
            .I(N__43836));
    LocalMux I__10027 (
            .O(N__43842),
            .I(N__43832));
    LocalMux I__10026 (
            .O(N__43839),
            .I(N__43829));
    LocalMux I__10025 (
            .O(N__43836),
            .I(N__43826));
    CascadeMux I__10024 (
            .O(N__43835),
            .I(N__43822));
    Span4Mux_v I__10023 (
            .O(N__43832),
            .I(N__43817));
    Span4Mux_v I__10022 (
            .O(N__43829),
            .I(N__43817));
    Span4Mux_h I__10021 (
            .O(N__43826),
            .I(N__43814));
    InMux I__10020 (
            .O(N__43825),
            .I(N__43811));
    InMux I__10019 (
            .O(N__43822),
            .I(N__43808));
    Span4Mux_h I__10018 (
            .O(N__43817),
            .I(N__43805));
    Span4Mux_h I__10017 (
            .O(N__43814),
            .I(N__43800));
    LocalMux I__10016 (
            .O(N__43811),
            .I(N__43800));
    LocalMux I__10015 (
            .O(N__43808),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__10014 (
            .O(N__43805),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__10013 (
            .O(N__43800),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    InMux I__10012 (
            .O(N__43793),
            .I(N__43789));
    InMux I__10011 (
            .O(N__43792),
            .I(N__43786));
    LocalMux I__10010 (
            .O(N__43789),
            .I(N__43783));
    LocalMux I__10009 (
            .O(N__43786),
            .I(N__43777));
    Span4Mux_h I__10008 (
            .O(N__43783),
            .I(N__43777));
    InMux I__10007 (
            .O(N__43782),
            .I(N__43774));
    Span4Mux_h I__10006 (
            .O(N__43777),
            .I(N__43769));
    LocalMux I__10005 (
            .O(N__43774),
            .I(N__43769));
    Span4Mux_v I__10004 (
            .O(N__43769),
            .I(N__43766));
    Odrv4 I__10003 (
            .O(N__43766),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO ));
    InMux I__10002 (
            .O(N__43763),
            .I(N__43759));
    InMux I__10001 (
            .O(N__43762),
            .I(N__43756));
    LocalMux I__10000 (
            .O(N__43759),
            .I(N__43753));
    LocalMux I__9999 (
            .O(N__43756),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    Odrv4 I__9998 (
            .O(N__43753),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    InMux I__9997 (
            .O(N__43748),
            .I(N__43745));
    LocalMux I__9996 (
            .O(N__43745),
            .I(N__43742));
    Span4Mux_h I__9995 (
            .O(N__43742),
            .I(N__43737));
    InMux I__9994 (
            .O(N__43741),
            .I(N__43734));
    InMux I__9993 (
            .O(N__43740),
            .I(N__43731));
    Span4Mux_h I__9992 (
            .O(N__43737),
            .I(N__43728));
    LocalMux I__9991 (
            .O(N__43734),
            .I(N__43725));
    LocalMux I__9990 (
            .O(N__43731),
            .I(N__43722));
    Span4Mux_v I__9989 (
            .O(N__43728),
            .I(N__43719));
    Span4Mux_v I__9988 (
            .O(N__43725),
            .I(N__43716));
    Span4Mux_v I__9987 (
            .O(N__43722),
            .I(N__43713));
    Sp12to4 I__9986 (
            .O(N__43719),
            .I(N__43710));
    Span4Mux_h I__9985 (
            .O(N__43716),
            .I(N__43707));
    Odrv4 I__9984 (
            .O(N__43713),
            .I(il_min_comp2_D2));
    Odrv12 I__9983 (
            .O(N__43710),
            .I(il_min_comp2_D2));
    Odrv4 I__9982 (
            .O(N__43707),
            .I(il_min_comp2_D2));
    InMux I__9981 (
            .O(N__43700),
            .I(N__43697));
    LocalMux I__9980 (
            .O(N__43697),
            .I(\phase_controller_inst2.start_timer_tr_0_sqmuxa ));
    InMux I__9979 (
            .O(N__43694),
            .I(N__43691));
    LocalMux I__9978 (
            .O(N__43691),
            .I(N__43688));
    Span4Mux_h I__9977 (
            .O(N__43688),
            .I(N__43685));
    Span4Mux_h I__9976 (
            .O(N__43685),
            .I(N__43682));
    Odrv4 I__9975 (
            .O(N__43682),
            .I(\phase_controller_inst2.time_passed_RNI9M3O ));
    CascadeMux I__9974 (
            .O(N__43679),
            .I(N__43674));
    CascadeMux I__9973 (
            .O(N__43678),
            .I(N__43671));
    InMux I__9972 (
            .O(N__43677),
            .I(N__43668));
    InMux I__9971 (
            .O(N__43674),
            .I(N__43665));
    InMux I__9970 (
            .O(N__43671),
            .I(N__43660));
    LocalMux I__9969 (
            .O(N__43668),
            .I(N__43657));
    LocalMux I__9968 (
            .O(N__43665),
            .I(N__43654));
    InMux I__9967 (
            .O(N__43664),
            .I(N__43651));
    InMux I__9966 (
            .O(N__43663),
            .I(N__43647));
    LocalMux I__9965 (
            .O(N__43660),
            .I(N__43644));
    Span4Mux_v I__9964 (
            .O(N__43657),
            .I(N__43641));
    Span4Mux_h I__9963 (
            .O(N__43654),
            .I(N__43636));
    LocalMux I__9962 (
            .O(N__43651),
            .I(N__43636));
    InMux I__9961 (
            .O(N__43650),
            .I(N__43633));
    LocalMux I__9960 (
            .O(N__43647),
            .I(N__43628));
    Span4Mux_h I__9959 (
            .O(N__43644),
            .I(N__43628));
    Span4Mux_v I__9958 (
            .O(N__43641),
            .I(N__43623));
    Span4Mux_h I__9957 (
            .O(N__43636),
            .I(N__43623));
    LocalMux I__9956 (
            .O(N__43633),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__9955 (
            .O(N__43628),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__9954 (
            .O(N__43623),
            .I(phase_controller_inst1_state_4));
    InMux I__9953 (
            .O(N__43616),
            .I(N__43613));
    LocalMux I__9952 (
            .O(N__43613),
            .I(N__43609));
    InMux I__9951 (
            .O(N__43612),
            .I(N__43605));
    Span4Mux_h I__9950 (
            .O(N__43609),
            .I(N__43602));
    InMux I__9949 (
            .O(N__43608),
            .I(N__43599));
    LocalMux I__9948 (
            .O(N__43605),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO ));
    Odrv4 I__9947 (
            .O(N__43602),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO ));
    LocalMux I__9946 (
            .O(N__43599),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO ));
    CascadeMux I__9945 (
            .O(N__43592),
            .I(N__43589));
    InMux I__9944 (
            .O(N__43589),
            .I(N__43586));
    LocalMux I__9943 (
            .O(N__43586),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIUMLHZ0Z1 ));
    CascadeMux I__9942 (
            .O(N__43583),
            .I(N__43580));
    InMux I__9941 (
            .O(N__43580),
            .I(N__43577));
    LocalMux I__9940 (
            .O(N__43577),
            .I(N__43574));
    Span4Mux_h I__9939 (
            .O(N__43574),
            .I(N__43569));
    InMux I__9938 (
            .O(N__43573),
            .I(N__43566));
    CascadeMux I__9937 (
            .O(N__43572),
            .I(N__43562));
    Span4Mux_h I__9936 (
            .O(N__43569),
            .I(N__43558));
    LocalMux I__9935 (
            .O(N__43566),
            .I(N__43555));
    InMux I__9934 (
            .O(N__43565),
            .I(N__43552));
    InMux I__9933 (
            .O(N__43562),
            .I(N__43547));
    InMux I__9932 (
            .O(N__43561),
            .I(N__43547));
    Odrv4 I__9931 (
            .O(N__43558),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__9930 (
            .O(N__43555),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__9929 (
            .O(N__43552),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__9928 (
            .O(N__43547),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    InMux I__9927 (
            .O(N__43538),
            .I(N__43532));
    InMux I__9926 (
            .O(N__43537),
            .I(N__43532));
    LocalMux I__9925 (
            .O(N__43532),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    InMux I__9924 (
            .O(N__43529),
            .I(N__43526));
    LocalMux I__9923 (
            .O(N__43526),
            .I(N__43520));
    InMux I__9922 (
            .O(N__43525),
            .I(N__43513));
    InMux I__9921 (
            .O(N__43524),
            .I(N__43513));
    InMux I__9920 (
            .O(N__43523),
            .I(N__43513));
    Odrv12 I__9919 (
            .O(N__43520),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__9918 (
            .O(N__43513),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    InMux I__9917 (
            .O(N__43508),
            .I(N__43505));
    LocalMux I__9916 (
            .O(N__43505),
            .I(N__43502));
    Span4Mux_h I__9915 (
            .O(N__43502),
            .I(N__43499));
    Span4Mux_h I__9914 (
            .O(N__43499),
            .I(N__43493));
    InMux I__9913 (
            .O(N__43498),
            .I(N__43488));
    InMux I__9912 (
            .O(N__43497),
            .I(N__43488));
    InMux I__9911 (
            .O(N__43496),
            .I(N__43485));
    Odrv4 I__9910 (
            .O(N__43493),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__9909 (
            .O(N__43488),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__9908 (
            .O(N__43485),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    CascadeMux I__9907 (
            .O(N__43478),
            .I(elapsed_time_ns_1_RNIVEIF91_0_25_cascade_));
    InMux I__9906 (
            .O(N__43475),
            .I(N__43471));
    InMux I__9905 (
            .O(N__43474),
            .I(N__43468));
    LocalMux I__9904 (
            .O(N__43471),
            .I(elapsed_time_ns_1_RNI0GIF91_0_26));
    LocalMux I__9903 (
            .O(N__43468),
            .I(elapsed_time_ns_1_RNI0GIF91_0_26));
    InMux I__9902 (
            .O(N__43463),
            .I(N__43460));
    LocalMux I__9901 (
            .O(N__43460),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15 ));
    InMux I__9900 (
            .O(N__43457),
            .I(N__43454));
    LocalMux I__9899 (
            .O(N__43454),
            .I(N__43450));
    InMux I__9898 (
            .O(N__43453),
            .I(N__43447));
    Span4Mux_h I__9897 (
            .O(N__43450),
            .I(N__43442));
    LocalMux I__9896 (
            .O(N__43447),
            .I(N__43442));
    Odrv4 I__9895 (
            .O(N__43442),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__9894 (
            .O(N__43439),
            .I(N__43433));
    InMux I__9893 (
            .O(N__43438),
            .I(N__43433));
    LocalMux I__9892 (
            .O(N__43433),
            .I(elapsed_time_ns_1_RNI2IIF91_0_28));
    InMux I__9891 (
            .O(N__43430),
            .I(N__43423));
    InMux I__9890 (
            .O(N__43429),
            .I(N__43420));
    InMux I__9889 (
            .O(N__43428),
            .I(N__43417));
    InMux I__9888 (
            .O(N__43427),
            .I(N__43414));
    InMux I__9887 (
            .O(N__43426),
            .I(N__43411));
    LocalMux I__9886 (
            .O(N__43423),
            .I(N__43408));
    LocalMux I__9885 (
            .O(N__43420),
            .I(N__43405));
    LocalMux I__9884 (
            .O(N__43417),
            .I(N__43398));
    LocalMux I__9883 (
            .O(N__43414),
            .I(N__43398));
    LocalMux I__9882 (
            .O(N__43411),
            .I(N__43398));
    Span4Mux_v I__9881 (
            .O(N__43408),
            .I(N__43393));
    Span4Mux_v I__9880 (
            .O(N__43405),
            .I(N__43393));
    Span4Mux_h I__9879 (
            .O(N__43398),
            .I(N__43390));
    Odrv4 I__9878 (
            .O(N__43393),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__9877 (
            .O(N__43390),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    CascadeMux I__9876 (
            .O(N__43385),
            .I(N__43382));
    InMux I__9875 (
            .O(N__43382),
            .I(N__43379));
    LocalMux I__9874 (
            .O(N__43379),
            .I(N__43374));
    InMux I__9873 (
            .O(N__43378),
            .I(N__43369));
    InMux I__9872 (
            .O(N__43377),
            .I(N__43369));
    Span4Mux_h I__9871 (
            .O(N__43374),
            .I(N__43366));
    LocalMux I__9870 (
            .O(N__43369),
            .I(\delay_measurement_inst.delay_tr_timer.N_378 ));
    Odrv4 I__9869 (
            .O(N__43366),
            .I(\delay_measurement_inst.delay_tr_timer.N_378 ));
    InMux I__9868 (
            .O(N__43361),
            .I(N__43358));
    LocalMux I__9867 (
            .O(N__43358),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0 ));
    InMux I__9866 (
            .O(N__43355),
            .I(N__43352));
    LocalMux I__9865 (
            .O(N__43352),
            .I(N__43348));
    InMux I__9864 (
            .O(N__43351),
            .I(N__43345));
    Odrv4 I__9863 (
            .O(N__43348),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    LocalMux I__9862 (
            .O(N__43345),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    CascadeMux I__9861 (
            .O(N__43340),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_ ));
    InMux I__9860 (
            .O(N__43337),
            .I(N__43333));
    InMux I__9859 (
            .O(N__43336),
            .I(N__43330));
    LocalMux I__9858 (
            .O(N__43333),
            .I(N__43324));
    LocalMux I__9857 (
            .O(N__43330),
            .I(N__43324));
    InMux I__9856 (
            .O(N__43329),
            .I(N__43320));
    Span4Mux_v I__9855 (
            .O(N__43324),
            .I(N__43317));
    InMux I__9854 (
            .O(N__43323),
            .I(N__43314));
    LocalMux I__9853 (
            .O(N__43320),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    Odrv4 I__9852 (
            .O(N__43317),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    LocalMux I__9851 (
            .O(N__43314),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    InMux I__9850 (
            .O(N__43307),
            .I(N__43303));
    CascadeMux I__9849 (
            .O(N__43306),
            .I(N__43300));
    LocalMux I__9848 (
            .O(N__43303),
            .I(N__43297));
    InMux I__9847 (
            .O(N__43300),
            .I(N__43294));
    Span4Mux_h I__9846 (
            .O(N__43297),
            .I(N__43289));
    LocalMux I__9845 (
            .O(N__43294),
            .I(N__43289));
    Odrv4 I__9844 (
            .O(N__43289),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    CascadeMux I__9843 (
            .O(N__43286),
            .I(N__43283));
    InMux I__9842 (
            .O(N__43283),
            .I(N__43280));
    LocalMux I__9841 (
            .O(N__43280),
            .I(N__43276));
    InMux I__9840 (
            .O(N__43279),
            .I(N__43273));
    Odrv4 I__9839 (
            .O(N__43276),
            .I(elapsed_time_ns_1_RNI1HIF91_0_27));
    LocalMux I__9838 (
            .O(N__43273),
            .I(elapsed_time_ns_1_RNI1HIF91_0_27));
    InMux I__9837 (
            .O(N__43268),
            .I(N__43264));
    CascadeMux I__9836 (
            .O(N__43267),
            .I(N__43261));
    LocalMux I__9835 (
            .O(N__43264),
            .I(N__43258));
    InMux I__9834 (
            .O(N__43261),
            .I(N__43255));
    Span4Mux_v I__9833 (
            .O(N__43258),
            .I(N__43252));
    LocalMux I__9832 (
            .O(N__43255),
            .I(N__43249));
    Odrv4 I__9831 (
            .O(N__43252),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    Odrv4 I__9830 (
            .O(N__43249),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    CascadeMux I__9829 (
            .O(N__43244),
            .I(N__43241));
    InMux I__9828 (
            .O(N__43241),
            .I(N__43237));
    InMux I__9827 (
            .O(N__43240),
            .I(N__43234));
    LocalMux I__9826 (
            .O(N__43237),
            .I(elapsed_time_ns_1_RNISBIF91_0_22));
    LocalMux I__9825 (
            .O(N__43234),
            .I(elapsed_time_ns_1_RNISBIF91_0_22));
    InMux I__9824 (
            .O(N__43229),
            .I(N__43225));
    InMux I__9823 (
            .O(N__43228),
            .I(N__43222));
    LocalMux I__9822 (
            .O(N__43225),
            .I(N__43219));
    LocalMux I__9821 (
            .O(N__43222),
            .I(N__43216));
    Span4Mux_v I__9820 (
            .O(N__43219),
            .I(N__43213));
    Span4Mux_h I__9819 (
            .O(N__43216),
            .I(N__43210));
    Odrv4 I__9818 (
            .O(N__43213),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    Odrv4 I__9817 (
            .O(N__43210),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__9816 (
            .O(N__43205),
            .I(N__43201));
    InMux I__9815 (
            .O(N__43204),
            .I(N__43198));
    LocalMux I__9814 (
            .O(N__43201),
            .I(elapsed_time_ns_1_RNIQ9IF91_0_20));
    LocalMux I__9813 (
            .O(N__43198),
            .I(elapsed_time_ns_1_RNIQ9IF91_0_20));
    InMux I__9812 (
            .O(N__43193),
            .I(N__43190));
    LocalMux I__9811 (
            .O(N__43190),
            .I(N__43186));
    InMux I__9810 (
            .O(N__43189),
            .I(N__43183));
    Span4Mux_v I__9809 (
            .O(N__43186),
            .I(N__43180));
    LocalMux I__9808 (
            .O(N__43183),
            .I(N__43177));
    Odrv4 I__9807 (
            .O(N__43180),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    Odrv4 I__9806 (
            .O(N__43177),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    CascadeMux I__9805 (
            .O(N__43172),
            .I(N__43164));
    CascadeMux I__9804 (
            .O(N__43171),
            .I(N__43161));
    CascadeMux I__9803 (
            .O(N__43170),
            .I(N__43158));
    CascadeMux I__9802 (
            .O(N__43169),
            .I(N__43153));
    InMux I__9801 (
            .O(N__43168),
            .I(N__43149));
    InMux I__9800 (
            .O(N__43167),
            .I(N__43142));
    InMux I__9799 (
            .O(N__43164),
            .I(N__43134));
    InMux I__9798 (
            .O(N__43161),
            .I(N__43127));
    InMux I__9797 (
            .O(N__43158),
            .I(N__43127));
    InMux I__9796 (
            .O(N__43157),
            .I(N__43127));
    InMux I__9795 (
            .O(N__43156),
            .I(N__43122));
    InMux I__9794 (
            .O(N__43153),
            .I(N__43122));
    InMux I__9793 (
            .O(N__43152),
            .I(N__43118));
    LocalMux I__9792 (
            .O(N__43149),
            .I(N__43115));
    InMux I__9791 (
            .O(N__43148),
            .I(N__43108));
    InMux I__9790 (
            .O(N__43147),
            .I(N__43108));
    InMux I__9789 (
            .O(N__43146),
            .I(N__43108));
    CascadeMux I__9788 (
            .O(N__43145),
            .I(N__43104));
    LocalMux I__9787 (
            .O(N__43142),
            .I(N__43096));
    InMux I__9786 (
            .O(N__43141),
            .I(N__43093));
    InMux I__9785 (
            .O(N__43140),
            .I(N__43090));
    InMux I__9784 (
            .O(N__43139),
            .I(N__43085));
    InMux I__9783 (
            .O(N__43138),
            .I(N__43085));
    InMux I__9782 (
            .O(N__43137),
            .I(N__43082));
    LocalMux I__9781 (
            .O(N__43134),
            .I(N__43079));
    LocalMux I__9780 (
            .O(N__43127),
            .I(N__43074));
    LocalMux I__9779 (
            .O(N__43122),
            .I(N__43074));
    CascadeMux I__9778 (
            .O(N__43121),
            .I(N__43066));
    LocalMux I__9777 (
            .O(N__43118),
            .I(N__43059));
    Span4Mux_v I__9776 (
            .O(N__43115),
            .I(N__43059));
    LocalMux I__9775 (
            .O(N__43108),
            .I(N__43059));
    InMux I__9774 (
            .O(N__43107),
            .I(N__43052));
    InMux I__9773 (
            .O(N__43104),
            .I(N__43052));
    InMux I__9772 (
            .O(N__43103),
            .I(N__43052));
    InMux I__9771 (
            .O(N__43102),
            .I(N__43049));
    InMux I__9770 (
            .O(N__43101),
            .I(N__43042));
    InMux I__9769 (
            .O(N__43100),
            .I(N__43042));
    InMux I__9768 (
            .O(N__43099),
            .I(N__43042));
    Span4Mux_h I__9767 (
            .O(N__43096),
            .I(N__43031));
    LocalMux I__9766 (
            .O(N__43093),
            .I(N__43031));
    LocalMux I__9765 (
            .O(N__43090),
            .I(N__43031));
    LocalMux I__9764 (
            .O(N__43085),
            .I(N__43031));
    LocalMux I__9763 (
            .O(N__43082),
            .I(N__43031));
    Span4Mux_h I__9762 (
            .O(N__43079),
            .I(N__43026));
    Span4Mux_v I__9761 (
            .O(N__43074),
            .I(N__43026));
    InMux I__9760 (
            .O(N__43073),
            .I(N__43013));
    InMux I__9759 (
            .O(N__43072),
            .I(N__43013));
    InMux I__9758 (
            .O(N__43071),
            .I(N__43013));
    InMux I__9757 (
            .O(N__43070),
            .I(N__43013));
    InMux I__9756 (
            .O(N__43069),
            .I(N__43013));
    InMux I__9755 (
            .O(N__43066),
            .I(N__43013));
    Span4Mux_h I__9754 (
            .O(N__43059),
            .I(N__43008));
    LocalMux I__9753 (
            .O(N__43052),
            .I(N__43008));
    LocalMux I__9752 (
            .O(N__43049),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__9751 (
            .O(N__43042),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__9750 (
            .O(N__43031),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__9749 (
            .O(N__43026),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__9748 (
            .O(N__43013),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__9747 (
            .O(N__43008),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    CascadeMux I__9746 (
            .O(N__42995),
            .I(N__42987));
    CascadeMux I__9745 (
            .O(N__42994),
            .I(N__42984));
    InMux I__9744 (
            .O(N__42993),
            .I(N__42979));
    CascadeMux I__9743 (
            .O(N__42992),
            .I(N__42976));
    CascadeMux I__9742 (
            .O(N__42991),
            .I(N__42972));
    InMux I__9741 (
            .O(N__42990),
            .I(N__42968));
    InMux I__9740 (
            .O(N__42987),
            .I(N__42963));
    InMux I__9739 (
            .O(N__42984),
            .I(N__42963));
    CascadeMux I__9738 (
            .O(N__42983),
            .I(N__42959));
    CascadeMux I__9737 (
            .O(N__42982),
            .I(N__42953));
    LocalMux I__9736 (
            .O(N__42979),
            .I(N__42947));
    InMux I__9735 (
            .O(N__42976),
            .I(N__42944));
    CascadeMux I__9734 (
            .O(N__42975),
            .I(N__42937));
    InMux I__9733 (
            .O(N__42972),
            .I(N__42934));
    InMux I__9732 (
            .O(N__42971),
            .I(N__42931));
    LocalMux I__9731 (
            .O(N__42968),
            .I(N__42926));
    LocalMux I__9730 (
            .O(N__42963),
            .I(N__42926));
    InMux I__9729 (
            .O(N__42962),
            .I(N__42923));
    InMux I__9728 (
            .O(N__42959),
            .I(N__42916));
    InMux I__9727 (
            .O(N__42958),
            .I(N__42916));
    InMux I__9726 (
            .O(N__42957),
            .I(N__42916));
    InMux I__9725 (
            .O(N__42956),
            .I(N__42913));
    InMux I__9724 (
            .O(N__42953),
            .I(N__42908));
    InMux I__9723 (
            .O(N__42952),
            .I(N__42908));
    InMux I__9722 (
            .O(N__42951),
            .I(N__42903));
    InMux I__9721 (
            .O(N__42950),
            .I(N__42903));
    Span4Mux_h I__9720 (
            .O(N__42947),
            .I(N__42898));
    LocalMux I__9719 (
            .O(N__42944),
            .I(N__42898));
    InMux I__9718 (
            .O(N__42943),
            .I(N__42889));
    InMux I__9717 (
            .O(N__42942),
            .I(N__42889));
    InMux I__9716 (
            .O(N__42941),
            .I(N__42889));
    InMux I__9715 (
            .O(N__42940),
            .I(N__42889));
    InMux I__9714 (
            .O(N__42937),
            .I(N__42886));
    LocalMux I__9713 (
            .O(N__42934),
            .I(N__42881));
    LocalMux I__9712 (
            .O(N__42931),
            .I(N__42881));
    Span4Mux_v I__9711 (
            .O(N__42926),
            .I(N__42878));
    LocalMux I__9710 (
            .O(N__42923),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__9709 (
            .O(N__42916),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__9708 (
            .O(N__42913),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__9707 (
            .O(N__42908),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__9706 (
            .O(N__42903),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    Odrv4 I__9705 (
            .O(N__42898),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__9704 (
            .O(N__42889),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__9703 (
            .O(N__42886),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    Odrv12 I__9702 (
            .O(N__42881),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    Odrv4 I__9701 (
            .O(N__42878),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    CascadeMux I__9700 (
            .O(N__42857),
            .I(N__42854));
    InMux I__9699 (
            .O(N__42854),
            .I(N__42850));
    InMux I__9698 (
            .O(N__42853),
            .I(N__42847));
    LocalMux I__9697 (
            .O(N__42850),
            .I(elapsed_time_ns_1_RNIRBJF91_0_30));
    LocalMux I__9696 (
            .O(N__42847),
            .I(elapsed_time_ns_1_RNIRBJF91_0_30));
    CascadeMux I__9695 (
            .O(N__42842),
            .I(N__42839));
    InMux I__9694 (
            .O(N__42839),
            .I(N__42835));
    InMux I__9693 (
            .O(N__42838),
            .I(N__42832));
    LocalMux I__9692 (
            .O(N__42835),
            .I(N__42827));
    LocalMux I__9691 (
            .O(N__42832),
            .I(N__42827));
    Odrv4 I__9690 (
            .O(N__42827),
            .I(\delay_measurement_inst.delay_tr_timer.N_367 ));
    InMux I__9689 (
            .O(N__42824),
            .I(N__42820));
    InMux I__9688 (
            .O(N__42823),
            .I(N__42817));
    LocalMux I__9687 (
            .O(N__42820),
            .I(N__42814));
    LocalMux I__9686 (
            .O(N__42817),
            .I(N__42811));
    Span4Mux_v I__9685 (
            .O(N__42814),
            .I(N__42807));
    Span4Mux_h I__9684 (
            .O(N__42811),
            .I(N__42804));
    InMux I__9683 (
            .O(N__42810),
            .I(N__42801));
    Odrv4 I__9682 (
            .O(N__42807),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ));
    Odrv4 I__9681 (
            .O(N__42804),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ));
    LocalMux I__9680 (
            .O(N__42801),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ));
    CascadeMux I__9679 (
            .O(N__42794),
            .I(N__42791));
    InMux I__9678 (
            .O(N__42791),
            .I(N__42786));
    CascadeMux I__9677 (
            .O(N__42790),
            .I(N__42782));
    CascadeMux I__9676 (
            .O(N__42789),
            .I(N__42779));
    LocalMux I__9675 (
            .O(N__42786),
            .I(N__42776));
    InMux I__9674 (
            .O(N__42785),
            .I(N__42771));
    InMux I__9673 (
            .O(N__42782),
            .I(N__42771));
    InMux I__9672 (
            .O(N__42779),
            .I(N__42768));
    Span4Mux_v I__9671 (
            .O(N__42776),
            .I(N__42765));
    LocalMux I__9670 (
            .O(N__42771),
            .I(N__42762));
    LocalMux I__9669 (
            .O(N__42768),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    Odrv4 I__9668 (
            .O(N__42765),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    Odrv4 I__9667 (
            .O(N__42762),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    InMux I__9666 (
            .O(N__42755),
            .I(N__42752));
    LocalMux I__9665 (
            .O(N__42752),
            .I(\delay_measurement_inst.delay_tr_timer.N_349 ));
    CascadeMux I__9664 (
            .O(N__42749),
            .I(\delay_measurement_inst.delay_tr_timer.N_363_cascade_ ));
    CascadeMux I__9663 (
            .O(N__42746),
            .I(N__42742));
    CascadeMux I__9662 (
            .O(N__42745),
            .I(N__42738));
    InMux I__9661 (
            .O(N__42742),
            .I(N__42730));
    InMux I__9660 (
            .O(N__42741),
            .I(N__42727));
    InMux I__9659 (
            .O(N__42738),
            .I(N__42724));
    InMux I__9658 (
            .O(N__42737),
            .I(N__42721));
    InMux I__9657 (
            .O(N__42736),
            .I(N__42716));
    InMux I__9656 (
            .O(N__42735),
            .I(N__42716));
    InMux I__9655 (
            .O(N__42734),
            .I(N__42713));
    InMux I__9654 (
            .O(N__42733),
            .I(N__42710));
    LocalMux I__9653 (
            .O(N__42730),
            .I(N__42699));
    LocalMux I__9652 (
            .O(N__42727),
            .I(N__42699));
    LocalMux I__9651 (
            .O(N__42724),
            .I(N__42699));
    LocalMux I__9650 (
            .O(N__42721),
            .I(N__42699));
    LocalMux I__9649 (
            .O(N__42716),
            .I(N__42699));
    LocalMux I__9648 (
            .O(N__42713),
            .I(N__42696));
    LocalMux I__9647 (
            .O(N__42710),
            .I(N__42690));
    Span4Mux_v I__9646 (
            .O(N__42699),
            .I(N__42690));
    Span4Mux_v I__9645 (
            .O(N__42696),
            .I(N__42687));
    InMux I__9644 (
            .O(N__42695),
            .I(N__42684));
    Span4Mux_h I__9643 (
            .O(N__42690),
            .I(N__42681));
    Odrv4 I__9642 (
            .O(N__42687),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9 ));
    LocalMux I__9641 (
            .O(N__42684),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9 ));
    Odrv4 I__9640 (
            .O(N__42681),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9 ));
    InMux I__9639 (
            .O(N__42674),
            .I(N__42671));
    LocalMux I__9638 (
            .O(N__42671),
            .I(N__42667));
    InMux I__9637 (
            .O(N__42670),
            .I(N__42664));
    Odrv4 I__9636 (
            .O(N__42667),
            .I(\delay_measurement_inst.delay_tr_timer.N_380 ));
    LocalMux I__9635 (
            .O(N__42664),
            .I(\delay_measurement_inst.delay_tr_timer.N_380 ));
    CascadeMux I__9634 (
            .O(N__42659),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9_cascade_ ));
    InMux I__9633 (
            .O(N__42656),
            .I(N__42653));
    LocalMux I__9632 (
            .O(N__42653),
            .I(N__42650));
    Odrv4 I__9631 (
            .O(N__42650),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6 ));
    CascadeMux I__9630 (
            .O(N__42647),
            .I(N__42644));
    InMux I__9629 (
            .O(N__42644),
            .I(N__42640));
    InMux I__9628 (
            .O(N__42643),
            .I(N__42637));
    LocalMux I__9627 (
            .O(N__42640),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8 ));
    LocalMux I__9626 (
            .O(N__42637),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8 ));
    InMux I__9625 (
            .O(N__42632),
            .I(N__42627));
    InMux I__9624 (
            .O(N__42631),
            .I(N__42622));
    InMux I__9623 (
            .O(N__42630),
            .I(N__42622));
    LocalMux I__9622 (
            .O(N__42627),
            .I(N__42617));
    LocalMux I__9621 (
            .O(N__42622),
            .I(N__42617));
    Odrv4 I__9620 (
            .O(N__42617),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7 ));
    InMux I__9619 (
            .O(N__42614),
            .I(N__42609));
    InMux I__9618 (
            .O(N__42613),
            .I(N__42604));
    InMux I__9617 (
            .O(N__42612),
            .I(N__42604));
    LocalMux I__9616 (
            .O(N__42609),
            .I(\delay_measurement_inst.delay_tr_timer.N_365 ));
    LocalMux I__9615 (
            .O(N__42604),
            .I(\delay_measurement_inst.delay_tr_timer.N_365 ));
    CascadeMux I__9614 (
            .O(N__42599),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8_cascade_ ));
    CascadeMux I__9613 (
            .O(N__42596),
            .I(N__42592));
    InMux I__9612 (
            .O(N__42595),
            .I(N__42589));
    InMux I__9611 (
            .O(N__42592),
            .I(N__42586));
    LocalMux I__9610 (
            .O(N__42589),
            .I(\delay_measurement_inst.delay_tr_timer.N_345 ));
    LocalMux I__9609 (
            .O(N__42586),
            .I(\delay_measurement_inst.delay_tr_timer.N_345 ));
    InMux I__9608 (
            .O(N__42581),
            .I(N__42575));
    InMux I__9607 (
            .O(N__42580),
            .I(N__42575));
    LocalMux I__9606 (
            .O(N__42575),
            .I(\delay_measurement_inst.delay_tr_timer.N_359_1 ));
    CascadeMux I__9605 (
            .O(N__42572),
            .I(N__42568));
    CascadeMux I__9604 (
            .O(N__42571),
            .I(N__42565));
    InMux I__9603 (
            .O(N__42568),
            .I(N__42560));
    InMux I__9602 (
            .O(N__42565),
            .I(N__42560));
    LocalMux I__9601 (
            .O(N__42560),
            .I(N__42557));
    Span4Mux_h I__9600 (
            .O(N__42557),
            .I(N__42554));
    Odrv4 I__9599 (
            .O(N__42554),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__9598 (
            .O(N__42551),
            .I(N__42548));
    LocalMux I__9597 (
            .O(N__42548),
            .I(N__42545));
    Span4Mux_v I__9596 (
            .O(N__42545),
            .I(N__42541));
    InMux I__9595 (
            .O(N__42544),
            .I(N__42538));
    Odrv4 I__9594 (
            .O(N__42541),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    LocalMux I__9593 (
            .O(N__42538),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    CascadeMux I__9592 (
            .O(N__42533),
            .I(N__42530));
    InMux I__9591 (
            .O(N__42530),
            .I(N__42526));
    InMux I__9590 (
            .O(N__42529),
            .I(N__42523));
    LocalMux I__9589 (
            .O(N__42526),
            .I(elapsed_time_ns_1_RNIUDIF91_0_24));
    LocalMux I__9588 (
            .O(N__42523),
            .I(elapsed_time_ns_1_RNIUDIF91_0_24));
    InMux I__9587 (
            .O(N__42518),
            .I(N__42514));
    InMux I__9586 (
            .O(N__42517),
            .I(N__42511));
    LocalMux I__9585 (
            .O(N__42514),
            .I(N__42508));
    LocalMux I__9584 (
            .O(N__42511),
            .I(N__42505));
    Span4Mux_h I__9583 (
            .O(N__42508),
            .I(N__42502));
    Span4Mux_h I__9582 (
            .O(N__42505),
            .I(N__42499));
    Odrv4 I__9581 (
            .O(N__42502),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    Odrv4 I__9580 (
            .O(N__42499),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__9579 (
            .O(N__42494),
            .I(N__42491));
    LocalMux I__9578 (
            .O(N__42491),
            .I(elapsed_time_ns_1_RNIVEIF91_0_25));
    InMux I__9577 (
            .O(N__42488),
            .I(N__42483));
    InMux I__9576 (
            .O(N__42487),
            .I(N__42480));
    InMux I__9575 (
            .O(N__42486),
            .I(N__42477));
    LocalMux I__9574 (
            .O(N__42483),
            .I(N__42474));
    LocalMux I__9573 (
            .O(N__42480),
            .I(N__42471));
    LocalMux I__9572 (
            .O(N__42477),
            .I(N__42468));
    Span4Mux_h I__9571 (
            .O(N__42474),
            .I(N__42464));
    Sp12to4 I__9570 (
            .O(N__42471),
            .I(N__42461));
    Span4Mux_h I__9569 (
            .O(N__42468),
            .I(N__42458));
    InMux I__9568 (
            .O(N__42467),
            .I(N__42455));
    Odrv4 I__9567 (
            .O(N__42464),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv12 I__9566 (
            .O(N__42461),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__9565 (
            .O(N__42458),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__9564 (
            .O(N__42455),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    CascadeMux I__9563 (
            .O(N__42446),
            .I(N__42442));
    CascadeMux I__9562 (
            .O(N__42445),
            .I(N__42438));
    InMux I__9561 (
            .O(N__42442),
            .I(N__42435));
    InMux I__9560 (
            .O(N__42441),
            .I(N__42432));
    InMux I__9559 (
            .O(N__42438),
            .I(N__42429));
    LocalMux I__9558 (
            .O(N__42435),
            .I(N__42426));
    LocalMux I__9557 (
            .O(N__42432),
            .I(N__42423));
    LocalMux I__9556 (
            .O(N__42429),
            .I(N__42420));
    Span4Mux_h I__9555 (
            .O(N__42426),
            .I(N__42415));
    Span4Mux_v I__9554 (
            .O(N__42423),
            .I(N__42415));
    Odrv4 I__9553 (
            .O(N__42420),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv4 I__9552 (
            .O(N__42415),
            .I(\current_shift_inst.un4_control_input1_13 ));
    CascadeMux I__9551 (
            .O(N__42410),
            .I(N__42407));
    InMux I__9550 (
            .O(N__42407),
            .I(N__42404));
    LocalMux I__9549 (
            .O(N__42404),
            .I(N__42401));
    Span4Mux_v I__9548 (
            .O(N__42401),
            .I(N__42398));
    Odrv4 I__9547 (
            .O(N__42398),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    InMux I__9546 (
            .O(N__42395),
            .I(N__42391));
    InMux I__9545 (
            .O(N__42394),
            .I(N__42388));
    LocalMux I__9544 (
            .O(N__42391),
            .I(N__42383));
    LocalMux I__9543 (
            .O(N__42388),
            .I(N__42380));
    InMux I__9542 (
            .O(N__42387),
            .I(N__42377));
    InMux I__9541 (
            .O(N__42386),
            .I(N__42374));
    Span4Mux_v I__9540 (
            .O(N__42383),
            .I(N__42371));
    Span4Mux_v I__9539 (
            .O(N__42380),
            .I(N__42368));
    LocalMux I__9538 (
            .O(N__42377),
            .I(N__42365));
    LocalMux I__9537 (
            .O(N__42374),
            .I(N__42362));
    Odrv4 I__9536 (
            .O(N__42371),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__9535 (
            .O(N__42368),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__9534 (
            .O(N__42365),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__9533 (
            .O(N__42362),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__9532 (
            .O(N__42353),
            .I(N__42350));
    LocalMux I__9531 (
            .O(N__42350),
            .I(N__42347));
    Span4Mux_h I__9530 (
            .O(N__42347),
            .I(N__42344));
    Odrv4 I__9529 (
            .O(N__42344),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    CascadeMux I__9528 (
            .O(N__42341),
            .I(N__42337));
    CascadeMux I__9527 (
            .O(N__42340),
            .I(N__42334));
    InMux I__9526 (
            .O(N__42337),
            .I(N__42331));
    InMux I__9525 (
            .O(N__42334),
            .I(N__42327));
    LocalMux I__9524 (
            .O(N__42331),
            .I(N__42324));
    InMux I__9523 (
            .O(N__42330),
            .I(N__42321));
    LocalMux I__9522 (
            .O(N__42327),
            .I(N__42318));
    Span4Mux_v I__9521 (
            .O(N__42324),
            .I(N__42315));
    LocalMux I__9520 (
            .O(N__42321),
            .I(N__42312));
    Span4Mux_v I__9519 (
            .O(N__42318),
            .I(N__42308));
    Span4Mux_v I__9518 (
            .O(N__42315),
            .I(N__42303));
    Span4Mux_h I__9517 (
            .O(N__42312),
            .I(N__42303));
    InMux I__9516 (
            .O(N__42311),
            .I(N__42300));
    Odrv4 I__9515 (
            .O(N__42308),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__9514 (
            .O(N__42303),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    LocalMux I__9513 (
            .O(N__42300),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__9512 (
            .O(N__42293),
            .I(N__42288));
    InMux I__9511 (
            .O(N__42292),
            .I(N__42285));
    InMux I__9510 (
            .O(N__42291),
            .I(N__42282));
    LocalMux I__9509 (
            .O(N__42288),
            .I(N__42279));
    LocalMux I__9508 (
            .O(N__42285),
            .I(N__42276));
    LocalMux I__9507 (
            .O(N__42282),
            .I(N__42271));
    Span4Mux_v I__9506 (
            .O(N__42279),
            .I(N__42271));
    Odrv4 I__9505 (
            .O(N__42276),
            .I(\current_shift_inst.un4_control_input1_23 ));
    Odrv4 I__9504 (
            .O(N__42271),
            .I(\current_shift_inst.un4_control_input1_23 ));
    CascadeMux I__9503 (
            .O(N__42266),
            .I(N__42263));
    InMux I__9502 (
            .O(N__42263),
            .I(N__42260));
    LocalMux I__9501 (
            .O(N__42260),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__9500 (
            .O(N__42257),
            .I(N__42242));
    InMux I__9499 (
            .O(N__42256),
            .I(N__42235));
    InMux I__9498 (
            .O(N__42255),
            .I(N__42232));
    InMux I__9497 (
            .O(N__42254),
            .I(N__42221));
    InMux I__9496 (
            .O(N__42253),
            .I(N__42221));
    InMux I__9495 (
            .O(N__42252),
            .I(N__42221));
    InMux I__9494 (
            .O(N__42251),
            .I(N__42221));
    InMux I__9493 (
            .O(N__42250),
            .I(N__42221));
    InMux I__9492 (
            .O(N__42249),
            .I(N__42205));
    InMux I__9491 (
            .O(N__42248),
            .I(N__42205));
    InMux I__9490 (
            .O(N__42247),
            .I(N__42205));
    InMux I__9489 (
            .O(N__42246),
            .I(N__42205));
    InMux I__9488 (
            .O(N__42245),
            .I(N__42205));
    LocalMux I__9487 (
            .O(N__42242),
            .I(N__42202));
    InMux I__9486 (
            .O(N__42241),
            .I(N__42193));
    InMux I__9485 (
            .O(N__42240),
            .I(N__42193));
    InMux I__9484 (
            .O(N__42239),
            .I(N__42193));
    InMux I__9483 (
            .O(N__42238),
            .I(N__42193));
    LocalMux I__9482 (
            .O(N__42235),
            .I(N__42185));
    LocalMux I__9481 (
            .O(N__42232),
            .I(N__42185));
    LocalMux I__9480 (
            .O(N__42221),
            .I(N__42182));
    InMux I__9479 (
            .O(N__42220),
            .I(N__42179));
    InMux I__9478 (
            .O(N__42219),
            .I(N__42174));
    InMux I__9477 (
            .O(N__42218),
            .I(N__42174));
    InMux I__9476 (
            .O(N__42217),
            .I(N__42169));
    InMux I__9475 (
            .O(N__42216),
            .I(N__42169));
    LocalMux I__9474 (
            .O(N__42205),
            .I(N__42162));
    Span4Mux_v I__9473 (
            .O(N__42202),
            .I(N__42162));
    LocalMux I__9472 (
            .O(N__42193),
            .I(N__42162));
    InMux I__9471 (
            .O(N__42192),
            .I(N__42159));
    InMux I__9470 (
            .O(N__42191),
            .I(N__42156));
    InMux I__9469 (
            .O(N__42190),
            .I(N__42153));
    Span4Mux_v I__9468 (
            .O(N__42185),
            .I(N__42148));
    Span4Mux_h I__9467 (
            .O(N__42182),
            .I(N__42148));
    LocalMux I__9466 (
            .O(N__42179),
            .I(N__42141));
    LocalMux I__9465 (
            .O(N__42174),
            .I(N__42141));
    LocalMux I__9464 (
            .O(N__42169),
            .I(N__42141));
    Span4Mux_h I__9463 (
            .O(N__42162),
            .I(N__42138));
    LocalMux I__9462 (
            .O(N__42159),
            .I(N__42133));
    LocalMux I__9461 (
            .O(N__42156),
            .I(N__42133));
    LocalMux I__9460 (
            .O(N__42153),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__9459 (
            .O(N__42148),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__9458 (
            .O(N__42141),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__9457 (
            .O(N__42138),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv12 I__9456 (
            .O(N__42133),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    CascadeMux I__9455 (
            .O(N__42122),
            .I(N__42118));
    InMux I__9454 (
            .O(N__42121),
            .I(N__42115));
    InMux I__9453 (
            .O(N__42118),
            .I(N__42112));
    LocalMux I__9452 (
            .O(N__42115),
            .I(N__42108));
    LocalMux I__9451 (
            .O(N__42112),
            .I(N__42105));
    InMux I__9450 (
            .O(N__42111),
            .I(N__42102));
    Span4Mux_v I__9449 (
            .O(N__42108),
            .I(N__42096));
    Span4Mux_h I__9448 (
            .O(N__42105),
            .I(N__42096));
    LocalMux I__9447 (
            .O(N__42102),
            .I(N__42093));
    InMux I__9446 (
            .O(N__42101),
            .I(N__42090));
    Odrv4 I__9445 (
            .O(N__42096),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv12 I__9444 (
            .O(N__42093),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    LocalMux I__9443 (
            .O(N__42090),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__9442 (
            .O(N__42083),
            .I(N__42078));
    InMux I__9441 (
            .O(N__42082),
            .I(N__42075));
    CascadeMux I__9440 (
            .O(N__42081),
            .I(N__42072));
    LocalMux I__9439 (
            .O(N__42078),
            .I(N__42067));
    LocalMux I__9438 (
            .O(N__42075),
            .I(N__42067));
    InMux I__9437 (
            .O(N__42072),
            .I(N__42064));
    Span4Mux_v I__9436 (
            .O(N__42067),
            .I(N__42061));
    LocalMux I__9435 (
            .O(N__42064),
            .I(\current_shift_inst.un4_control_input1_9 ));
    Odrv4 I__9434 (
            .O(N__42061),
            .I(\current_shift_inst.un4_control_input1_9 ));
    CascadeMux I__9433 (
            .O(N__42056),
            .I(N__42053));
    InMux I__9432 (
            .O(N__42053),
            .I(N__42050));
    LocalMux I__9431 (
            .O(N__42050),
            .I(N__42047));
    Odrv4 I__9430 (
            .O(N__42047),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__9429 (
            .O(N__42044),
            .I(N__42040));
    InMux I__9428 (
            .O(N__42043),
            .I(N__42035));
    LocalMux I__9427 (
            .O(N__42040),
            .I(N__42032));
    InMux I__9426 (
            .O(N__42039),
            .I(N__42027));
    InMux I__9425 (
            .O(N__42038),
            .I(N__42027));
    LocalMux I__9424 (
            .O(N__42035),
            .I(N__42024));
    Span4Mux_v I__9423 (
            .O(N__42032),
            .I(N__42019));
    LocalMux I__9422 (
            .O(N__42027),
            .I(N__42019));
    Odrv4 I__9421 (
            .O(N__42024),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv4 I__9420 (
            .O(N__42019),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__9419 (
            .O(N__42014),
            .I(N__42011));
    LocalMux I__9418 (
            .O(N__42011),
            .I(N__42007));
    InMux I__9417 (
            .O(N__42010),
            .I(N__42004));
    Span4Mux_h I__9416 (
            .O(N__42007),
            .I(N__42000));
    LocalMux I__9415 (
            .O(N__42004),
            .I(N__41997));
    InMux I__9414 (
            .O(N__42003),
            .I(N__41994));
    Odrv4 I__9413 (
            .O(N__42000),
            .I(\current_shift_inst.un4_control_input1_4 ));
    Odrv4 I__9412 (
            .O(N__41997),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__9411 (
            .O(N__41994),
            .I(\current_shift_inst.un4_control_input1_4 ));
    CascadeMux I__9410 (
            .O(N__41987),
            .I(N__41983));
    InMux I__9409 (
            .O(N__41986),
            .I(N__41979));
    InMux I__9408 (
            .O(N__41983),
            .I(N__41976));
    InMux I__9407 (
            .O(N__41982),
            .I(N__41973));
    LocalMux I__9406 (
            .O(N__41979),
            .I(N__41969));
    LocalMux I__9405 (
            .O(N__41976),
            .I(N__41966));
    LocalMux I__9404 (
            .O(N__41973),
            .I(N__41963));
    InMux I__9403 (
            .O(N__41972),
            .I(N__41959));
    Span4Mux_v I__9402 (
            .O(N__41969),
            .I(N__41956));
    Span4Mux_h I__9401 (
            .O(N__41966),
            .I(N__41953));
    Span4Mux_h I__9400 (
            .O(N__41963),
            .I(N__41950));
    InMux I__9399 (
            .O(N__41962),
            .I(N__41947));
    LocalMux I__9398 (
            .O(N__41959),
            .I(N__41943));
    Span4Mux_h I__9397 (
            .O(N__41956),
            .I(N__41938));
    Span4Mux_v I__9396 (
            .O(N__41953),
            .I(N__41938));
    Span4Mux_v I__9395 (
            .O(N__41950),
            .I(N__41935));
    LocalMux I__9394 (
            .O(N__41947),
            .I(N__41932));
    InMux I__9393 (
            .O(N__41946),
            .I(N__41929));
    Span4Mux_v I__9392 (
            .O(N__41943),
            .I(N__41926));
    Span4Mux_v I__9391 (
            .O(N__41938),
            .I(N__41923));
    Sp12to4 I__9390 (
            .O(N__41935),
            .I(N__41918));
    Span12Mux_h I__9389 (
            .O(N__41932),
            .I(N__41918));
    LocalMux I__9388 (
            .O(N__41929),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__9387 (
            .O(N__41926),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__9386 (
            .O(N__41923),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv12 I__9385 (
            .O(N__41918),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    IoInMux I__9384 (
            .O(N__41909),
            .I(N__41906));
    LocalMux I__9383 (
            .O(N__41906),
            .I(N__41903));
    IoSpan4Mux I__9382 (
            .O(N__41903),
            .I(N__41900));
    Sp12to4 I__9381 (
            .O(N__41900),
            .I(N__41896));
    InMux I__9380 (
            .O(N__41899),
            .I(N__41893));
    Odrv12 I__9379 (
            .O(N__41896),
            .I(T01_c));
    LocalMux I__9378 (
            .O(N__41893),
            .I(T01_c));
    InMux I__9377 (
            .O(N__41888),
            .I(N__41884));
    InMux I__9376 (
            .O(N__41887),
            .I(N__41881));
    LocalMux I__9375 (
            .O(N__41884),
            .I(N__41876));
    LocalMux I__9374 (
            .O(N__41881),
            .I(N__41873));
    InMux I__9373 (
            .O(N__41880),
            .I(N__41868));
    InMux I__9372 (
            .O(N__41879),
            .I(N__41868));
    Span4Mux_h I__9371 (
            .O(N__41876),
            .I(N__41865));
    Odrv12 I__9370 (
            .O(N__41873),
            .I(\phase_controller_inst2.hc_time_passed ));
    LocalMux I__9369 (
            .O(N__41868),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv4 I__9368 (
            .O(N__41865),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__9367 (
            .O(N__41858),
            .I(N__41854));
    InMux I__9366 (
            .O(N__41857),
            .I(N__41851));
    LocalMux I__9365 (
            .O(N__41854),
            .I(N__41847));
    LocalMux I__9364 (
            .O(N__41851),
            .I(N__41843));
    InMux I__9363 (
            .O(N__41850),
            .I(N__41840));
    Span4Mux_v I__9362 (
            .O(N__41847),
            .I(N__41837));
    InMux I__9361 (
            .O(N__41846),
            .I(N__41834));
    Span4Mux_h I__9360 (
            .O(N__41843),
            .I(N__41831));
    LocalMux I__9359 (
            .O(N__41840),
            .I(N__41827));
    Sp12to4 I__9358 (
            .O(N__41837),
            .I(N__41822));
    LocalMux I__9357 (
            .O(N__41834),
            .I(N__41822));
    Span4Mux_h I__9356 (
            .O(N__41831),
            .I(N__41819));
    InMux I__9355 (
            .O(N__41830),
            .I(N__41816));
    Span4Mux_v I__9354 (
            .O(N__41827),
            .I(N__41813));
    Odrv12 I__9353 (
            .O(N__41822),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    Odrv4 I__9352 (
            .O(N__41819),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__9351 (
            .O(N__41816),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    Odrv4 I__9350 (
            .O(N__41813),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    IoInMux I__9349 (
            .O(N__41804),
            .I(N__41801));
    LocalMux I__9348 (
            .O(N__41801),
            .I(N__41798));
    Span4Mux_s3_v I__9347 (
            .O(N__41798),
            .I(N__41794));
    InMux I__9346 (
            .O(N__41797),
            .I(N__41791));
    Odrv4 I__9345 (
            .O(N__41794),
            .I(T12_c));
    LocalMux I__9344 (
            .O(N__41791),
            .I(T12_c));
    InMux I__9343 (
            .O(N__41786),
            .I(N__41782));
    InMux I__9342 (
            .O(N__41785),
            .I(N__41779));
    LocalMux I__9341 (
            .O(N__41782),
            .I(N__41775));
    LocalMux I__9340 (
            .O(N__41779),
            .I(N__41772));
    InMux I__9339 (
            .O(N__41778),
            .I(N__41769));
    Span4Mux_v I__9338 (
            .O(N__41775),
            .I(N__41765));
    Span4Mux_v I__9337 (
            .O(N__41772),
            .I(N__41760));
    LocalMux I__9336 (
            .O(N__41769),
            .I(N__41760));
    InMux I__9335 (
            .O(N__41768),
            .I(N__41757));
    Odrv4 I__9334 (
            .O(N__41765),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__9333 (
            .O(N__41760),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    LocalMux I__9332 (
            .O(N__41757),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    CascadeMux I__9331 (
            .O(N__41750),
            .I(N__41746));
    CascadeMux I__9330 (
            .O(N__41749),
            .I(N__41743));
    InMux I__9329 (
            .O(N__41746),
            .I(N__41740));
    InMux I__9328 (
            .O(N__41743),
            .I(N__41737));
    LocalMux I__9327 (
            .O(N__41740),
            .I(N__41734));
    LocalMux I__9326 (
            .O(N__41737),
            .I(N__41730));
    Span4Mux_h I__9325 (
            .O(N__41734),
            .I(N__41727));
    InMux I__9324 (
            .O(N__41733),
            .I(N__41724));
    Odrv4 I__9323 (
            .O(N__41730),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__9322 (
            .O(N__41727),
            .I(\current_shift_inst.un4_control_input1_15 ));
    LocalMux I__9321 (
            .O(N__41724),
            .I(\current_shift_inst.un4_control_input1_15 ));
    InMux I__9320 (
            .O(N__41717),
            .I(N__41712));
    InMux I__9319 (
            .O(N__41716),
            .I(N__41705));
    InMux I__9318 (
            .O(N__41715),
            .I(N__41705));
    LocalMux I__9317 (
            .O(N__41712),
            .I(N__41685));
    InMux I__9316 (
            .O(N__41711),
            .I(N__41682));
    InMux I__9315 (
            .O(N__41710),
            .I(N__41679));
    LocalMux I__9314 (
            .O(N__41705),
            .I(N__41676));
    InMux I__9313 (
            .O(N__41704),
            .I(N__41671));
    InMux I__9312 (
            .O(N__41703),
            .I(N__41671));
    InMux I__9311 (
            .O(N__41702),
            .I(N__41668));
    InMux I__9310 (
            .O(N__41701),
            .I(N__41663));
    InMux I__9309 (
            .O(N__41700),
            .I(N__41663));
    InMux I__9308 (
            .O(N__41699),
            .I(N__41656));
    InMux I__9307 (
            .O(N__41698),
            .I(N__41656));
    InMux I__9306 (
            .O(N__41697),
            .I(N__41656));
    InMux I__9305 (
            .O(N__41696),
            .I(N__41649));
    InMux I__9304 (
            .O(N__41695),
            .I(N__41649));
    InMux I__9303 (
            .O(N__41694),
            .I(N__41649));
    InMux I__9302 (
            .O(N__41693),
            .I(N__41638));
    InMux I__9301 (
            .O(N__41692),
            .I(N__41638));
    InMux I__9300 (
            .O(N__41691),
            .I(N__41638));
    InMux I__9299 (
            .O(N__41690),
            .I(N__41638));
    InMux I__9298 (
            .O(N__41689),
            .I(N__41638));
    InMux I__9297 (
            .O(N__41688),
            .I(N__41635));
    Span12Mux_v I__9296 (
            .O(N__41685),
            .I(N__41630));
    LocalMux I__9295 (
            .O(N__41682),
            .I(N__41630));
    LocalMux I__9294 (
            .O(N__41679),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    Odrv4 I__9293 (
            .O(N__41676),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__9292 (
            .O(N__41671),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__9291 (
            .O(N__41668),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__9290 (
            .O(N__41663),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__9289 (
            .O(N__41656),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__9288 (
            .O(N__41649),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__9287 (
            .O(N__41638),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    LocalMux I__9286 (
            .O(N__41635),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    Odrv12 I__9285 (
            .O(N__41630),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ));
    InMux I__9284 (
            .O(N__41609),
            .I(N__41606));
    LocalMux I__9283 (
            .O(N__41606),
            .I(N__41602));
    CascadeMux I__9282 (
            .O(N__41605),
            .I(N__41598));
    Span12Mux_v I__9281 (
            .O(N__41602),
            .I(N__41595));
    InMux I__9280 (
            .O(N__41601),
            .I(N__41590));
    InMux I__9279 (
            .O(N__41598),
            .I(N__41590));
    Span12Mux_h I__9278 (
            .O(N__41595),
            .I(N__41587));
    LocalMux I__9277 (
            .O(N__41590),
            .I(N__41584));
    Odrv12 I__9276 (
            .O(N__41587),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    Odrv12 I__9275 (
            .O(N__41584),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    CascadeMux I__9274 (
            .O(N__41579),
            .I(N__41576));
    InMux I__9273 (
            .O(N__41576),
            .I(N__41570));
    InMux I__9272 (
            .O(N__41575),
            .I(N__41558));
    InMux I__9271 (
            .O(N__41574),
            .I(N__41558));
    CascadeMux I__9270 (
            .O(N__41573),
            .I(N__41555));
    LocalMux I__9269 (
            .O(N__41570),
            .I(N__41552));
    InMux I__9268 (
            .O(N__41569),
            .I(N__41546));
    InMux I__9267 (
            .O(N__41568),
            .I(N__41541));
    InMux I__9266 (
            .O(N__41567),
            .I(N__41534));
    InMux I__9265 (
            .O(N__41566),
            .I(N__41534));
    InMux I__9264 (
            .O(N__41565),
            .I(N__41534));
    CascadeMux I__9263 (
            .O(N__41564),
            .I(N__41531));
    CascadeMux I__9262 (
            .O(N__41563),
            .I(N__41527));
    LocalMux I__9261 (
            .O(N__41558),
            .I(N__41524));
    InMux I__9260 (
            .O(N__41555),
            .I(N__41515));
    Span4Mux_h I__9259 (
            .O(N__41552),
            .I(N__41512));
    CascadeMux I__9258 (
            .O(N__41551),
            .I(N__41508));
    CascadeMux I__9257 (
            .O(N__41550),
            .I(N__41505));
    CascadeMux I__9256 (
            .O(N__41549),
            .I(N__41501));
    LocalMux I__9255 (
            .O(N__41546),
            .I(N__41493));
    InMux I__9254 (
            .O(N__41545),
            .I(N__41490));
    InMux I__9253 (
            .O(N__41544),
            .I(N__41487));
    LocalMux I__9252 (
            .O(N__41541),
            .I(N__41484));
    LocalMux I__9251 (
            .O(N__41534),
            .I(N__41481));
    InMux I__9250 (
            .O(N__41531),
            .I(N__41478));
    InMux I__9249 (
            .O(N__41530),
            .I(N__41475));
    InMux I__9248 (
            .O(N__41527),
            .I(N__41472));
    Span4Mux_h I__9247 (
            .O(N__41524),
            .I(N__41469));
    InMux I__9246 (
            .O(N__41523),
            .I(N__41464));
    InMux I__9245 (
            .O(N__41522),
            .I(N__41464));
    InMux I__9244 (
            .O(N__41521),
            .I(N__41461));
    InMux I__9243 (
            .O(N__41520),
            .I(N__41454));
    InMux I__9242 (
            .O(N__41519),
            .I(N__41454));
    InMux I__9241 (
            .O(N__41518),
            .I(N__41454));
    LocalMux I__9240 (
            .O(N__41515),
            .I(N__41449));
    Span4Mux_h I__9239 (
            .O(N__41512),
            .I(N__41449));
    InMux I__9238 (
            .O(N__41511),
            .I(N__41444));
    InMux I__9237 (
            .O(N__41508),
            .I(N__41444));
    InMux I__9236 (
            .O(N__41505),
            .I(N__41441));
    InMux I__9235 (
            .O(N__41504),
            .I(N__41434));
    InMux I__9234 (
            .O(N__41501),
            .I(N__41434));
    InMux I__9233 (
            .O(N__41500),
            .I(N__41434));
    InMux I__9232 (
            .O(N__41499),
            .I(N__41425));
    InMux I__9231 (
            .O(N__41498),
            .I(N__41425));
    InMux I__9230 (
            .O(N__41497),
            .I(N__41425));
    InMux I__9229 (
            .O(N__41496),
            .I(N__41425));
    Span4Mux_v I__9228 (
            .O(N__41493),
            .I(N__41416));
    LocalMux I__9227 (
            .O(N__41490),
            .I(N__41416));
    LocalMux I__9226 (
            .O(N__41487),
            .I(N__41416));
    Span4Mux_v I__9225 (
            .O(N__41484),
            .I(N__41416));
    Odrv12 I__9224 (
            .O(N__41481),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__9223 (
            .O(N__41478),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__9222 (
            .O(N__41475),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__9221 (
            .O(N__41472),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    Odrv4 I__9220 (
            .O(N__41469),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__9219 (
            .O(N__41464),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__9218 (
            .O(N__41461),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__9217 (
            .O(N__41454),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    Odrv4 I__9216 (
            .O(N__41449),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__9215 (
            .O(N__41444),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__9214 (
            .O(N__41441),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__9213 (
            .O(N__41434),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    LocalMux I__9212 (
            .O(N__41425),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    Odrv4 I__9211 (
            .O(N__41416),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i ));
    InMux I__9210 (
            .O(N__41387),
            .I(N__41383));
    InMux I__9209 (
            .O(N__41386),
            .I(N__41380));
    LocalMux I__9208 (
            .O(N__41383),
            .I(N__41377));
    LocalMux I__9207 (
            .O(N__41380),
            .I(N__41374));
    Span4Mux_v I__9206 (
            .O(N__41377),
            .I(N__41370));
    Span4Mux_v I__9205 (
            .O(N__41374),
            .I(N__41367));
    InMux I__9204 (
            .O(N__41373),
            .I(N__41364));
    Sp12to4 I__9203 (
            .O(N__41370),
            .I(N__41359));
    Sp12to4 I__9202 (
            .O(N__41367),
            .I(N__41359));
    LocalMux I__9201 (
            .O(N__41364),
            .I(elapsed_time_ns_1_RNI81DJ11_0_2));
    Odrv12 I__9200 (
            .O(N__41359),
            .I(elapsed_time_ns_1_RNI81DJ11_0_2));
    CascadeMux I__9199 (
            .O(N__41354),
            .I(N__41350));
    CascadeMux I__9198 (
            .O(N__41353),
            .I(N__41347));
    InMux I__9197 (
            .O(N__41350),
            .I(N__41344));
    InMux I__9196 (
            .O(N__41347),
            .I(N__41341));
    LocalMux I__9195 (
            .O(N__41344),
            .I(N__41337));
    LocalMux I__9194 (
            .O(N__41341),
            .I(N__41334));
    InMux I__9193 (
            .O(N__41340),
            .I(N__41331));
    Span4Mux_v I__9192 (
            .O(N__41337),
            .I(N__41328));
    Span4Mux_v I__9191 (
            .O(N__41334),
            .I(N__41325));
    LocalMux I__9190 (
            .O(N__41331),
            .I(N__41322));
    Span4Mux_v I__9189 (
            .O(N__41328),
            .I(N__41318));
    Span4Mux_v I__9188 (
            .O(N__41325),
            .I(N__41313));
    Span4Mux_h I__9187 (
            .O(N__41322),
            .I(N__41313));
    InMux I__9186 (
            .O(N__41321),
            .I(N__41310));
    Odrv4 I__9185 (
            .O(N__41318),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    Odrv4 I__9184 (
            .O(N__41313),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__9183 (
            .O(N__41310),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__9182 (
            .O(N__41303),
            .I(N__41299));
    InMux I__9181 (
            .O(N__41302),
            .I(N__41296));
    LocalMux I__9180 (
            .O(N__41299),
            .I(N__41293));
    LocalMux I__9179 (
            .O(N__41296),
            .I(N__41289));
    Span4Mux_h I__9178 (
            .O(N__41293),
            .I(N__41286));
    InMux I__9177 (
            .O(N__41292),
            .I(N__41283));
    Odrv12 I__9176 (
            .O(N__41289),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv4 I__9175 (
            .O(N__41286),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__9174 (
            .O(N__41283),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__9173 (
            .O(N__41276),
            .I(N__41273));
    LocalMux I__9172 (
            .O(N__41273),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    CascadeMux I__9171 (
            .O(N__41270),
            .I(N__41267));
    InMux I__9170 (
            .O(N__41267),
            .I(N__41264));
    LocalMux I__9169 (
            .O(N__41264),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    InMux I__9168 (
            .O(N__41261),
            .I(N__41257));
    CascadeMux I__9167 (
            .O(N__41260),
            .I(N__41254));
    LocalMux I__9166 (
            .O(N__41257),
            .I(N__41250));
    InMux I__9165 (
            .O(N__41254),
            .I(N__41247));
    InMux I__9164 (
            .O(N__41253),
            .I(N__41244));
    Span4Mux_h I__9163 (
            .O(N__41250),
            .I(N__41241));
    LocalMux I__9162 (
            .O(N__41247),
            .I(N__41236));
    LocalMux I__9161 (
            .O(N__41244),
            .I(N__41236));
    Odrv4 I__9160 (
            .O(N__41241),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__9159 (
            .O(N__41236),
            .I(\current_shift_inst.un4_control_input1_18 ));
    CascadeMux I__9158 (
            .O(N__41231),
            .I(N__41228));
    InMux I__9157 (
            .O(N__41228),
            .I(N__41223));
    InMux I__9156 (
            .O(N__41227),
            .I(N__41218));
    InMux I__9155 (
            .O(N__41226),
            .I(N__41218));
    LocalMux I__9154 (
            .O(N__41223),
            .I(N__41215));
    LocalMux I__9153 (
            .O(N__41218),
            .I(N__41212));
    Span4Mux_v I__9152 (
            .O(N__41215),
            .I(N__41206));
    Span4Mux_h I__9151 (
            .O(N__41212),
            .I(N__41206));
    InMux I__9150 (
            .O(N__41211),
            .I(N__41203));
    Odrv4 I__9149 (
            .O(N__41206),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    LocalMux I__9148 (
            .O(N__41203),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__9147 (
            .O(N__41198),
            .I(N__41189));
    InMux I__9146 (
            .O(N__41197),
            .I(N__41189));
    InMux I__9145 (
            .O(N__41196),
            .I(N__41189));
    LocalMux I__9144 (
            .O(N__41189),
            .I(N__41186));
    Span4Mux_v I__9143 (
            .O(N__41186),
            .I(N__41183));
    Span4Mux_v I__9142 (
            .O(N__41183),
            .I(N__41179));
    InMux I__9141 (
            .O(N__41182),
            .I(N__41176));
    Odrv4 I__9140 (
            .O(N__41179),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__9139 (
            .O(N__41176),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    CascadeMux I__9138 (
            .O(N__41171),
            .I(N__41168));
    InMux I__9137 (
            .O(N__41168),
            .I(N__41159));
    InMux I__9136 (
            .O(N__41167),
            .I(N__41159));
    InMux I__9135 (
            .O(N__41166),
            .I(N__41159));
    LocalMux I__9134 (
            .O(N__41159),
            .I(N__41156));
    Span4Mux_h I__9133 (
            .O(N__41156),
            .I(N__41153));
    Odrv4 I__9132 (
            .O(N__41153),
            .I(\current_shift_inst.un4_control_input1_29 ));
    CascadeMux I__9131 (
            .O(N__41150),
            .I(N__41147));
    InMux I__9130 (
            .O(N__41147),
            .I(N__41144));
    LocalMux I__9129 (
            .O(N__41144),
            .I(N__41141));
    Odrv4 I__9128 (
            .O(N__41141),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__9127 (
            .O(N__41138),
            .I(N__41135));
    LocalMux I__9126 (
            .O(N__41135),
            .I(N__41132));
    Odrv4 I__9125 (
            .O(N__41132),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    InMux I__9124 (
            .O(N__41129),
            .I(N__41126));
    LocalMux I__9123 (
            .O(N__41126),
            .I(N__41123));
    Span4Mux_h I__9122 (
            .O(N__41123),
            .I(N__41120));
    Odrv4 I__9121 (
            .O(N__41120),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__9120 (
            .O(N__41117),
            .I(N__41108));
    InMux I__9119 (
            .O(N__41116),
            .I(N__41108));
    InMux I__9118 (
            .O(N__41115),
            .I(N__41108));
    LocalMux I__9117 (
            .O(N__41108),
            .I(N__41105));
    Span4Mux_h I__9116 (
            .O(N__41105),
            .I(N__41102));
    Span4Mux_v I__9115 (
            .O(N__41102),
            .I(N__41098));
    InMux I__9114 (
            .O(N__41101),
            .I(N__41095));
    Odrv4 I__9113 (
            .O(N__41098),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__9112 (
            .O(N__41095),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    CascadeMux I__9111 (
            .O(N__41090),
            .I(N__41087));
    InMux I__9110 (
            .O(N__41087),
            .I(N__41078));
    InMux I__9109 (
            .O(N__41086),
            .I(N__41078));
    InMux I__9108 (
            .O(N__41085),
            .I(N__41078));
    LocalMux I__9107 (
            .O(N__41078),
            .I(N__41075));
    Span4Mux_h I__9106 (
            .O(N__41075),
            .I(N__41072));
    Odrv4 I__9105 (
            .O(N__41072),
            .I(\current_shift_inst.un4_control_input1_22 ));
    CascadeMux I__9104 (
            .O(N__41069),
            .I(N__41066));
    InMux I__9103 (
            .O(N__41066),
            .I(N__41063));
    LocalMux I__9102 (
            .O(N__41063),
            .I(N__41060));
    Odrv4 I__9101 (
            .O(N__41060),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    InMux I__9100 (
            .O(N__41057),
            .I(N__41054));
    LocalMux I__9099 (
            .O(N__41054),
            .I(N__41049));
    InMux I__9098 (
            .O(N__41053),
            .I(N__41046));
    InMux I__9097 (
            .O(N__41052),
            .I(N__41043));
    Span4Mux_h I__9096 (
            .O(N__41049),
            .I(N__41038));
    LocalMux I__9095 (
            .O(N__41046),
            .I(N__41038));
    LocalMux I__9094 (
            .O(N__41043),
            .I(N__41035));
    Span4Mux_v I__9093 (
            .O(N__41038),
            .I(N__41030));
    Span4Mux_h I__9092 (
            .O(N__41035),
            .I(N__41030));
    Span4Mux_v I__9091 (
            .O(N__41030),
            .I(N__41027));
    Odrv4 I__9090 (
            .O(N__41027),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    CEMux I__9089 (
            .O(N__41024),
            .I(N__40997));
    CEMux I__9088 (
            .O(N__41023),
            .I(N__40997));
    CEMux I__9087 (
            .O(N__41022),
            .I(N__40997));
    CEMux I__9086 (
            .O(N__41021),
            .I(N__40997));
    CEMux I__9085 (
            .O(N__41020),
            .I(N__40997));
    CEMux I__9084 (
            .O(N__41019),
            .I(N__40997));
    CEMux I__9083 (
            .O(N__41018),
            .I(N__40997));
    CEMux I__9082 (
            .O(N__41017),
            .I(N__40997));
    CEMux I__9081 (
            .O(N__41016),
            .I(N__40997));
    GlobalMux I__9080 (
            .O(N__40997),
            .I(N__40994));
    gio2CtrlBuf I__9079 (
            .O(N__40994),
            .I(\current_shift_inst.timer_s1.N_166_i_g ));
    InMux I__9078 (
            .O(N__40991),
            .I(N__40988));
    LocalMux I__9077 (
            .O(N__40988),
            .I(N__40985));
    Span4Mux_h I__9076 (
            .O(N__40985),
            .I(N__40982));
    Odrv4 I__9075 (
            .O(N__40982),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__9074 (
            .O(N__40979),
            .I(N__40976));
    LocalMux I__9073 (
            .O(N__40976),
            .I(N__40973));
    Odrv4 I__9072 (
            .O(N__40973),
            .I(\current_shift_inst.control_input_1_axb_6 ));
    InMux I__9071 (
            .O(N__40970),
            .I(N__40967));
    LocalMux I__9070 (
            .O(N__40967),
            .I(N__40964));
    Span4Mux_v I__9069 (
            .O(N__40964),
            .I(N__40961));
    Odrv4 I__9068 (
            .O(N__40961),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__9067 (
            .O(N__40958),
            .I(N__40955));
    LocalMux I__9066 (
            .O(N__40955),
            .I(N__40952));
    Odrv4 I__9065 (
            .O(N__40952),
            .I(\current_shift_inst.control_input_1_axb_8 ));
    InMux I__9064 (
            .O(N__40949),
            .I(N__40946));
    LocalMux I__9063 (
            .O(N__40946),
            .I(N__40943));
    Span4Mux_v I__9062 (
            .O(N__40943),
            .I(N__40940));
    Odrv4 I__9061 (
            .O(N__40940),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__9060 (
            .O(N__40937),
            .I(N__40922));
    InMux I__9059 (
            .O(N__40936),
            .I(N__40913));
    InMux I__9058 (
            .O(N__40935),
            .I(N__40913));
    InMux I__9057 (
            .O(N__40934),
            .I(N__40913));
    InMux I__9056 (
            .O(N__40933),
            .I(N__40913));
    InMux I__9055 (
            .O(N__40932),
            .I(N__40902));
    InMux I__9054 (
            .O(N__40931),
            .I(N__40902));
    InMux I__9053 (
            .O(N__40930),
            .I(N__40902));
    InMux I__9052 (
            .O(N__40929),
            .I(N__40902));
    InMux I__9051 (
            .O(N__40928),
            .I(N__40902));
    InMux I__9050 (
            .O(N__40927),
            .I(N__40895));
    InMux I__9049 (
            .O(N__40926),
            .I(N__40895));
    InMux I__9048 (
            .O(N__40925),
            .I(N__40895));
    LocalMux I__9047 (
            .O(N__40922),
            .I(N__40888));
    LocalMux I__9046 (
            .O(N__40913),
            .I(N__40888));
    LocalMux I__9045 (
            .O(N__40902),
            .I(N__40888));
    LocalMux I__9044 (
            .O(N__40895),
            .I(N__40885));
    Span4Mux_v I__9043 (
            .O(N__40888),
            .I(N__40882));
    Odrv4 I__9042 (
            .O(N__40885),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__9041 (
            .O(N__40882),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__9040 (
            .O(N__40877),
            .I(N__40874));
    LocalMux I__9039 (
            .O(N__40874),
            .I(N__40871));
    Odrv4 I__9038 (
            .O(N__40871),
            .I(\current_shift_inst.control_input_1_axb_9 ));
    InMux I__9037 (
            .O(N__40868),
            .I(N__40864));
    InMux I__9036 (
            .O(N__40867),
            .I(N__40861));
    LocalMux I__9035 (
            .O(N__40864),
            .I(N__40858));
    LocalMux I__9034 (
            .O(N__40861),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__9033 (
            .O(N__40858),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__9032 (
            .O(N__40853),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__9031 (
            .O(N__40850),
            .I(N__40847));
    LocalMux I__9030 (
            .O(N__40847),
            .I(N__40843));
    InMux I__9029 (
            .O(N__40846),
            .I(N__40840));
    Span4Mux_h I__9028 (
            .O(N__40843),
            .I(N__40837));
    LocalMux I__9027 (
            .O(N__40840),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__9026 (
            .O(N__40837),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__9025 (
            .O(N__40832),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__9024 (
            .O(N__40829),
            .I(N__40825));
    InMux I__9023 (
            .O(N__40828),
            .I(N__40822));
    LocalMux I__9022 (
            .O(N__40825),
            .I(N__40819));
    LocalMux I__9021 (
            .O(N__40822),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv12 I__9020 (
            .O(N__40819),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__9019 (
            .O(N__40814),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__9018 (
            .O(N__40811),
            .I(N__40807));
    InMux I__9017 (
            .O(N__40810),
            .I(N__40804));
    LocalMux I__9016 (
            .O(N__40807),
            .I(N__40801));
    LocalMux I__9015 (
            .O(N__40804),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__9014 (
            .O(N__40801),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__9013 (
            .O(N__40796),
            .I(bfn_17_16_0_));
    InMux I__9012 (
            .O(N__40793),
            .I(N__40789));
    InMux I__9011 (
            .O(N__40792),
            .I(N__40786));
    LocalMux I__9010 (
            .O(N__40789),
            .I(N__40783));
    LocalMux I__9009 (
            .O(N__40786),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__9008 (
            .O(N__40783),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__9007 (
            .O(N__40778),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__9006 (
            .O(N__40775),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__9005 (
            .O(N__40772),
            .I(N__40768));
    InMux I__9004 (
            .O(N__40771),
            .I(N__40765));
    LocalMux I__9003 (
            .O(N__40768),
            .I(N__40762));
    LocalMux I__9002 (
            .O(N__40765),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__9001 (
            .O(N__40762),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    CascadeMux I__9000 (
            .O(N__40757),
            .I(N__40754));
    InMux I__8999 (
            .O(N__40754),
            .I(N__40751));
    LocalMux I__8998 (
            .O(N__40751),
            .I(N__40748));
    Odrv4 I__8997 (
            .O(N__40748),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    InMux I__8996 (
            .O(N__40745),
            .I(N__40741));
    InMux I__8995 (
            .O(N__40744),
            .I(N__40738));
    LocalMux I__8994 (
            .O(N__40741),
            .I(N__40735));
    LocalMux I__8993 (
            .O(N__40738),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__8992 (
            .O(N__40735),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__8991 (
            .O(N__40730),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__8990 (
            .O(N__40727),
            .I(N__40723));
    InMux I__8989 (
            .O(N__40726),
            .I(N__40720));
    LocalMux I__8988 (
            .O(N__40723),
            .I(N__40717));
    LocalMux I__8987 (
            .O(N__40720),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__8986 (
            .O(N__40717),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__8985 (
            .O(N__40712),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__8984 (
            .O(N__40709),
            .I(N__40705));
    InMux I__8983 (
            .O(N__40708),
            .I(N__40702));
    LocalMux I__8982 (
            .O(N__40705),
            .I(N__40699));
    LocalMux I__8981 (
            .O(N__40702),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv12 I__8980 (
            .O(N__40699),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__8979 (
            .O(N__40694),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__8978 (
            .O(N__40691),
            .I(N__40687));
    InMux I__8977 (
            .O(N__40690),
            .I(N__40684));
    LocalMux I__8976 (
            .O(N__40687),
            .I(N__40681));
    LocalMux I__8975 (
            .O(N__40684),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv12 I__8974 (
            .O(N__40681),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__8973 (
            .O(N__40676),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__8972 (
            .O(N__40673),
            .I(N__40669));
    InMux I__8971 (
            .O(N__40672),
            .I(N__40666));
    LocalMux I__8970 (
            .O(N__40669),
            .I(N__40663));
    LocalMux I__8969 (
            .O(N__40666),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__8968 (
            .O(N__40663),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__8967 (
            .O(N__40658),
            .I(bfn_17_15_0_));
    InMux I__8966 (
            .O(N__40655),
            .I(N__40651));
    InMux I__8965 (
            .O(N__40654),
            .I(N__40648));
    LocalMux I__8964 (
            .O(N__40651),
            .I(N__40645));
    LocalMux I__8963 (
            .O(N__40648),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__8962 (
            .O(N__40645),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__8961 (
            .O(N__40640),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__8960 (
            .O(N__40637),
            .I(N__40633));
    InMux I__8959 (
            .O(N__40636),
            .I(N__40630));
    LocalMux I__8958 (
            .O(N__40633),
            .I(N__40627));
    LocalMux I__8957 (
            .O(N__40630),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__8956 (
            .O(N__40627),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__8955 (
            .O(N__40622),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__8954 (
            .O(N__40619),
            .I(N__40615));
    InMux I__8953 (
            .O(N__40618),
            .I(N__40612));
    LocalMux I__8952 (
            .O(N__40615),
            .I(N__40609));
    LocalMux I__8951 (
            .O(N__40612),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__8950 (
            .O(N__40609),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__8949 (
            .O(N__40604),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__8948 (
            .O(N__40601),
            .I(N__40597));
    InMux I__8947 (
            .O(N__40600),
            .I(N__40594));
    LocalMux I__8946 (
            .O(N__40597),
            .I(N__40591));
    LocalMux I__8945 (
            .O(N__40594),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__8944 (
            .O(N__40591),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__8943 (
            .O(N__40586),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__8942 (
            .O(N__40583),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_19 ));
    InMux I__8941 (
            .O(N__40580),
            .I(N__40577));
    LocalMux I__8940 (
            .O(N__40577),
            .I(N__40573));
    InMux I__8939 (
            .O(N__40576),
            .I(N__40570));
    Span4Mux_s1_v I__8938 (
            .O(N__40573),
            .I(N__40565));
    LocalMux I__8937 (
            .O(N__40570),
            .I(N__40565));
    Span4Mux_v I__8936 (
            .O(N__40565),
            .I(N__40561));
    InMux I__8935 (
            .O(N__40564),
            .I(N__40558));
    Span4Mux_h I__8934 (
            .O(N__40561),
            .I(N__40555));
    LocalMux I__8933 (
            .O(N__40558),
            .I(N__40552));
    Sp12to4 I__8932 (
            .O(N__40555),
            .I(N__40548));
    Span4Mux_v I__8931 (
            .O(N__40552),
            .I(N__40545));
    InMux I__8930 (
            .O(N__40551),
            .I(N__40542));
    Span12Mux_v I__8929 (
            .O(N__40548),
            .I(N__40539));
    Span4Mux_h I__8928 (
            .O(N__40545),
            .I(N__40534));
    LocalMux I__8927 (
            .O(N__40542),
            .I(N__40534));
    Span12Mux_v I__8926 (
            .O(N__40539),
            .I(N__40531));
    Span4Mux_v I__8925 (
            .O(N__40534),
            .I(N__40528));
    Span12Mux_h I__8924 (
            .O(N__40531),
            .I(N__40525));
    Sp12to4 I__8923 (
            .O(N__40528),
            .I(N__40522));
    Odrv12 I__8922 (
            .O(N__40525),
            .I(start_stop_c));
    Odrv12 I__8921 (
            .O(N__40522),
            .I(start_stop_c));
    InMux I__8920 (
            .O(N__40517),
            .I(N__40514));
    LocalMux I__8919 (
            .O(N__40514),
            .I(N__40510));
    InMux I__8918 (
            .O(N__40513),
            .I(N__40507));
    Span4Mux_v I__8917 (
            .O(N__40510),
            .I(N__40502));
    LocalMux I__8916 (
            .O(N__40507),
            .I(N__40502));
    Span4Mux_h I__8915 (
            .O(N__40502),
            .I(N__40499));
    Odrv4 I__8914 (
            .O(N__40499),
            .I(state_ns_i_a3_1));
    InMux I__8913 (
            .O(N__40496),
            .I(N__40493));
    LocalMux I__8912 (
            .O(N__40493),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ));
    InMux I__8911 (
            .O(N__40490),
            .I(N__40486));
    InMux I__8910 (
            .O(N__40489),
            .I(N__40483));
    LocalMux I__8909 (
            .O(N__40486),
            .I(N__40480));
    LocalMux I__8908 (
            .O(N__40483),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__8907 (
            .O(N__40480),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__8906 (
            .O(N__40475),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ));
    InMux I__8905 (
            .O(N__40472),
            .I(N__40468));
    InMux I__8904 (
            .O(N__40471),
            .I(N__40465));
    LocalMux I__8903 (
            .O(N__40468),
            .I(N__40462));
    LocalMux I__8902 (
            .O(N__40465),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__8901 (
            .O(N__40462),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__8900 (
            .O(N__40457),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__8899 (
            .O(N__40454),
            .I(N__40450));
    InMux I__8898 (
            .O(N__40453),
            .I(N__40447));
    LocalMux I__8897 (
            .O(N__40450),
            .I(N__40444));
    LocalMux I__8896 (
            .O(N__40447),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__8895 (
            .O(N__40444),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__8894 (
            .O(N__40439),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__8893 (
            .O(N__40436),
            .I(N__40433));
    LocalMux I__8892 (
            .O(N__40433),
            .I(N__40430));
    Span4Mux_h I__8891 (
            .O(N__40430),
            .I(N__40427));
    Odrv4 I__8890 (
            .O(N__40427),
            .I(\phase_controller_inst2.stoper_tr.un6_running_12 ));
    CascadeMux I__8889 (
            .O(N__40424),
            .I(N__40421));
    InMux I__8888 (
            .O(N__40421),
            .I(N__40418));
    LocalMux I__8887 (
            .O(N__40418),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    InMux I__8886 (
            .O(N__40415),
            .I(N__40412));
    LocalMux I__8885 (
            .O(N__40412),
            .I(N__40409));
    Span4Mux_h I__8884 (
            .O(N__40409),
            .I(N__40406));
    Odrv4 I__8883 (
            .O(N__40406),
            .I(\phase_controller_inst2.stoper_tr.un6_running_13 ));
    CascadeMux I__8882 (
            .O(N__40403),
            .I(N__40400));
    InMux I__8881 (
            .O(N__40400),
            .I(N__40397));
    LocalMux I__8880 (
            .O(N__40397),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    InMux I__8879 (
            .O(N__40394),
            .I(N__40391));
    LocalMux I__8878 (
            .O(N__40391),
            .I(N__40388));
    Span4Mux_h I__8877 (
            .O(N__40388),
            .I(N__40385));
    Odrv4 I__8876 (
            .O(N__40385),
            .I(\phase_controller_inst2.stoper_tr.un6_running_14 ));
    CascadeMux I__8875 (
            .O(N__40382),
            .I(N__40379));
    InMux I__8874 (
            .O(N__40379),
            .I(N__40376));
    LocalMux I__8873 (
            .O(N__40376),
            .I(N__40373));
    Odrv4 I__8872 (
            .O(N__40373),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    InMux I__8871 (
            .O(N__40370),
            .I(N__40367));
    LocalMux I__8870 (
            .O(N__40367),
            .I(N__40364));
    Span4Mux_v I__8869 (
            .O(N__40364),
            .I(N__40361));
    Odrv4 I__8868 (
            .O(N__40361),
            .I(\phase_controller_inst2.stoper_tr.un6_running_15 ));
    CascadeMux I__8867 (
            .O(N__40358),
            .I(N__40355));
    InMux I__8866 (
            .O(N__40355),
            .I(N__40352));
    LocalMux I__8865 (
            .O(N__40352),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    InMux I__8864 (
            .O(N__40349),
            .I(N__40346));
    LocalMux I__8863 (
            .O(N__40346),
            .I(N__40343));
    Span12Mux_h I__8862 (
            .O(N__40343),
            .I(N__40340));
    Odrv12 I__8861 (
            .O(N__40340),
            .I(\phase_controller_inst2.stoper_tr.un6_running_16 ));
    CascadeMux I__8860 (
            .O(N__40337),
            .I(N__40334));
    InMux I__8859 (
            .O(N__40334),
            .I(N__40331));
    LocalMux I__8858 (
            .O(N__40331),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_16 ));
    InMux I__8857 (
            .O(N__40328),
            .I(N__40325));
    LocalMux I__8856 (
            .O(N__40325),
            .I(N__40322));
    Span4Mux_h I__8855 (
            .O(N__40322),
            .I(N__40319));
    Odrv4 I__8854 (
            .O(N__40319),
            .I(\phase_controller_inst2.stoper_tr.un6_running_17 ));
    CascadeMux I__8853 (
            .O(N__40316),
            .I(N__40313));
    InMux I__8852 (
            .O(N__40313),
            .I(N__40310));
    LocalMux I__8851 (
            .O(N__40310),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_17 ));
    InMux I__8850 (
            .O(N__40307),
            .I(N__40304));
    LocalMux I__8849 (
            .O(N__40304),
            .I(N__40301));
    Span4Mux_h I__8848 (
            .O(N__40301),
            .I(N__40298));
    Odrv4 I__8847 (
            .O(N__40298),
            .I(\phase_controller_inst2.stoper_tr.un6_running_18 ));
    CascadeMux I__8846 (
            .O(N__40295),
            .I(N__40292));
    InMux I__8845 (
            .O(N__40292),
            .I(N__40289));
    LocalMux I__8844 (
            .O(N__40289),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_18 ));
    InMux I__8843 (
            .O(N__40286),
            .I(N__40283));
    LocalMux I__8842 (
            .O(N__40283),
            .I(N__40280));
    Span4Mux_v I__8841 (
            .O(N__40280),
            .I(N__40277));
    Odrv4 I__8840 (
            .O(N__40277),
            .I(\phase_controller_inst2.stoper_tr.un6_running_19 ));
    CascadeMux I__8839 (
            .O(N__40274),
            .I(N__40271));
    InMux I__8838 (
            .O(N__40271),
            .I(N__40268));
    LocalMux I__8837 (
            .O(N__40268),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_19 ));
    InMux I__8836 (
            .O(N__40265),
            .I(N__40262));
    LocalMux I__8835 (
            .O(N__40262),
            .I(N__40259));
    Span4Mux_v I__8834 (
            .O(N__40259),
            .I(N__40256));
    Odrv4 I__8833 (
            .O(N__40256),
            .I(\phase_controller_inst2.stoper_tr.un6_running_4 ));
    CascadeMux I__8832 (
            .O(N__40253),
            .I(N__40250));
    InMux I__8831 (
            .O(N__40250),
            .I(N__40247));
    LocalMux I__8830 (
            .O(N__40247),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    InMux I__8829 (
            .O(N__40244),
            .I(N__40241));
    LocalMux I__8828 (
            .O(N__40241),
            .I(N__40238));
    Span4Mux_v I__8827 (
            .O(N__40238),
            .I(N__40235));
    Odrv4 I__8826 (
            .O(N__40235),
            .I(\phase_controller_inst2.stoper_tr.un6_running_5 ));
    CascadeMux I__8825 (
            .O(N__40232),
            .I(N__40229));
    InMux I__8824 (
            .O(N__40229),
            .I(N__40226));
    LocalMux I__8823 (
            .O(N__40226),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    InMux I__8822 (
            .O(N__40223),
            .I(N__40220));
    LocalMux I__8821 (
            .O(N__40220),
            .I(N__40217));
    Span4Mux_h I__8820 (
            .O(N__40217),
            .I(N__40214));
    Odrv4 I__8819 (
            .O(N__40214),
            .I(\phase_controller_inst2.stoper_tr.un6_running_6 ));
    CascadeMux I__8818 (
            .O(N__40211),
            .I(N__40208));
    InMux I__8817 (
            .O(N__40208),
            .I(N__40205));
    LocalMux I__8816 (
            .O(N__40205),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    InMux I__8815 (
            .O(N__40202),
            .I(N__40199));
    LocalMux I__8814 (
            .O(N__40199),
            .I(N__40196));
    Span4Mux_v I__8813 (
            .O(N__40196),
            .I(N__40193));
    Odrv4 I__8812 (
            .O(N__40193),
            .I(\phase_controller_inst2.stoper_tr.un6_running_7 ));
    CascadeMux I__8811 (
            .O(N__40190),
            .I(N__40187));
    InMux I__8810 (
            .O(N__40187),
            .I(N__40184));
    LocalMux I__8809 (
            .O(N__40184),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    InMux I__8808 (
            .O(N__40181),
            .I(N__40178));
    LocalMux I__8807 (
            .O(N__40178),
            .I(N__40175));
    Span4Mux_h I__8806 (
            .O(N__40175),
            .I(N__40172));
    Odrv4 I__8805 (
            .O(N__40172),
            .I(\phase_controller_inst2.stoper_tr.un6_running_8 ));
    CascadeMux I__8804 (
            .O(N__40169),
            .I(N__40166));
    InMux I__8803 (
            .O(N__40166),
            .I(N__40163));
    LocalMux I__8802 (
            .O(N__40163),
            .I(N__40160));
    Odrv4 I__8801 (
            .O(N__40160),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    InMux I__8800 (
            .O(N__40157),
            .I(N__40154));
    LocalMux I__8799 (
            .O(N__40154),
            .I(N__40151));
    Span4Mux_h I__8798 (
            .O(N__40151),
            .I(N__40148));
    Odrv4 I__8797 (
            .O(N__40148),
            .I(\phase_controller_inst2.stoper_tr.un6_running_9 ));
    CascadeMux I__8796 (
            .O(N__40145),
            .I(N__40142));
    InMux I__8795 (
            .O(N__40142),
            .I(N__40139));
    LocalMux I__8794 (
            .O(N__40139),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    InMux I__8793 (
            .O(N__40136),
            .I(N__40133));
    LocalMux I__8792 (
            .O(N__40133),
            .I(N__40130));
    Span4Mux_h I__8791 (
            .O(N__40130),
            .I(N__40127));
    Odrv4 I__8790 (
            .O(N__40127),
            .I(\phase_controller_inst2.stoper_tr.un6_running_10 ));
    CascadeMux I__8789 (
            .O(N__40124),
            .I(N__40121));
    InMux I__8788 (
            .O(N__40121),
            .I(N__40118));
    LocalMux I__8787 (
            .O(N__40118),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    InMux I__8786 (
            .O(N__40115),
            .I(N__40112));
    LocalMux I__8785 (
            .O(N__40112),
            .I(N__40109));
    Span4Mux_h I__8784 (
            .O(N__40109),
            .I(N__40106));
    Odrv4 I__8783 (
            .O(N__40106),
            .I(\phase_controller_inst2.stoper_tr.un6_running_11 ));
    CascadeMux I__8782 (
            .O(N__40103),
            .I(N__40100));
    InMux I__8781 (
            .O(N__40100),
            .I(N__40097));
    LocalMux I__8780 (
            .O(N__40097),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__8779 (
            .O(N__40094),
            .I(elapsed_time_ns_1_RNI3JIF91_0_29_cascade_));
    InMux I__8778 (
            .O(N__40091),
            .I(N__40088));
    LocalMux I__8777 (
            .O(N__40088),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15 ));
    CascadeMux I__8776 (
            .O(N__40085),
            .I(N__40082));
    InMux I__8775 (
            .O(N__40082),
            .I(N__40077));
    InMux I__8774 (
            .O(N__40081),
            .I(N__40070));
    InMux I__8773 (
            .O(N__40080),
            .I(N__40070));
    LocalMux I__8772 (
            .O(N__40077),
            .I(N__40067));
    InMux I__8771 (
            .O(N__40076),
            .I(N__40062));
    InMux I__8770 (
            .O(N__40075),
            .I(N__40062));
    LocalMux I__8769 (
            .O(N__40070),
            .I(N__40059));
    Odrv4 I__8768 (
            .O(N__40067),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14));
    LocalMux I__8767 (
            .O(N__40062),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14));
    Odrv4 I__8766 (
            .O(N__40059),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14));
    InMux I__8765 (
            .O(N__40052),
            .I(N__40049));
    LocalMux I__8764 (
            .O(N__40049),
            .I(N__40046));
    Span4Mux_h I__8763 (
            .O(N__40046),
            .I(N__40043));
    Odrv4 I__8762 (
            .O(N__40043),
            .I(\phase_controller_inst1.stoper_tr.un6_running_14 ));
    InMux I__8761 (
            .O(N__40040),
            .I(N__40036));
    InMux I__8760 (
            .O(N__40039),
            .I(N__40033));
    LocalMux I__8759 (
            .O(N__40036),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    LocalMux I__8758 (
            .O(N__40033),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    CascadeMux I__8757 (
            .O(N__40028),
            .I(N__40025));
    InMux I__8756 (
            .O(N__40025),
            .I(N__40021));
    InMux I__8755 (
            .O(N__40024),
            .I(N__40018));
    LocalMux I__8754 (
            .O(N__40021),
            .I(N__40014));
    LocalMux I__8753 (
            .O(N__40018),
            .I(N__40011));
    InMux I__8752 (
            .O(N__40017),
            .I(N__40008));
    Odrv4 I__8751 (
            .O(N__40014),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    Odrv4 I__8750 (
            .O(N__40011),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    LocalMux I__8749 (
            .O(N__40008),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    CascadeMux I__8748 (
            .O(N__40001),
            .I(N__39994));
    CascadeMux I__8747 (
            .O(N__40000),
            .I(N__39985));
    CascadeMux I__8746 (
            .O(N__39999),
            .I(N__39982));
    InMux I__8745 (
            .O(N__39998),
            .I(N__39977));
    InMux I__8744 (
            .O(N__39997),
            .I(N__39977));
    InMux I__8743 (
            .O(N__39994),
            .I(N__39974));
    InMux I__8742 (
            .O(N__39993),
            .I(N__39971));
    InMux I__8741 (
            .O(N__39992),
            .I(N__39964));
    InMux I__8740 (
            .O(N__39991),
            .I(N__39964));
    InMux I__8739 (
            .O(N__39990),
            .I(N__39964));
    InMux I__8738 (
            .O(N__39989),
            .I(N__39955));
    InMux I__8737 (
            .O(N__39988),
            .I(N__39955));
    InMux I__8736 (
            .O(N__39985),
            .I(N__39955));
    InMux I__8735 (
            .O(N__39982),
            .I(N__39955));
    LocalMux I__8734 (
            .O(N__39977),
            .I(N__39950));
    LocalMux I__8733 (
            .O(N__39974),
            .I(N__39950));
    LocalMux I__8732 (
            .O(N__39971),
            .I(\phase_controller_inst1.stoper_tr.N_241 ));
    LocalMux I__8731 (
            .O(N__39964),
            .I(\phase_controller_inst1.stoper_tr.N_241 ));
    LocalMux I__8730 (
            .O(N__39955),
            .I(\phase_controller_inst1.stoper_tr.N_241 ));
    Odrv12 I__8729 (
            .O(N__39950),
            .I(\phase_controller_inst1.stoper_tr.N_241 ));
    CascadeMux I__8728 (
            .O(N__39941),
            .I(elapsed_time_ns_1_RNISAHF91_0_13_cascade_));
    InMux I__8727 (
            .O(N__39938),
            .I(N__39935));
    LocalMux I__8726 (
            .O(N__39935),
            .I(N__39932));
    Span4Mux_h I__8725 (
            .O(N__39932),
            .I(N__39929));
    Odrv4 I__8724 (
            .O(N__39929),
            .I(\phase_controller_inst1.stoper_tr.un6_running_13 ));
    InMux I__8723 (
            .O(N__39926),
            .I(N__39923));
    LocalMux I__8722 (
            .O(N__39923),
            .I(N__39920));
    Span4Mux_h I__8721 (
            .O(N__39920),
            .I(N__39914));
    InMux I__8720 (
            .O(N__39919),
            .I(N__39911));
    InMux I__8719 (
            .O(N__39918),
            .I(N__39906));
    InMux I__8718 (
            .O(N__39917),
            .I(N__39906));
    Odrv4 I__8717 (
            .O(N__39914),
            .I(elapsed_time_ns_1_RNIIJ4DM1_0_19));
    LocalMux I__8716 (
            .O(N__39911),
            .I(elapsed_time_ns_1_RNIIJ4DM1_0_19));
    LocalMux I__8715 (
            .O(N__39906),
            .I(elapsed_time_ns_1_RNIIJ4DM1_0_19));
    InMux I__8714 (
            .O(N__39899),
            .I(N__39866));
    InMux I__8713 (
            .O(N__39898),
            .I(N__39866));
    InMux I__8712 (
            .O(N__39897),
            .I(N__39866));
    InMux I__8711 (
            .O(N__39896),
            .I(N__39853));
    InMux I__8710 (
            .O(N__39895),
            .I(N__39853));
    InMux I__8709 (
            .O(N__39894),
            .I(N__39844));
    InMux I__8708 (
            .O(N__39893),
            .I(N__39844));
    InMux I__8707 (
            .O(N__39892),
            .I(N__39844));
    InMux I__8706 (
            .O(N__39891),
            .I(N__39844));
    InMux I__8705 (
            .O(N__39890),
            .I(N__39841));
    InMux I__8704 (
            .O(N__39889),
            .I(N__39836));
    InMux I__8703 (
            .O(N__39888),
            .I(N__39836));
    InMux I__8702 (
            .O(N__39887),
            .I(N__39829));
    InMux I__8701 (
            .O(N__39886),
            .I(N__39829));
    InMux I__8700 (
            .O(N__39885),
            .I(N__39829));
    InMux I__8699 (
            .O(N__39884),
            .I(N__39822));
    InMux I__8698 (
            .O(N__39883),
            .I(N__39822));
    InMux I__8697 (
            .O(N__39882),
            .I(N__39822));
    InMux I__8696 (
            .O(N__39881),
            .I(N__39807));
    InMux I__8695 (
            .O(N__39880),
            .I(N__39807));
    InMux I__8694 (
            .O(N__39879),
            .I(N__39807));
    InMux I__8693 (
            .O(N__39878),
            .I(N__39807));
    InMux I__8692 (
            .O(N__39877),
            .I(N__39807));
    InMux I__8691 (
            .O(N__39876),
            .I(N__39807));
    InMux I__8690 (
            .O(N__39875),
            .I(N__39807));
    InMux I__8689 (
            .O(N__39874),
            .I(N__39802));
    InMux I__8688 (
            .O(N__39873),
            .I(N__39802));
    LocalMux I__8687 (
            .O(N__39866),
            .I(N__39799));
    InMux I__8686 (
            .O(N__39865),
            .I(N__39788));
    InMux I__8685 (
            .O(N__39864),
            .I(N__39788));
    InMux I__8684 (
            .O(N__39863),
            .I(N__39788));
    InMux I__8683 (
            .O(N__39862),
            .I(N__39788));
    InMux I__8682 (
            .O(N__39861),
            .I(N__39788));
    InMux I__8681 (
            .O(N__39860),
            .I(N__39781));
    InMux I__8680 (
            .O(N__39859),
            .I(N__39781));
    InMux I__8679 (
            .O(N__39858),
            .I(N__39781));
    LocalMux I__8678 (
            .O(N__39853),
            .I(N__39772));
    LocalMux I__8677 (
            .O(N__39844),
            .I(N__39772));
    LocalMux I__8676 (
            .O(N__39841),
            .I(N__39772));
    LocalMux I__8675 (
            .O(N__39836),
            .I(N__39772));
    LocalMux I__8674 (
            .O(N__39829),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__8673 (
            .O(N__39822),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__8672 (
            .O(N__39807),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__8671 (
            .O(N__39802),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    Odrv4 I__8670 (
            .O(N__39799),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__8669 (
            .O(N__39788),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__8668 (
            .O(N__39781),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    Odrv4 I__8667 (
            .O(N__39772),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    CascadeMux I__8666 (
            .O(N__39755),
            .I(N__39748));
    CascadeMux I__8665 (
            .O(N__39754),
            .I(N__39745));
    InMux I__8664 (
            .O(N__39753),
            .I(N__39717));
    InMux I__8663 (
            .O(N__39752),
            .I(N__39717));
    InMux I__8662 (
            .O(N__39751),
            .I(N__39717));
    InMux I__8661 (
            .O(N__39748),
            .I(N__39717));
    InMux I__8660 (
            .O(N__39745),
            .I(N__39717));
    InMux I__8659 (
            .O(N__39744),
            .I(N__39703));
    InMux I__8658 (
            .O(N__39743),
            .I(N__39703));
    InMux I__8657 (
            .O(N__39742),
            .I(N__39703));
    InMux I__8656 (
            .O(N__39741),
            .I(N__39703));
    InMux I__8655 (
            .O(N__39740),
            .I(N__39703));
    InMux I__8654 (
            .O(N__39739),
            .I(N__39698));
    InMux I__8653 (
            .O(N__39738),
            .I(N__39698));
    InMux I__8652 (
            .O(N__39737),
            .I(N__39691));
    InMux I__8651 (
            .O(N__39736),
            .I(N__39691));
    InMux I__8650 (
            .O(N__39735),
            .I(N__39691));
    InMux I__8649 (
            .O(N__39734),
            .I(N__39688));
    InMux I__8648 (
            .O(N__39733),
            .I(N__39685));
    InMux I__8647 (
            .O(N__39732),
            .I(N__39678));
    InMux I__8646 (
            .O(N__39731),
            .I(N__39678));
    InMux I__8645 (
            .O(N__39730),
            .I(N__39678));
    CascadeMux I__8644 (
            .O(N__39729),
            .I(N__39674));
    CascadeMux I__8643 (
            .O(N__39728),
            .I(N__39670));
    LocalMux I__8642 (
            .O(N__39717),
            .I(N__39667));
    InMux I__8641 (
            .O(N__39716),
            .I(N__39660));
    InMux I__8640 (
            .O(N__39715),
            .I(N__39660));
    InMux I__8639 (
            .O(N__39714),
            .I(N__39660));
    LocalMux I__8638 (
            .O(N__39703),
            .I(N__39653));
    LocalMux I__8637 (
            .O(N__39698),
            .I(N__39653));
    LocalMux I__8636 (
            .O(N__39691),
            .I(N__39653));
    LocalMux I__8635 (
            .O(N__39688),
            .I(N__39646));
    LocalMux I__8634 (
            .O(N__39685),
            .I(N__39646));
    LocalMux I__8633 (
            .O(N__39678),
            .I(N__39646));
    InMux I__8632 (
            .O(N__39677),
            .I(N__39643));
    InMux I__8631 (
            .O(N__39674),
            .I(N__39636));
    InMux I__8630 (
            .O(N__39673),
            .I(N__39636));
    InMux I__8629 (
            .O(N__39670),
            .I(N__39636));
    Span4Mux_v I__8628 (
            .O(N__39667),
            .I(N__39633));
    LocalMux I__8627 (
            .O(N__39660),
            .I(N__39628));
    Span4Mux_h I__8626 (
            .O(N__39653),
            .I(N__39628));
    Span4Mux_v I__8625 (
            .O(N__39646),
            .I(N__39623));
    LocalMux I__8624 (
            .O(N__39643),
            .I(N__39623));
    LocalMux I__8623 (
            .O(N__39636),
            .I(N__39620));
    Odrv4 I__8622 (
            .O(N__39633),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    Odrv4 I__8621 (
            .O(N__39628),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    Odrv4 I__8620 (
            .O(N__39623),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    Odrv12 I__8619 (
            .O(N__39620),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    InMux I__8618 (
            .O(N__39611),
            .I(N__39608));
    LocalMux I__8617 (
            .O(N__39608),
            .I(N__39605));
    Span4Mux_h I__8616 (
            .O(N__39605),
            .I(N__39602));
    Odrv4 I__8615 (
            .O(N__39602),
            .I(\phase_controller_inst1.stoper_tr.un6_running_19 ));
    CEMux I__8614 (
            .O(N__39599),
            .I(N__39594));
    CEMux I__8613 (
            .O(N__39598),
            .I(N__39591));
    CEMux I__8612 (
            .O(N__39597),
            .I(N__39582));
    LocalMux I__8611 (
            .O(N__39594),
            .I(N__39575));
    LocalMux I__8610 (
            .O(N__39591),
            .I(N__39572));
    InMux I__8609 (
            .O(N__39590),
            .I(N__39563));
    InMux I__8608 (
            .O(N__39589),
            .I(N__39563));
    InMux I__8607 (
            .O(N__39588),
            .I(N__39563));
    InMux I__8606 (
            .O(N__39587),
            .I(N__39563));
    InMux I__8605 (
            .O(N__39586),
            .I(N__39560));
    CEMux I__8604 (
            .O(N__39585),
            .I(N__39557));
    LocalMux I__8603 (
            .O(N__39582),
            .I(N__39554));
    InMux I__8602 (
            .O(N__39581),
            .I(N__39535));
    InMux I__8601 (
            .O(N__39580),
            .I(N__39535));
    InMux I__8600 (
            .O(N__39579),
            .I(N__39535));
    InMux I__8599 (
            .O(N__39578),
            .I(N__39535));
    Span4Mux_v I__8598 (
            .O(N__39575),
            .I(N__39532));
    Span4Mux_h I__8597 (
            .O(N__39572),
            .I(N__39529));
    LocalMux I__8596 (
            .O(N__39563),
            .I(N__39524));
    LocalMux I__8595 (
            .O(N__39560),
            .I(N__39524));
    LocalMux I__8594 (
            .O(N__39557),
            .I(N__39519));
    Span4Mux_h I__8593 (
            .O(N__39554),
            .I(N__39519));
    InMux I__8592 (
            .O(N__39553),
            .I(N__39512));
    InMux I__8591 (
            .O(N__39552),
            .I(N__39512));
    InMux I__8590 (
            .O(N__39551),
            .I(N__39512));
    InMux I__8589 (
            .O(N__39550),
            .I(N__39509));
    InMux I__8588 (
            .O(N__39549),
            .I(N__39504));
    InMux I__8587 (
            .O(N__39548),
            .I(N__39504));
    InMux I__8586 (
            .O(N__39547),
            .I(N__39495));
    InMux I__8585 (
            .O(N__39546),
            .I(N__39495));
    InMux I__8584 (
            .O(N__39545),
            .I(N__39495));
    InMux I__8583 (
            .O(N__39544),
            .I(N__39495));
    LocalMux I__8582 (
            .O(N__39535),
            .I(N__39490));
    Span4Mux_h I__8581 (
            .O(N__39532),
            .I(N__39490));
    Span4Mux_v I__8580 (
            .O(N__39529),
            .I(N__39485));
    Span4Mux_h I__8579 (
            .O(N__39524),
            .I(N__39485));
    Span4Mux_h I__8578 (
            .O(N__39519),
            .I(N__39482));
    LocalMux I__8577 (
            .O(N__39512),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    LocalMux I__8576 (
            .O(N__39509),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    LocalMux I__8575 (
            .O(N__39504),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    LocalMux I__8574 (
            .O(N__39495),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__8573 (
            .O(N__39490),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__8572 (
            .O(N__39485),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__8571 (
            .O(N__39482),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    InMux I__8570 (
            .O(N__39467),
            .I(N__39464));
    LocalMux I__8569 (
            .O(N__39464),
            .I(N__39461));
    Span4Mux_h I__8568 (
            .O(N__39461),
            .I(N__39458));
    Odrv4 I__8567 (
            .O(N__39458),
            .I(\phase_controller_inst2.stoper_tr.un6_running_1 ));
    CascadeMux I__8566 (
            .O(N__39455),
            .I(N__39452));
    InMux I__8565 (
            .O(N__39452),
            .I(N__39449));
    LocalMux I__8564 (
            .O(N__39449),
            .I(N__39446));
    Odrv4 I__8563 (
            .O(N__39446),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    InMux I__8562 (
            .O(N__39443),
            .I(N__39440));
    LocalMux I__8561 (
            .O(N__39440),
            .I(N__39437));
    Span4Mux_h I__8560 (
            .O(N__39437),
            .I(N__39434));
    Odrv4 I__8559 (
            .O(N__39434),
            .I(\phase_controller_inst2.stoper_tr.un6_running_2 ));
    CascadeMux I__8558 (
            .O(N__39431),
            .I(N__39428));
    InMux I__8557 (
            .O(N__39428),
            .I(N__39425));
    LocalMux I__8556 (
            .O(N__39425),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    InMux I__8555 (
            .O(N__39422),
            .I(N__39419));
    LocalMux I__8554 (
            .O(N__39419),
            .I(N__39416));
    Span4Mux_v I__8553 (
            .O(N__39416),
            .I(N__39413));
    Odrv4 I__8552 (
            .O(N__39413),
            .I(\phase_controller_inst2.stoper_tr.un6_running_3 ));
    CascadeMux I__8551 (
            .O(N__39410),
            .I(N__39407));
    InMux I__8550 (
            .O(N__39407),
            .I(N__39404));
    LocalMux I__8549 (
            .O(N__39404),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__8548 (
            .O(N__39401),
            .I(elapsed_time_ns_1_RNITCIF91_0_23_cascade_));
    InMux I__8547 (
            .O(N__39398),
            .I(N__39394));
    InMux I__8546 (
            .O(N__39397),
            .I(N__39391));
    LocalMux I__8545 (
            .O(N__39394),
            .I(elapsed_time_ns_1_RNIRAIF91_0_21));
    LocalMux I__8544 (
            .O(N__39391),
            .I(elapsed_time_ns_1_RNIRAIF91_0_21));
    CascadeMux I__8543 (
            .O(N__39386),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15_cascade_ ));
    InMux I__8542 (
            .O(N__39383),
            .I(N__39379));
    InMux I__8541 (
            .O(N__39382),
            .I(N__39376));
    LocalMux I__8540 (
            .O(N__39379),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    LocalMux I__8539 (
            .O(N__39376),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__8538 (
            .O(N__39371),
            .I(N__39367));
    InMux I__8537 (
            .O(N__39370),
            .I(N__39364));
    LocalMux I__8536 (
            .O(N__39367),
            .I(N__39360));
    LocalMux I__8535 (
            .O(N__39364),
            .I(N__39357));
    CascadeMux I__8534 (
            .O(N__39363),
            .I(N__39353));
    Span4Mux_v I__8533 (
            .O(N__39360),
            .I(N__39348));
    Span4Mux_v I__8532 (
            .O(N__39357),
            .I(N__39348));
    InMux I__8531 (
            .O(N__39356),
            .I(N__39345));
    InMux I__8530 (
            .O(N__39353),
            .I(N__39342));
    Sp12to4 I__8529 (
            .O(N__39348),
            .I(N__39337));
    LocalMux I__8528 (
            .O(N__39345),
            .I(N__39337));
    LocalMux I__8527 (
            .O(N__39342),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    Odrv12 I__8526 (
            .O(N__39337),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    CascadeMux I__8525 (
            .O(N__39332),
            .I(N__39328));
    InMux I__8524 (
            .O(N__39331),
            .I(N__39325));
    InMux I__8523 (
            .O(N__39328),
            .I(N__39322));
    LocalMux I__8522 (
            .O(N__39325),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    LocalMux I__8521 (
            .O(N__39322),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__8520 (
            .O(N__39317),
            .I(N__39311));
    InMux I__8519 (
            .O(N__39316),
            .I(N__39311));
    LocalMux I__8518 (
            .O(N__39311),
            .I(\delay_measurement_inst.delay_tr_timer.N_347 ));
    InMux I__8517 (
            .O(N__39308),
            .I(N__39305));
    LocalMux I__8516 (
            .O(N__39305),
            .I(N__39301));
    InMux I__8515 (
            .O(N__39304),
            .I(N__39298));
    Odrv4 I__8514 (
            .O(N__39301),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    LocalMux I__8513 (
            .O(N__39298),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    CascadeMux I__8512 (
            .O(N__39293),
            .I(N__39290));
    InMux I__8511 (
            .O(N__39290),
            .I(N__39287));
    LocalMux I__8510 (
            .O(N__39287),
            .I(N__39283));
    InMux I__8509 (
            .O(N__39286),
            .I(N__39280));
    Odrv4 I__8508 (
            .O(N__39283),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    LocalMux I__8507 (
            .O(N__39280),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__8506 (
            .O(N__39275),
            .I(N__39269));
    InMux I__8505 (
            .O(N__39274),
            .I(N__39269));
    LocalMux I__8504 (
            .O(N__39269),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    CascadeMux I__8503 (
            .O(N__39266),
            .I(N__39263));
    InMux I__8502 (
            .O(N__39263),
            .I(N__39259));
    InMux I__8501 (
            .O(N__39262),
            .I(N__39256));
    LocalMux I__8500 (
            .O(N__39259),
            .I(N__39253));
    LocalMux I__8499 (
            .O(N__39256),
            .I(N__39247));
    Span4Mux_v I__8498 (
            .O(N__39253),
            .I(N__39247));
    InMux I__8497 (
            .O(N__39252),
            .I(N__39244));
    Odrv4 I__8496 (
            .O(N__39247),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    LocalMux I__8495 (
            .O(N__39244),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    CascadeMux I__8494 (
            .O(N__39239),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11_cascade_));
    CascadeMux I__8493 (
            .O(N__39236),
            .I(N__39233));
    InMux I__8492 (
            .O(N__39233),
            .I(N__39228));
    InMux I__8491 (
            .O(N__39232),
            .I(N__39225));
    CascadeMux I__8490 (
            .O(N__39231),
            .I(N__39222));
    LocalMux I__8489 (
            .O(N__39228),
            .I(N__39217));
    LocalMux I__8488 (
            .O(N__39225),
            .I(N__39217));
    InMux I__8487 (
            .O(N__39222),
            .I(N__39213));
    Span4Mux_v I__8486 (
            .O(N__39217),
            .I(N__39210));
    InMux I__8485 (
            .O(N__39216),
            .I(N__39207));
    LocalMux I__8484 (
            .O(N__39213),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    Odrv4 I__8483 (
            .O(N__39210),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    LocalMux I__8482 (
            .O(N__39207),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    CascadeMux I__8481 (
            .O(N__39200),
            .I(N__39195));
    InMux I__8480 (
            .O(N__39199),
            .I(N__39192));
    InMux I__8479 (
            .O(N__39198),
            .I(N__39189));
    InMux I__8478 (
            .O(N__39195),
            .I(N__39186));
    LocalMux I__8477 (
            .O(N__39192),
            .I(N__39181));
    LocalMux I__8476 (
            .O(N__39189),
            .I(N__39181));
    LocalMux I__8475 (
            .O(N__39186),
            .I(N__39178));
    Span4Mux_v I__8474 (
            .O(N__39181),
            .I(N__39173));
    Span4Mux_v I__8473 (
            .O(N__39178),
            .I(N__39173));
    Odrv4 I__8472 (
            .O(N__39173),
            .I(\phase_controller_inst1.stoper_tr.N_244 ));
    InMux I__8471 (
            .O(N__39170),
            .I(N__39164));
    InMux I__8470 (
            .O(N__39169),
            .I(N__39164));
    LocalMux I__8469 (
            .O(N__39164),
            .I(N__39161));
    Odrv4 I__8468 (
            .O(N__39161),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__8467 (
            .O(N__39158),
            .I(N__39155));
    LocalMux I__8466 (
            .O(N__39155),
            .I(elapsed_time_ns_1_RNI3JIF91_0_29));
    CascadeMux I__8465 (
            .O(N__39152),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ));
    CascadeMux I__8464 (
            .O(N__39149),
            .I(\delay_measurement_inst.delay_tr_timer.N_358_cascade_ ));
    InMux I__8463 (
            .O(N__39146),
            .I(N__39143));
    LocalMux I__8462 (
            .O(N__39143),
            .I(\delay_measurement_inst.delay_tr_timer.N_381 ));
    InMux I__8461 (
            .O(N__39140),
            .I(N__39130));
    InMux I__8460 (
            .O(N__39139),
            .I(N__39127));
    InMux I__8459 (
            .O(N__39138),
            .I(N__39124));
    InMux I__8458 (
            .O(N__39137),
            .I(N__39121));
    InMux I__8457 (
            .O(N__39136),
            .I(N__39118));
    InMux I__8456 (
            .O(N__39135),
            .I(N__39113));
    InMux I__8455 (
            .O(N__39134),
            .I(N__39113));
    InMux I__8454 (
            .O(N__39133),
            .I(N__39110));
    LocalMux I__8453 (
            .O(N__39130),
            .I(N__39104));
    LocalMux I__8452 (
            .O(N__39127),
            .I(N__39104));
    LocalMux I__8451 (
            .O(N__39124),
            .I(N__39099));
    LocalMux I__8450 (
            .O(N__39121),
            .I(N__39099));
    LocalMux I__8449 (
            .O(N__39118),
            .I(N__39094));
    LocalMux I__8448 (
            .O(N__39113),
            .I(N__39094));
    LocalMux I__8447 (
            .O(N__39110),
            .I(N__39091));
    InMux I__8446 (
            .O(N__39109),
            .I(N__39088));
    Span4Mux_h I__8445 (
            .O(N__39104),
            .I(N__39085));
    Span4Mux_h I__8444 (
            .O(N__39099),
            .I(N__39082));
    Span4Mux_h I__8443 (
            .O(N__39094),
            .I(N__39079));
    Odrv12 I__8442 (
            .O(N__39091),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    LocalMux I__8441 (
            .O(N__39088),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    Odrv4 I__8440 (
            .O(N__39085),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    Odrv4 I__8439 (
            .O(N__39082),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    Odrv4 I__8438 (
            .O(N__39079),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    InMux I__8437 (
            .O(N__39068),
            .I(N__39065));
    LocalMux I__8436 (
            .O(N__39065),
            .I(N__39059));
    InMux I__8435 (
            .O(N__39064),
            .I(N__39056));
    InMux I__8434 (
            .O(N__39063),
            .I(N__39051));
    InMux I__8433 (
            .O(N__39062),
            .I(N__39051));
    Odrv4 I__8432 (
            .O(N__39059),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    LocalMux I__8431 (
            .O(N__39056),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    LocalMux I__8430 (
            .O(N__39051),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    InMux I__8429 (
            .O(N__39044),
            .I(N__39041));
    LocalMux I__8428 (
            .O(N__39041),
            .I(N__39037));
    CascadeMux I__8427 (
            .O(N__39040),
            .I(N__39034));
    Span4Mux_v I__8426 (
            .O(N__39037),
            .I(N__39030));
    InMux I__8425 (
            .O(N__39034),
            .I(N__39025));
    InMux I__8424 (
            .O(N__39033),
            .I(N__39025));
    Odrv4 I__8423 (
            .O(N__39030),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    LocalMux I__8422 (
            .O(N__39025),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    CascadeMux I__8421 (
            .O(N__39020),
            .I(\delay_measurement_inst.delay_tr_timer.N_348_cascade_ ));
    InMux I__8420 (
            .O(N__39017),
            .I(N__39014));
    LocalMux I__8419 (
            .O(N__39014),
            .I(N__39008));
    InMux I__8418 (
            .O(N__39013),
            .I(N__39005));
    InMux I__8417 (
            .O(N__39012),
            .I(N__39000));
    InMux I__8416 (
            .O(N__39011),
            .I(N__39000));
    Odrv4 I__8415 (
            .O(N__39008),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    LocalMux I__8414 (
            .O(N__39005),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    LocalMux I__8413 (
            .O(N__39000),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    InMux I__8412 (
            .O(N__38993),
            .I(N__38984));
    InMux I__8411 (
            .O(N__38992),
            .I(N__38984));
    InMux I__8410 (
            .O(N__38991),
            .I(N__38984));
    LocalMux I__8409 (
            .O(N__38984),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__8408 (
            .O(N__38981),
            .I(N__38978));
    LocalMux I__8407 (
            .O(N__38978),
            .I(N__38973));
    InMux I__8406 (
            .O(N__38977),
            .I(N__38970));
    InMux I__8405 (
            .O(N__38976),
            .I(N__38967));
    Span4Mux_h I__8404 (
            .O(N__38973),
            .I(N__38961));
    LocalMux I__8403 (
            .O(N__38970),
            .I(N__38961));
    LocalMux I__8402 (
            .O(N__38967),
            .I(N__38958));
    InMux I__8401 (
            .O(N__38966),
            .I(N__38955));
    Span4Mux_v I__8400 (
            .O(N__38961),
            .I(N__38952));
    Span4Mux_v I__8399 (
            .O(N__38958),
            .I(N__38949));
    LocalMux I__8398 (
            .O(N__38955),
            .I(N__38946));
    Odrv4 I__8397 (
            .O(N__38952),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    Odrv4 I__8396 (
            .O(N__38949),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    Odrv12 I__8395 (
            .O(N__38946),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    InMux I__8394 (
            .O(N__38939),
            .I(N__38936));
    LocalMux I__8393 (
            .O(N__38936),
            .I(elapsed_time_ns_1_RNITCIF91_0_23));
    CascadeMux I__8392 (
            .O(N__38933),
            .I(N__38930));
    InMux I__8391 (
            .O(N__38930),
            .I(N__38926));
    InMux I__8390 (
            .O(N__38929),
            .I(N__38923));
    LocalMux I__8389 (
            .O(N__38926),
            .I(N__38920));
    LocalMux I__8388 (
            .O(N__38923),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__8387 (
            .O(N__38920),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__8386 (
            .O(N__38915),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__8385 (
            .O(N__38912),
            .I(N__38888));
    InMux I__8384 (
            .O(N__38911),
            .I(N__38888));
    InMux I__8383 (
            .O(N__38910),
            .I(N__38888));
    InMux I__8382 (
            .O(N__38909),
            .I(N__38888));
    InMux I__8381 (
            .O(N__38908),
            .I(N__38879));
    InMux I__8380 (
            .O(N__38907),
            .I(N__38879));
    InMux I__8379 (
            .O(N__38906),
            .I(N__38879));
    InMux I__8378 (
            .O(N__38905),
            .I(N__38879));
    InMux I__8377 (
            .O(N__38904),
            .I(N__38856));
    InMux I__8376 (
            .O(N__38903),
            .I(N__38856));
    InMux I__8375 (
            .O(N__38902),
            .I(N__38856));
    InMux I__8374 (
            .O(N__38901),
            .I(N__38856));
    InMux I__8373 (
            .O(N__38900),
            .I(N__38847));
    InMux I__8372 (
            .O(N__38899),
            .I(N__38847));
    InMux I__8371 (
            .O(N__38898),
            .I(N__38847));
    InMux I__8370 (
            .O(N__38897),
            .I(N__38847));
    LocalMux I__8369 (
            .O(N__38888),
            .I(N__38844));
    LocalMux I__8368 (
            .O(N__38879),
            .I(N__38841));
    InMux I__8367 (
            .O(N__38878),
            .I(N__38836));
    InMux I__8366 (
            .O(N__38877),
            .I(N__38836));
    InMux I__8365 (
            .O(N__38876),
            .I(N__38827));
    InMux I__8364 (
            .O(N__38875),
            .I(N__38827));
    InMux I__8363 (
            .O(N__38874),
            .I(N__38827));
    InMux I__8362 (
            .O(N__38873),
            .I(N__38827));
    InMux I__8361 (
            .O(N__38872),
            .I(N__38818));
    InMux I__8360 (
            .O(N__38871),
            .I(N__38818));
    InMux I__8359 (
            .O(N__38870),
            .I(N__38818));
    InMux I__8358 (
            .O(N__38869),
            .I(N__38818));
    InMux I__8357 (
            .O(N__38868),
            .I(N__38809));
    InMux I__8356 (
            .O(N__38867),
            .I(N__38809));
    InMux I__8355 (
            .O(N__38866),
            .I(N__38809));
    InMux I__8354 (
            .O(N__38865),
            .I(N__38809));
    LocalMux I__8353 (
            .O(N__38856),
            .I(N__38804));
    LocalMux I__8352 (
            .O(N__38847),
            .I(N__38804));
    Span4Mux_h I__8351 (
            .O(N__38844),
            .I(N__38799));
    Span4Mux_h I__8350 (
            .O(N__38841),
            .I(N__38799));
    LocalMux I__8349 (
            .O(N__38836),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__8348 (
            .O(N__38827),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__8347 (
            .O(N__38818),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__8346 (
            .O(N__38809),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__8345 (
            .O(N__38804),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__8344 (
            .O(N__38799),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__8343 (
            .O(N__38786),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    InMux I__8342 (
            .O(N__38783),
            .I(N__38779));
    InMux I__8341 (
            .O(N__38782),
            .I(N__38776));
    LocalMux I__8340 (
            .O(N__38779),
            .I(N__38773));
    LocalMux I__8339 (
            .O(N__38776),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__8338 (
            .O(N__38773),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__8337 (
            .O(N__38768),
            .I(N__38763));
    CEMux I__8336 (
            .O(N__38767),
            .I(N__38760));
    CEMux I__8335 (
            .O(N__38766),
            .I(N__38757));
    LocalMux I__8334 (
            .O(N__38763),
            .I(N__38754));
    LocalMux I__8333 (
            .O(N__38760),
            .I(N__38751));
    LocalMux I__8332 (
            .O(N__38757),
            .I(N__38747));
    Span4Mux_v I__8331 (
            .O(N__38754),
            .I(N__38742));
    Span4Mux_h I__8330 (
            .O(N__38751),
            .I(N__38742));
    CEMux I__8329 (
            .O(N__38750),
            .I(N__38739));
    Span4Mux_v I__8328 (
            .O(N__38747),
            .I(N__38732));
    Span4Mux_h I__8327 (
            .O(N__38742),
            .I(N__38732));
    LocalMux I__8326 (
            .O(N__38739),
            .I(N__38732));
    Span4Mux_v I__8325 (
            .O(N__38732),
            .I(N__38729));
    Odrv4 I__8324 (
            .O(N__38729),
            .I(\current_shift_inst.timer_s1.N_167_i ));
    CascadeMux I__8323 (
            .O(N__38726),
            .I(N__38722));
    InMux I__8322 (
            .O(N__38725),
            .I(N__38719));
    InMux I__8321 (
            .O(N__38722),
            .I(N__38716));
    LocalMux I__8320 (
            .O(N__38719),
            .I(N__38710));
    LocalMux I__8319 (
            .O(N__38716),
            .I(N__38710));
    InMux I__8318 (
            .O(N__38715),
            .I(N__38707));
    Span4Mux_v I__8317 (
            .O(N__38710),
            .I(N__38704));
    LocalMux I__8316 (
            .O(N__38707),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    Odrv4 I__8315 (
            .O(N__38704),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    CEMux I__8314 (
            .O(N__38699),
            .I(N__38681));
    CEMux I__8313 (
            .O(N__38698),
            .I(N__38681));
    CEMux I__8312 (
            .O(N__38697),
            .I(N__38681));
    CEMux I__8311 (
            .O(N__38696),
            .I(N__38681));
    CEMux I__8310 (
            .O(N__38695),
            .I(N__38681));
    CEMux I__8309 (
            .O(N__38694),
            .I(N__38681));
    GlobalMux I__8308 (
            .O(N__38681),
            .I(N__38678));
    gio2CtrlBuf I__8307 (
            .O(N__38678),
            .I(\delay_measurement_inst.delay_tr_timer.N_434_i_g ));
    CascadeMux I__8306 (
            .O(N__38675),
            .I(N__38671));
    InMux I__8305 (
            .O(N__38674),
            .I(N__38665));
    InMux I__8304 (
            .O(N__38671),
            .I(N__38665));
    InMux I__8303 (
            .O(N__38670),
            .I(N__38662));
    LocalMux I__8302 (
            .O(N__38665),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__8301 (
            .O(N__38662),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    InMux I__8300 (
            .O(N__38657),
            .I(N__38654));
    LocalMux I__8299 (
            .O(N__38654),
            .I(N__38650));
    CascadeMux I__8298 (
            .O(N__38653),
            .I(N__38647));
    Span4Mux_h I__8297 (
            .O(N__38650),
            .I(N__38644));
    InMux I__8296 (
            .O(N__38647),
            .I(N__38641));
    Odrv4 I__8295 (
            .O(N__38644),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    LocalMux I__8294 (
            .O(N__38641),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    InMux I__8293 (
            .O(N__38636),
            .I(N__38632));
    InMux I__8292 (
            .O(N__38635),
            .I(N__38629));
    LocalMux I__8291 (
            .O(N__38632),
            .I(\delay_measurement_inst.delay_tr_timer.N_341 ));
    LocalMux I__8290 (
            .O(N__38629),
            .I(\delay_measurement_inst.delay_tr_timer.N_341 ));
    CascadeMux I__8289 (
            .O(N__38624),
            .I(N__38620));
    InMux I__8288 (
            .O(N__38623),
            .I(N__38616));
    InMux I__8287 (
            .O(N__38620),
            .I(N__38611));
    InMux I__8286 (
            .O(N__38619),
            .I(N__38611));
    LocalMux I__8285 (
            .O(N__38616),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    LocalMux I__8284 (
            .O(N__38611),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    CascadeMux I__8283 (
            .O(N__38606),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ));
    InMux I__8282 (
            .O(N__38603),
            .I(N__38600));
    LocalMux I__8281 (
            .O(N__38600),
            .I(N__38596));
    InMux I__8280 (
            .O(N__38599),
            .I(N__38593));
    Span4Mux_v I__8279 (
            .O(N__38596),
            .I(N__38585));
    LocalMux I__8278 (
            .O(N__38593),
            .I(N__38585));
    InMux I__8277 (
            .O(N__38592),
            .I(N__38580));
    InMux I__8276 (
            .O(N__38591),
            .I(N__38580));
    InMux I__8275 (
            .O(N__38590),
            .I(N__38577));
    Span4Mux_h I__8274 (
            .O(N__38585),
            .I(N__38574));
    LocalMux I__8273 (
            .O(N__38580),
            .I(N__38571));
    LocalMux I__8272 (
            .O(N__38577),
            .I(elapsed_time_ns_1_RNIRHL2M1_0_3));
    Odrv4 I__8271 (
            .O(N__38574),
            .I(elapsed_time_ns_1_RNIRHL2M1_0_3));
    Odrv12 I__8270 (
            .O(N__38571),
            .I(elapsed_time_ns_1_RNIRHL2M1_0_3));
    CascadeMux I__8269 (
            .O(N__38564),
            .I(\delay_measurement_inst.delay_tr_timer.N_381_cascade_ ));
    InMux I__8268 (
            .O(N__38561),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    CascadeMux I__8267 (
            .O(N__38558),
            .I(N__38554));
    InMux I__8266 (
            .O(N__38557),
            .I(N__38550));
    InMux I__8265 (
            .O(N__38554),
            .I(N__38547));
    InMux I__8264 (
            .O(N__38553),
            .I(N__38544));
    LocalMux I__8263 (
            .O(N__38550),
            .I(N__38539));
    LocalMux I__8262 (
            .O(N__38547),
            .I(N__38539));
    LocalMux I__8261 (
            .O(N__38544),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__8260 (
            .O(N__38539),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__8259 (
            .O(N__38534),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    CascadeMux I__8258 (
            .O(N__38531),
            .I(N__38528));
    InMux I__8257 (
            .O(N__38528),
            .I(N__38523));
    InMux I__8256 (
            .O(N__38527),
            .I(N__38520));
    InMux I__8255 (
            .O(N__38526),
            .I(N__38517));
    LocalMux I__8254 (
            .O(N__38523),
            .I(N__38512));
    LocalMux I__8253 (
            .O(N__38520),
            .I(N__38512));
    LocalMux I__8252 (
            .O(N__38517),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__8251 (
            .O(N__38512),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__8250 (
            .O(N__38507),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    CascadeMux I__8249 (
            .O(N__38504),
            .I(N__38500));
    CascadeMux I__8248 (
            .O(N__38503),
            .I(N__38497));
    InMux I__8247 (
            .O(N__38500),
            .I(N__38491));
    InMux I__8246 (
            .O(N__38497),
            .I(N__38491));
    InMux I__8245 (
            .O(N__38496),
            .I(N__38488));
    LocalMux I__8244 (
            .O(N__38491),
            .I(N__38485));
    LocalMux I__8243 (
            .O(N__38488),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__8242 (
            .O(N__38485),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__8241 (
            .O(N__38480),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__8240 (
            .O(N__38477),
            .I(N__38470));
    InMux I__8239 (
            .O(N__38476),
            .I(N__38470));
    InMux I__8238 (
            .O(N__38475),
            .I(N__38467));
    LocalMux I__8237 (
            .O(N__38470),
            .I(N__38464));
    LocalMux I__8236 (
            .O(N__38467),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__8235 (
            .O(N__38464),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__8234 (
            .O(N__38459),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    CascadeMux I__8233 (
            .O(N__38456),
            .I(N__38453));
    InMux I__8232 (
            .O(N__38453),
            .I(N__38448));
    InMux I__8231 (
            .O(N__38452),
            .I(N__38445));
    InMux I__8230 (
            .O(N__38451),
            .I(N__38442));
    LocalMux I__8229 (
            .O(N__38448),
            .I(N__38437));
    LocalMux I__8228 (
            .O(N__38445),
            .I(N__38437));
    LocalMux I__8227 (
            .O(N__38442),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__8226 (
            .O(N__38437),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__8225 (
            .O(N__38432),
            .I(bfn_16_25_0_));
    CascadeMux I__8224 (
            .O(N__38429),
            .I(N__38425));
    CascadeMux I__8223 (
            .O(N__38428),
            .I(N__38422));
    InMux I__8222 (
            .O(N__38425),
            .I(N__38418));
    InMux I__8221 (
            .O(N__38422),
            .I(N__38415));
    InMux I__8220 (
            .O(N__38421),
            .I(N__38412));
    LocalMux I__8219 (
            .O(N__38418),
            .I(N__38407));
    LocalMux I__8218 (
            .O(N__38415),
            .I(N__38407));
    LocalMux I__8217 (
            .O(N__38412),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__8216 (
            .O(N__38407),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__8215 (
            .O(N__38402),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    InMux I__8214 (
            .O(N__38399),
            .I(N__38392));
    InMux I__8213 (
            .O(N__38398),
            .I(N__38392));
    InMux I__8212 (
            .O(N__38397),
            .I(N__38389));
    LocalMux I__8211 (
            .O(N__38392),
            .I(N__38386));
    LocalMux I__8210 (
            .O(N__38389),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv4 I__8209 (
            .O(N__38386),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__8208 (
            .O(N__38381),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    CascadeMux I__8207 (
            .O(N__38378),
            .I(N__38375));
    InMux I__8206 (
            .O(N__38375),
            .I(N__38370));
    InMux I__8205 (
            .O(N__38374),
            .I(N__38367));
    InMux I__8204 (
            .O(N__38373),
            .I(N__38364));
    LocalMux I__8203 (
            .O(N__38370),
            .I(N__38359));
    LocalMux I__8202 (
            .O(N__38367),
            .I(N__38359));
    LocalMux I__8201 (
            .O(N__38364),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv4 I__8200 (
            .O(N__38359),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__8199 (
            .O(N__38354),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    CascadeMux I__8198 (
            .O(N__38351),
            .I(N__38348));
    InMux I__8197 (
            .O(N__38348),
            .I(N__38343));
    InMux I__8196 (
            .O(N__38347),
            .I(N__38340));
    InMux I__8195 (
            .O(N__38346),
            .I(N__38337));
    LocalMux I__8194 (
            .O(N__38343),
            .I(N__38332));
    LocalMux I__8193 (
            .O(N__38340),
            .I(N__38332));
    LocalMux I__8192 (
            .O(N__38337),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv4 I__8191 (
            .O(N__38332),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__8190 (
            .O(N__38327),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    CascadeMux I__8189 (
            .O(N__38324),
            .I(N__38320));
    InMux I__8188 (
            .O(N__38323),
            .I(N__38316));
    InMux I__8187 (
            .O(N__38320),
            .I(N__38313));
    InMux I__8186 (
            .O(N__38319),
            .I(N__38310));
    LocalMux I__8185 (
            .O(N__38316),
            .I(N__38305));
    LocalMux I__8184 (
            .O(N__38313),
            .I(N__38305));
    LocalMux I__8183 (
            .O(N__38310),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__8182 (
            .O(N__38305),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__8181 (
            .O(N__38300),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__8180 (
            .O(N__38297),
            .I(N__38294));
    InMux I__8179 (
            .O(N__38294),
            .I(N__38289));
    InMux I__8178 (
            .O(N__38293),
            .I(N__38286));
    InMux I__8177 (
            .O(N__38292),
            .I(N__38283));
    LocalMux I__8176 (
            .O(N__38289),
            .I(N__38278));
    LocalMux I__8175 (
            .O(N__38286),
            .I(N__38278));
    LocalMux I__8174 (
            .O(N__38283),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__8173 (
            .O(N__38278),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__8172 (
            .O(N__38273),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    CascadeMux I__8171 (
            .O(N__38270),
            .I(N__38266));
    CascadeMux I__8170 (
            .O(N__38269),
            .I(N__38263));
    InMux I__8169 (
            .O(N__38266),
            .I(N__38257));
    InMux I__8168 (
            .O(N__38263),
            .I(N__38257));
    InMux I__8167 (
            .O(N__38262),
            .I(N__38254));
    LocalMux I__8166 (
            .O(N__38257),
            .I(N__38251));
    LocalMux I__8165 (
            .O(N__38254),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__8164 (
            .O(N__38251),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__8163 (
            .O(N__38246),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__8162 (
            .O(N__38243),
            .I(N__38236));
    InMux I__8161 (
            .O(N__38242),
            .I(N__38236));
    InMux I__8160 (
            .O(N__38241),
            .I(N__38233));
    LocalMux I__8159 (
            .O(N__38236),
            .I(N__38230));
    LocalMux I__8158 (
            .O(N__38233),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__8157 (
            .O(N__38230),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__8156 (
            .O(N__38225),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__8155 (
            .O(N__38222),
            .I(N__38219));
    InMux I__8154 (
            .O(N__38219),
            .I(N__38214));
    InMux I__8153 (
            .O(N__38218),
            .I(N__38211));
    InMux I__8152 (
            .O(N__38217),
            .I(N__38208));
    LocalMux I__8151 (
            .O(N__38214),
            .I(N__38203));
    LocalMux I__8150 (
            .O(N__38211),
            .I(N__38203));
    LocalMux I__8149 (
            .O(N__38208),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__8148 (
            .O(N__38203),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__8147 (
            .O(N__38198),
            .I(bfn_16_24_0_));
    CascadeMux I__8146 (
            .O(N__38195),
            .I(N__38191));
    CascadeMux I__8145 (
            .O(N__38194),
            .I(N__38188));
    InMux I__8144 (
            .O(N__38191),
            .I(N__38185));
    InMux I__8143 (
            .O(N__38188),
            .I(N__38181));
    LocalMux I__8142 (
            .O(N__38185),
            .I(N__38178));
    InMux I__8141 (
            .O(N__38184),
            .I(N__38175));
    LocalMux I__8140 (
            .O(N__38181),
            .I(N__38170));
    Span4Mux_h I__8139 (
            .O(N__38178),
            .I(N__38170));
    LocalMux I__8138 (
            .O(N__38175),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__8137 (
            .O(N__38170),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__8136 (
            .O(N__38165),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__8135 (
            .O(N__38162),
            .I(N__38155));
    InMux I__8134 (
            .O(N__38161),
            .I(N__38155));
    InMux I__8133 (
            .O(N__38160),
            .I(N__38152));
    LocalMux I__8132 (
            .O(N__38155),
            .I(N__38149));
    LocalMux I__8131 (
            .O(N__38152),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__8130 (
            .O(N__38149),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__8129 (
            .O(N__38144),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    CascadeMux I__8128 (
            .O(N__38141),
            .I(N__38138));
    InMux I__8127 (
            .O(N__38138),
            .I(N__38133));
    InMux I__8126 (
            .O(N__38137),
            .I(N__38130));
    InMux I__8125 (
            .O(N__38136),
            .I(N__38127));
    LocalMux I__8124 (
            .O(N__38133),
            .I(N__38122));
    LocalMux I__8123 (
            .O(N__38130),
            .I(N__38122));
    LocalMux I__8122 (
            .O(N__38127),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv4 I__8121 (
            .O(N__38122),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    CascadeMux I__8120 (
            .O(N__38117),
            .I(N__38114));
    InMux I__8119 (
            .O(N__38114),
            .I(N__38109));
    InMux I__8118 (
            .O(N__38113),
            .I(N__38106));
    InMux I__8117 (
            .O(N__38112),
            .I(N__38103));
    LocalMux I__8116 (
            .O(N__38109),
            .I(N__38098));
    LocalMux I__8115 (
            .O(N__38106),
            .I(N__38098));
    LocalMux I__8114 (
            .O(N__38103),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__8113 (
            .O(N__38098),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__8112 (
            .O(N__38093),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    InMux I__8111 (
            .O(N__38090),
            .I(N__38083));
    InMux I__8110 (
            .O(N__38089),
            .I(N__38083));
    InMux I__8109 (
            .O(N__38088),
            .I(N__38080));
    LocalMux I__8108 (
            .O(N__38083),
            .I(N__38077));
    LocalMux I__8107 (
            .O(N__38080),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__8106 (
            .O(N__38077),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__8105 (
            .O(N__38072),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__8104 (
            .O(N__38069),
            .I(N__38066));
    InMux I__8103 (
            .O(N__38066),
            .I(N__38061));
    InMux I__8102 (
            .O(N__38065),
            .I(N__38058));
    InMux I__8101 (
            .O(N__38064),
            .I(N__38055));
    LocalMux I__8100 (
            .O(N__38061),
            .I(N__38050));
    LocalMux I__8099 (
            .O(N__38058),
            .I(N__38050));
    LocalMux I__8098 (
            .O(N__38055),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__8097 (
            .O(N__38050),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__8096 (
            .O(N__38045),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    CascadeMux I__8095 (
            .O(N__38042),
            .I(N__38038));
    CascadeMux I__8094 (
            .O(N__38041),
            .I(N__38035));
    InMux I__8093 (
            .O(N__38038),
            .I(N__38029));
    InMux I__8092 (
            .O(N__38035),
            .I(N__38029));
    InMux I__8091 (
            .O(N__38034),
            .I(N__38026));
    LocalMux I__8090 (
            .O(N__38029),
            .I(N__38023));
    LocalMux I__8089 (
            .O(N__38026),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__8088 (
            .O(N__38023),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__8087 (
            .O(N__38018),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__8086 (
            .O(N__38015),
            .I(N__38008));
    InMux I__8085 (
            .O(N__38014),
            .I(N__38008));
    InMux I__8084 (
            .O(N__38013),
            .I(N__38005));
    LocalMux I__8083 (
            .O(N__38008),
            .I(N__38002));
    LocalMux I__8082 (
            .O(N__38005),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__8081 (
            .O(N__38002),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__8080 (
            .O(N__37997),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__8079 (
            .O(N__37994),
            .I(N__37991));
    InMux I__8078 (
            .O(N__37991),
            .I(N__37986));
    InMux I__8077 (
            .O(N__37990),
            .I(N__37983));
    InMux I__8076 (
            .O(N__37989),
            .I(N__37980));
    LocalMux I__8075 (
            .O(N__37986),
            .I(N__37975));
    LocalMux I__8074 (
            .O(N__37983),
            .I(N__37975));
    LocalMux I__8073 (
            .O(N__37980),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__8072 (
            .O(N__37975),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__8071 (
            .O(N__37970),
            .I(bfn_16_23_0_));
    CascadeMux I__8070 (
            .O(N__37967),
            .I(N__37963));
    CascadeMux I__8069 (
            .O(N__37966),
            .I(N__37960));
    InMux I__8068 (
            .O(N__37963),
            .I(N__37956));
    InMux I__8067 (
            .O(N__37960),
            .I(N__37953));
    InMux I__8066 (
            .O(N__37959),
            .I(N__37950));
    LocalMux I__8065 (
            .O(N__37956),
            .I(N__37945));
    LocalMux I__8064 (
            .O(N__37953),
            .I(N__37945));
    LocalMux I__8063 (
            .O(N__37950),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__8062 (
            .O(N__37945),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__8061 (
            .O(N__37940),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    InMux I__8060 (
            .O(N__37937),
            .I(N__37930));
    InMux I__8059 (
            .O(N__37936),
            .I(N__37930));
    InMux I__8058 (
            .O(N__37935),
            .I(N__37927));
    LocalMux I__8057 (
            .O(N__37930),
            .I(N__37924));
    LocalMux I__8056 (
            .O(N__37927),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__8055 (
            .O(N__37924),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__8054 (
            .O(N__37919),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    CascadeMux I__8053 (
            .O(N__37916),
            .I(N__37908));
    CascadeMux I__8052 (
            .O(N__37915),
            .I(N__37904));
    CascadeMux I__8051 (
            .O(N__37914),
            .I(N__37900));
    CascadeMux I__8050 (
            .O(N__37913),
            .I(N__37892));
    CascadeMux I__8049 (
            .O(N__37912),
            .I(N__37888));
    InMux I__8048 (
            .O(N__37911),
            .I(N__37864));
    InMux I__8047 (
            .O(N__37908),
            .I(N__37864));
    InMux I__8046 (
            .O(N__37907),
            .I(N__37864));
    InMux I__8045 (
            .O(N__37904),
            .I(N__37864));
    InMux I__8044 (
            .O(N__37903),
            .I(N__37864));
    InMux I__8043 (
            .O(N__37900),
            .I(N__37864));
    InMux I__8042 (
            .O(N__37899),
            .I(N__37864));
    InMux I__8041 (
            .O(N__37898),
            .I(N__37859));
    InMux I__8040 (
            .O(N__37897),
            .I(N__37859));
    InMux I__8039 (
            .O(N__37896),
            .I(N__37846));
    InMux I__8038 (
            .O(N__37895),
            .I(N__37846));
    InMux I__8037 (
            .O(N__37892),
            .I(N__37846));
    InMux I__8036 (
            .O(N__37891),
            .I(N__37846));
    InMux I__8035 (
            .O(N__37888),
            .I(N__37846));
    InMux I__8034 (
            .O(N__37887),
            .I(N__37846));
    CascadeMux I__8033 (
            .O(N__37886),
            .I(N__37843));
    CascadeMux I__8032 (
            .O(N__37885),
            .I(N__37839));
    CascadeMux I__8031 (
            .O(N__37884),
            .I(N__37835));
    CascadeMux I__8030 (
            .O(N__37883),
            .I(N__37831));
    CascadeMux I__8029 (
            .O(N__37882),
            .I(N__37826));
    CascadeMux I__8028 (
            .O(N__37881),
            .I(N__37822));
    CascadeMux I__8027 (
            .O(N__37880),
            .I(N__37818));
    InMux I__8026 (
            .O(N__37879),
            .I(N__37814));
    LocalMux I__8025 (
            .O(N__37864),
            .I(N__37796));
    LocalMux I__8024 (
            .O(N__37859),
            .I(N__37796));
    LocalMux I__8023 (
            .O(N__37846),
            .I(N__37796));
    InMux I__8022 (
            .O(N__37843),
            .I(N__37779));
    InMux I__8021 (
            .O(N__37842),
            .I(N__37779));
    InMux I__8020 (
            .O(N__37839),
            .I(N__37779));
    InMux I__8019 (
            .O(N__37838),
            .I(N__37779));
    InMux I__8018 (
            .O(N__37835),
            .I(N__37779));
    InMux I__8017 (
            .O(N__37834),
            .I(N__37779));
    InMux I__8016 (
            .O(N__37831),
            .I(N__37779));
    InMux I__8015 (
            .O(N__37830),
            .I(N__37779));
    InMux I__8014 (
            .O(N__37829),
            .I(N__37764));
    InMux I__8013 (
            .O(N__37826),
            .I(N__37764));
    InMux I__8012 (
            .O(N__37825),
            .I(N__37764));
    InMux I__8011 (
            .O(N__37822),
            .I(N__37764));
    InMux I__8010 (
            .O(N__37821),
            .I(N__37764));
    InMux I__8009 (
            .O(N__37818),
            .I(N__37764));
    InMux I__8008 (
            .O(N__37817),
            .I(N__37764));
    LocalMux I__8007 (
            .O(N__37814),
            .I(N__37759));
    InMux I__8006 (
            .O(N__37813),
            .I(N__37756));
    InMux I__8005 (
            .O(N__37812),
            .I(N__37753));
    InMux I__8004 (
            .O(N__37811),
            .I(N__37750));
    InMux I__8003 (
            .O(N__37810),
            .I(N__37747));
    InMux I__8002 (
            .O(N__37809),
            .I(N__37740));
    InMux I__8001 (
            .O(N__37808),
            .I(N__37740));
    InMux I__8000 (
            .O(N__37807),
            .I(N__37740));
    InMux I__7999 (
            .O(N__37806),
            .I(N__37731));
    InMux I__7998 (
            .O(N__37805),
            .I(N__37731));
    InMux I__7997 (
            .O(N__37804),
            .I(N__37731));
    InMux I__7996 (
            .O(N__37803),
            .I(N__37731));
    Span4Mux_v I__7995 (
            .O(N__37796),
            .I(N__37715));
    LocalMux I__7994 (
            .O(N__37779),
            .I(N__37715));
    LocalMux I__7993 (
            .O(N__37764),
            .I(N__37715));
    InMux I__7992 (
            .O(N__37763),
            .I(N__37710));
    InMux I__7991 (
            .O(N__37762),
            .I(N__37710));
    Span12Mux_s2_h I__7990 (
            .O(N__37759),
            .I(N__37707));
    LocalMux I__7989 (
            .O(N__37756),
            .I(N__37700));
    LocalMux I__7988 (
            .O(N__37753),
            .I(N__37700));
    LocalMux I__7987 (
            .O(N__37750),
            .I(N__37700));
    LocalMux I__7986 (
            .O(N__37747),
            .I(N__37693));
    LocalMux I__7985 (
            .O(N__37740),
            .I(N__37693));
    LocalMux I__7984 (
            .O(N__37731),
            .I(N__37693));
    InMux I__7983 (
            .O(N__37730),
            .I(N__37690));
    InMux I__7982 (
            .O(N__37729),
            .I(N__37683));
    InMux I__7981 (
            .O(N__37728),
            .I(N__37683));
    InMux I__7980 (
            .O(N__37727),
            .I(N__37683));
    InMux I__7979 (
            .O(N__37726),
            .I(N__37674));
    InMux I__7978 (
            .O(N__37725),
            .I(N__37674));
    InMux I__7977 (
            .O(N__37724),
            .I(N__37674));
    InMux I__7976 (
            .O(N__37723),
            .I(N__37674));
    CascadeMux I__7975 (
            .O(N__37722),
            .I(N__37670));
    Span4Mux_v I__7974 (
            .O(N__37715),
            .I(N__37664));
    LocalMux I__7973 (
            .O(N__37710),
            .I(N__37664));
    Span12Mux_v I__7972 (
            .O(N__37707),
            .I(N__37661));
    Span12Mux_s8_v I__7971 (
            .O(N__37700),
            .I(N__37650));
    Span12Mux_s9_v I__7970 (
            .O(N__37693),
            .I(N__37650));
    LocalMux I__7969 (
            .O(N__37690),
            .I(N__37650));
    LocalMux I__7968 (
            .O(N__37683),
            .I(N__37650));
    LocalMux I__7967 (
            .O(N__37674),
            .I(N__37650));
    InMux I__7966 (
            .O(N__37673),
            .I(N__37643));
    InMux I__7965 (
            .O(N__37670),
            .I(N__37643));
    InMux I__7964 (
            .O(N__37669),
            .I(N__37643));
    Span4Mux_v I__7963 (
            .O(N__37664),
            .I(N__37640));
    Span12Mux_h I__7962 (
            .O(N__37661),
            .I(N__37637));
    Span12Mux_v I__7961 (
            .O(N__37650),
            .I(N__37632));
    LocalMux I__7960 (
            .O(N__37643),
            .I(N__37632));
    Span4Mux_h I__7959 (
            .O(N__37640),
            .I(N__37629));
    Odrv12 I__7958 (
            .O(N__37637),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__7957 (
            .O(N__37632),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__7956 (
            .O(N__37629),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__7955 (
            .O(N__37622),
            .I(N__37619));
    InMux I__7954 (
            .O(N__37619),
            .I(N__37616));
    LocalMux I__7953 (
            .O(N__37616),
            .I(N__37613));
    Span4Mux_h I__7952 (
            .O(N__37613),
            .I(N__37610));
    Odrv4 I__7951 (
            .O(N__37610),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__7950 (
            .O(N__37607),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    InMux I__7949 (
            .O(N__37604),
            .I(N__37601));
    LocalMux I__7948 (
            .O(N__37601),
            .I(N__37598));
    Odrv4 I__7947 (
            .O(N__37598),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    CascadeMux I__7946 (
            .O(N__37595),
            .I(N__37592));
    InMux I__7945 (
            .O(N__37592),
            .I(N__37589));
    LocalMux I__7944 (
            .O(N__37589),
            .I(N__37586));
    Odrv4 I__7943 (
            .O(N__37586),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__7942 (
            .O(N__37583),
            .I(N__37580));
    LocalMux I__7941 (
            .O(N__37580),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    InMux I__7940 (
            .O(N__37577),
            .I(N__37574));
    LocalMux I__7939 (
            .O(N__37574),
            .I(N__37571));
    Span4Mux_h I__7938 (
            .O(N__37571),
            .I(N__37568));
    Odrv4 I__7937 (
            .O(N__37568),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__7936 (
            .O(N__37565),
            .I(N__37562));
    LocalMux I__7935 (
            .O(N__37562),
            .I(N__37559));
    Span4Mux_v I__7934 (
            .O(N__37559),
            .I(N__37555));
    InMux I__7933 (
            .O(N__37558),
            .I(N__37551));
    Span4Mux_h I__7932 (
            .O(N__37555),
            .I(N__37548));
    InMux I__7931 (
            .O(N__37554),
            .I(N__37545));
    LocalMux I__7930 (
            .O(N__37551),
            .I(N__37542));
    Odrv4 I__7929 (
            .O(N__37548),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__7928 (
            .O(N__37545),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv4 I__7927 (
            .O(N__37542),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__7926 (
            .O(N__37535),
            .I(bfn_16_22_0_));
    InMux I__7925 (
            .O(N__37532),
            .I(N__37529));
    LocalMux I__7924 (
            .O(N__37529),
            .I(N__37525));
    CascadeMux I__7923 (
            .O(N__37528),
            .I(N__37522));
    Span4Mux_v I__7922 (
            .O(N__37525),
            .I(N__37519));
    InMux I__7921 (
            .O(N__37522),
            .I(N__37515));
    Span4Mux_h I__7920 (
            .O(N__37519),
            .I(N__37512));
    InMux I__7919 (
            .O(N__37518),
            .I(N__37509));
    LocalMux I__7918 (
            .O(N__37515),
            .I(N__37506));
    Odrv4 I__7917 (
            .O(N__37512),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__7916 (
            .O(N__37509),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__7915 (
            .O(N__37506),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__7914 (
            .O(N__37499),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    CascadeMux I__7913 (
            .O(N__37496),
            .I(N__37492));
    CascadeMux I__7912 (
            .O(N__37495),
            .I(N__37489));
    InMux I__7911 (
            .O(N__37492),
            .I(N__37484));
    InMux I__7910 (
            .O(N__37489),
            .I(N__37484));
    LocalMux I__7909 (
            .O(N__37484),
            .I(N__37480));
    InMux I__7908 (
            .O(N__37483),
            .I(N__37477));
    Span12Mux_h I__7907 (
            .O(N__37480),
            .I(N__37474));
    LocalMux I__7906 (
            .O(N__37477),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv12 I__7905 (
            .O(N__37474),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__7904 (
            .O(N__37469),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    CascadeMux I__7903 (
            .O(N__37466),
            .I(N__37463));
    InMux I__7902 (
            .O(N__37463),
            .I(N__37460));
    LocalMux I__7901 (
            .O(N__37460),
            .I(N__37457));
    Span4Mux_v I__7900 (
            .O(N__37457),
            .I(N__37454));
    Span4Mux_h I__7899 (
            .O(N__37454),
            .I(N__37451));
    Odrv4 I__7898 (
            .O(N__37451),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__7897 (
            .O(N__37448),
            .I(N__37445));
    LocalMux I__7896 (
            .O(N__37445),
            .I(N__37442));
    Span4Mux_h I__7895 (
            .O(N__37442),
            .I(N__37439));
    Span4Mux_v I__7894 (
            .O(N__37439),
            .I(N__37436));
    Odrv4 I__7893 (
            .O(N__37436),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    InMux I__7892 (
            .O(N__37433),
            .I(N__37430));
    LocalMux I__7891 (
            .O(N__37430),
            .I(N__37427));
    Span4Mux_h I__7890 (
            .O(N__37427),
            .I(N__37424));
    Odrv4 I__7889 (
            .O(N__37424),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    CascadeMux I__7888 (
            .O(N__37421),
            .I(N__37418));
    InMux I__7887 (
            .O(N__37418),
            .I(N__37415));
    LocalMux I__7886 (
            .O(N__37415),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__7885 (
            .O(N__37412),
            .I(N__37409));
    LocalMux I__7884 (
            .O(N__37409),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    CascadeMux I__7883 (
            .O(N__37406),
            .I(N__37403));
    InMux I__7882 (
            .O(N__37403),
            .I(N__37400));
    LocalMux I__7881 (
            .O(N__37400),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    CascadeMux I__7880 (
            .O(N__37397),
            .I(N__37394));
    InMux I__7879 (
            .O(N__37394),
            .I(N__37391));
    LocalMux I__7878 (
            .O(N__37391),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    InMux I__7877 (
            .O(N__37388),
            .I(N__37385));
    LocalMux I__7876 (
            .O(N__37385),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    CascadeMux I__7875 (
            .O(N__37382),
            .I(N__37379));
    InMux I__7874 (
            .O(N__37379),
            .I(N__37376));
    LocalMux I__7873 (
            .O(N__37376),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    InMux I__7872 (
            .O(N__37373),
            .I(N__37370));
    LocalMux I__7871 (
            .O(N__37370),
            .I(N__37367));
    Span4Mux_h I__7870 (
            .O(N__37367),
            .I(N__37364));
    Odrv4 I__7869 (
            .O(N__37364),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    CascadeMux I__7868 (
            .O(N__37361),
            .I(N__37358));
    InMux I__7867 (
            .O(N__37358),
            .I(N__37355));
    LocalMux I__7866 (
            .O(N__37355),
            .I(N__37352));
    Span12Mux_v I__7865 (
            .O(N__37352),
            .I(N__37349));
    Odrv12 I__7864 (
            .O(N__37349),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__7863 (
            .O(N__37346),
            .I(N__37343));
    LocalMux I__7862 (
            .O(N__37343),
            .I(N__37340));
    Span4Mux_v I__7861 (
            .O(N__37340),
            .I(N__37337));
    Odrv4 I__7860 (
            .O(N__37337),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    CascadeMux I__7859 (
            .O(N__37334),
            .I(N__37331));
    InMux I__7858 (
            .O(N__37331),
            .I(N__37328));
    LocalMux I__7857 (
            .O(N__37328),
            .I(N__37325));
    Span4Mux_h I__7856 (
            .O(N__37325),
            .I(N__37322));
    Odrv4 I__7855 (
            .O(N__37322),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    InMux I__7854 (
            .O(N__37319),
            .I(N__37316));
    LocalMux I__7853 (
            .O(N__37316),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    CascadeMux I__7852 (
            .O(N__37313),
            .I(N__37310));
    InMux I__7851 (
            .O(N__37310),
            .I(N__37307));
    LocalMux I__7850 (
            .O(N__37307),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    InMux I__7849 (
            .O(N__37304),
            .I(N__37301));
    LocalMux I__7848 (
            .O(N__37301),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    InMux I__7847 (
            .O(N__37298),
            .I(N__37295));
    LocalMux I__7846 (
            .O(N__37295),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    CascadeMux I__7845 (
            .O(N__37292),
            .I(N__37289));
    InMux I__7844 (
            .O(N__37289),
            .I(N__37286));
    LocalMux I__7843 (
            .O(N__37286),
            .I(\current_shift_inst.control_input_1_axb_1 ));
    InMux I__7842 (
            .O(N__37283),
            .I(N__37280));
    LocalMux I__7841 (
            .O(N__37280),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__7840 (
            .O(N__37277),
            .I(N__37274));
    LocalMux I__7839 (
            .O(N__37274),
            .I(\current_shift_inst.control_input_1_axb_7 ));
    InMux I__7838 (
            .O(N__37271),
            .I(N__37268));
    LocalMux I__7837 (
            .O(N__37268),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__7836 (
            .O(N__37265),
            .I(N__37262));
    LocalMux I__7835 (
            .O(N__37262),
            .I(\current_shift_inst.control_input_1_axb_10 ));
    InMux I__7834 (
            .O(N__37259),
            .I(N__37256));
    LocalMux I__7833 (
            .O(N__37256),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__7832 (
            .O(N__37253),
            .I(N__37250));
    LocalMux I__7831 (
            .O(N__37250),
            .I(\current_shift_inst.control_input_1_axb_2 ));
    InMux I__7830 (
            .O(N__37247),
            .I(N__37244));
    LocalMux I__7829 (
            .O(N__37244),
            .I(N__37241));
    Span4Mux_h I__7828 (
            .O(N__37241),
            .I(N__37237));
    InMux I__7827 (
            .O(N__37240),
            .I(N__37234));
    Span4Mux_v I__7826 (
            .O(N__37237),
            .I(N__37231));
    LocalMux I__7825 (
            .O(N__37234),
            .I(N__37228));
    Odrv4 I__7824 (
            .O(N__37231),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    Odrv12 I__7823 (
            .O(N__37228),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    CascadeMux I__7822 (
            .O(N__37223),
            .I(N__37220));
    InMux I__7821 (
            .O(N__37220),
            .I(N__37217));
    LocalMux I__7820 (
            .O(N__37217),
            .I(N__37212));
    InMux I__7819 (
            .O(N__37216),
            .I(N__37207));
    InMux I__7818 (
            .O(N__37215),
            .I(N__37207));
    Odrv12 I__7817 (
            .O(N__37212),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    LocalMux I__7816 (
            .O(N__37207),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    CascadeMux I__7815 (
            .O(N__37202),
            .I(N__37199));
    InMux I__7814 (
            .O(N__37199),
            .I(N__37196));
    LocalMux I__7813 (
            .O(N__37196),
            .I(N__37193));
    Odrv12 I__7812 (
            .O(N__37193),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__7811 (
            .O(N__37190),
            .I(N__37187));
    LocalMux I__7810 (
            .O(N__37187),
            .I(N__37184));
    Span4Mux_h I__7809 (
            .O(N__37184),
            .I(N__37181));
    Odrv4 I__7808 (
            .O(N__37181),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    CascadeMux I__7807 (
            .O(N__37178),
            .I(N__37175));
    InMux I__7806 (
            .O(N__37175),
            .I(N__37172));
    LocalMux I__7805 (
            .O(N__37172),
            .I(N__37169));
    Odrv4 I__7804 (
            .O(N__37169),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__7803 (
            .O(N__37166),
            .I(N__37163));
    LocalMux I__7802 (
            .O(N__37163),
            .I(N__37160));
    Odrv12 I__7801 (
            .O(N__37160),
            .I(\current_shift_inst.control_inputZ0Z_3 ));
    InMux I__7800 (
            .O(N__37157),
            .I(\current_shift_inst.control_input_1_cry_2 ));
    InMux I__7799 (
            .O(N__37154),
            .I(N__37151));
    LocalMux I__7798 (
            .O(N__37151),
            .I(\current_shift_inst.control_input_1_axb_4 ));
    InMux I__7797 (
            .O(N__37148),
            .I(N__37145));
    LocalMux I__7796 (
            .O(N__37145),
            .I(N__37142));
    Span12Mux_v I__7795 (
            .O(N__37142),
            .I(N__37139));
    Odrv12 I__7794 (
            .O(N__37139),
            .I(\current_shift_inst.control_inputZ0Z_4 ));
    InMux I__7793 (
            .O(N__37136),
            .I(\current_shift_inst.control_input_1_cry_3 ));
    InMux I__7792 (
            .O(N__37133),
            .I(N__37130));
    LocalMux I__7791 (
            .O(N__37130),
            .I(\current_shift_inst.control_input_1_axb_5 ));
    InMux I__7790 (
            .O(N__37127),
            .I(N__37124));
    LocalMux I__7789 (
            .O(N__37124),
            .I(N__37121));
    Span4Mux_v I__7788 (
            .O(N__37121),
            .I(N__37118));
    Span4Mux_h I__7787 (
            .O(N__37118),
            .I(N__37115));
    Odrv4 I__7786 (
            .O(N__37115),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    InMux I__7785 (
            .O(N__37112),
            .I(\current_shift_inst.control_input_1_cry_4 ));
    InMux I__7784 (
            .O(N__37109),
            .I(N__37106));
    LocalMux I__7783 (
            .O(N__37106),
            .I(N__37103));
    Odrv12 I__7782 (
            .O(N__37103),
            .I(\current_shift_inst.control_inputZ0Z_6 ));
    InMux I__7781 (
            .O(N__37100),
            .I(\current_shift_inst.control_input_1_cry_5 ));
    InMux I__7780 (
            .O(N__37097),
            .I(N__37094));
    LocalMux I__7779 (
            .O(N__37094),
            .I(N__37091));
    Span4Mux_h I__7778 (
            .O(N__37091),
            .I(N__37088));
    Span4Mux_h I__7777 (
            .O(N__37088),
            .I(N__37085));
    Odrv4 I__7776 (
            .O(N__37085),
            .I(\current_shift_inst.control_inputZ0Z_7 ));
    InMux I__7775 (
            .O(N__37082),
            .I(\current_shift_inst.control_input_1_cry_6 ));
    InMux I__7774 (
            .O(N__37079),
            .I(N__37076));
    LocalMux I__7773 (
            .O(N__37076),
            .I(N__37073));
    Span4Mux_h I__7772 (
            .O(N__37073),
            .I(N__37070));
    Odrv4 I__7771 (
            .O(N__37070),
            .I(\current_shift_inst.control_inputZ0Z_8 ));
    InMux I__7770 (
            .O(N__37067),
            .I(bfn_16_16_0_));
    InMux I__7769 (
            .O(N__37064),
            .I(\current_shift_inst.control_input_1_cry_8 ));
    InMux I__7768 (
            .O(N__37061),
            .I(N__37058));
    LocalMux I__7767 (
            .O(N__37058),
            .I(N__37055));
    Span4Mux_v I__7766 (
            .O(N__37055),
            .I(N__37052));
    Odrv4 I__7765 (
            .O(N__37052),
            .I(\current_shift_inst.control_inputZ0Z_10 ));
    InMux I__7764 (
            .O(N__37049),
            .I(\current_shift_inst.control_input_1_cry_9 ));
    InMux I__7763 (
            .O(N__37046),
            .I(N__37043));
    LocalMux I__7762 (
            .O(N__37043),
            .I(\current_shift_inst.control_input_1_axb_11 ));
    InMux I__7761 (
            .O(N__37040),
            .I(\current_shift_inst.control_input_1_cry_10 ));
    InMux I__7760 (
            .O(N__37037),
            .I(N__37034));
    LocalMux I__7759 (
            .O(N__37034),
            .I(N__37030));
    InMux I__7758 (
            .O(N__37033),
            .I(N__37027));
    Span12Mux_s9_h I__7757 (
            .O(N__37030),
            .I(N__37024));
    LocalMux I__7756 (
            .O(N__37027),
            .I(N__37021));
    Odrv12 I__7755 (
            .O(N__37024),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    Odrv4 I__7754 (
            .O(N__37021),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    InMux I__7753 (
            .O(N__37016),
            .I(N__37013));
    LocalMux I__7752 (
            .O(N__37013),
            .I(N__37010));
    Odrv4 I__7751 (
            .O(N__37010),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__7750 (
            .O(N__37007),
            .I(N__37004));
    LocalMux I__7749 (
            .O(N__37004),
            .I(N__37001));
    Odrv4 I__7748 (
            .O(N__37001),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__7747 (
            .O(N__36998),
            .I(N__36995));
    LocalMux I__7746 (
            .O(N__36995),
            .I(N__36992));
    Span12Mux_v I__7745 (
            .O(N__36992),
            .I(N__36989));
    Odrv12 I__7744 (
            .O(N__36989),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    CascadeMux I__7743 (
            .O(N__36986),
            .I(N__36982));
    InMux I__7742 (
            .O(N__36985),
            .I(N__36978));
    InMux I__7741 (
            .O(N__36982),
            .I(N__36975));
    InMux I__7740 (
            .O(N__36981),
            .I(N__36972));
    LocalMux I__7739 (
            .O(N__36978),
            .I(N__36969));
    LocalMux I__7738 (
            .O(N__36975),
            .I(N__36966));
    LocalMux I__7737 (
            .O(N__36972),
            .I(N__36963));
    Span4Mux_h I__7736 (
            .O(N__36969),
            .I(N__36960));
    Span4Mux_v I__7735 (
            .O(N__36966),
            .I(N__36955));
    Span4Mux_h I__7734 (
            .O(N__36963),
            .I(N__36955));
    Odrv4 I__7733 (
            .O(N__36960),
            .I(\current_shift_inst.un4_control_input1_8 ));
    Odrv4 I__7732 (
            .O(N__36955),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__7731 (
            .O(N__36950),
            .I(N__36947));
    LocalMux I__7730 (
            .O(N__36947),
            .I(N__36944));
    Odrv4 I__7729 (
            .O(N__36944),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__7728 (
            .O(N__36941),
            .I(N__36938));
    LocalMux I__7727 (
            .O(N__36938),
            .I(\current_shift_inst.control_input_1_axb_0 ));
    InMux I__7726 (
            .O(N__36935),
            .I(N__36931));
    CascadeMux I__7725 (
            .O(N__36934),
            .I(N__36928));
    LocalMux I__7724 (
            .O(N__36931),
            .I(N__36925));
    InMux I__7723 (
            .O(N__36928),
            .I(N__36922));
    Odrv4 I__7722 (
            .O(N__36925),
            .I(\current_shift_inst.N_1572_i ));
    LocalMux I__7721 (
            .O(N__36922),
            .I(\current_shift_inst.N_1572_i ));
    InMux I__7720 (
            .O(N__36917),
            .I(N__36913));
    InMux I__7719 (
            .O(N__36916),
            .I(N__36910));
    LocalMux I__7718 (
            .O(N__36913),
            .I(N__36905));
    LocalMux I__7717 (
            .O(N__36910),
            .I(N__36905));
    Span12Mux_h I__7716 (
            .O(N__36905),
            .I(N__36902));
    Odrv12 I__7715 (
            .O(N__36902),
            .I(\current_shift_inst.control_inputZ0Z_0 ));
    InMux I__7714 (
            .O(N__36899),
            .I(N__36896));
    LocalMux I__7713 (
            .O(N__36896),
            .I(N__36893));
    Span4Mux_h I__7712 (
            .O(N__36893),
            .I(N__36890));
    Span4Mux_h I__7711 (
            .O(N__36890),
            .I(N__36887));
    Span4Mux_h I__7710 (
            .O(N__36887),
            .I(N__36884));
    Odrv4 I__7709 (
            .O(N__36884),
            .I(\current_shift_inst.control_inputZ0Z_1 ));
    InMux I__7708 (
            .O(N__36881),
            .I(\current_shift_inst.control_input_1_cry_0 ));
    InMux I__7707 (
            .O(N__36878),
            .I(N__36875));
    LocalMux I__7706 (
            .O(N__36875),
            .I(N__36872));
    Span4Mux_v I__7705 (
            .O(N__36872),
            .I(N__36869));
    Span4Mux_h I__7704 (
            .O(N__36869),
            .I(N__36866));
    Odrv4 I__7703 (
            .O(N__36866),
            .I(\current_shift_inst.control_inputZ0Z_2 ));
    InMux I__7702 (
            .O(N__36863),
            .I(\current_shift_inst.control_input_1_cry_1 ));
    InMux I__7701 (
            .O(N__36860),
            .I(N__36857));
    LocalMux I__7700 (
            .O(N__36857),
            .I(\current_shift_inst.control_input_1_axb_3 ));
    InMux I__7699 (
            .O(N__36854),
            .I(N__36850));
    InMux I__7698 (
            .O(N__36853),
            .I(N__36847));
    LocalMux I__7697 (
            .O(N__36850),
            .I(N__36844));
    LocalMux I__7696 (
            .O(N__36847),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    Odrv4 I__7695 (
            .O(N__36844),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__7694 (
            .O(N__36839),
            .I(N__36836));
    InMux I__7693 (
            .O(N__36836),
            .I(N__36831));
    InMux I__7692 (
            .O(N__36835),
            .I(N__36828));
    InMux I__7691 (
            .O(N__36834),
            .I(N__36825));
    LocalMux I__7690 (
            .O(N__36831),
            .I(N__36820));
    LocalMux I__7689 (
            .O(N__36828),
            .I(N__36820));
    LocalMux I__7688 (
            .O(N__36825),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    Odrv4 I__7687 (
            .O(N__36820),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__7686 (
            .O(N__36815),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__7685 (
            .O(N__36812),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    IoInMux I__7684 (
            .O(N__36809),
            .I(N__36806));
    LocalMux I__7683 (
            .O(N__36806),
            .I(N__36803));
    Span12Mux_s8_v I__7682 (
            .O(N__36803),
            .I(N__36799));
    InMux I__7681 (
            .O(N__36802),
            .I(N__36796));
    Odrv12 I__7680 (
            .O(N__36799),
            .I(T45_c));
    LocalMux I__7679 (
            .O(N__36796),
            .I(T45_c));
    CascadeMux I__7678 (
            .O(N__36791),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ));
    InMux I__7677 (
            .O(N__36788),
            .I(N__36785));
    LocalMux I__7676 (
            .O(N__36785),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    InMux I__7675 (
            .O(N__36782),
            .I(N__36779));
    LocalMux I__7674 (
            .O(N__36779),
            .I(N__36776));
    Odrv4 I__7673 (
            .O(N__36776),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    CascadeMux I__7672 (
            .O(N__36773),
            .I(N__36769));
    InMux I__7671 (
            .O(N__36772),
            .I(N__36765));
    InMux I__7670 (
            .O(N__36769),
            .I(N__36762));
    InMux I__7669 (
            .O(N__36768),
            .I(N__36759));
    LocalMux I__7668 (
            .O(N__36765),
            .I(N__36756));
    LocalMux I__7667 (
            .O(N__36762),
            .I(N__36751));
    LocalMux I__7666 (
            .O(N__36759),
            .I(N__36751));
    Span4Mux_v I__7665 (
            .O(N__36756),
            .I(N__36747));
    Span4Mux_h I__7664 (
            .O(N__36751),
            .I(N__36744));
    InMux I__7663 (
            .O(N__36750),
            .I(N__36741));
    Odrv4 I__7662 (
            .O(N__36747),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__7661 (
            .O(N__36744),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    LocalMux I__7660 (
            .O(N__36741),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__7659 (
            .O(N__36734),
            .I(N__36731));
    LocalMux I__7658 (
            .O(N__36731),
            .I(N__36728));
    Span4Mux_v I__7657 (
            .O(N__36728),
            .I(N__36723));
    InMux I__7656 (
            .O(N__36727),
            .I(N__36718));
    InMux I__7655 (
            .O(N__36726),
            .I(N__36718));
    Odrv4 I__7654 (
            .O(N__36723),
            .I(\current_shift_inst.un4_control_input1_7 ));
    LocalMux I__7653 (
            .O(N__36718),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__7652 (
            .O(N__36713),
            .I(N__36706));
    InMux I__7651 (
            .O(N__36712),
            .I(N__36706));
    InMux I__7650 (
            .O(N__36711),
            .I(N__36703));
    LocalMux I__7649 (
            .O(N__36706),
            .I(N__36700));
    LocalMux I__7648 (
            .O(N__36703),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    Odrv4 I__7647 (
            .O(N__36700),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__7646 (
            .O(N__36695),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__7645 (
            .O(N__36692),
            .I(N__36685));
    InMux I__7644 (
            .O(N__36691),
            .I(N__36685));
    InMux I__7643 (
            .O(N__36690),
            .I(N__36682));
    LocalMux I__7642 (
            .O(N__36685),
            .I(N__36679));
    LocalMux I__7641 (
            .O(N__36682),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    Odrv4 I__7640 (
            .O(N__36679),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__7639 (
            .O(N__36674),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__7638 (
            .O(N__36671),
            .I(N__36667));
    InMux I__7637 (
            .O(N__36670),
            .I(N__36663));
    InMux I__7636 (
            .O(N__36667),
            .I(N__36660));
    InMux I__7635 (
            .O(N__36666),
            .I(N__36657));
    LocalMux I__7634 (
            .O(N__36663),
            .I(N__36652));
    LocalMux I__7633 (
            .O(N__36660),
            .I(N__36652));
    LocalMux I__7632 (
            .O(N__36657),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    Odrv4 I__7631 (
            .O(N__36652),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__7630 (
            .O(N__36647),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__7629 (
            .O(N__36644),
            .I(N__36640));
    InMux I__7628 (
            .O(N__36643),
            .I(N__36636));
    InMux I__7627 (
            .O(N__36640),
            .I(N__36633));
    InMux I__7626 (
            .O(N__36639),
            .I(N__36630));
    LocalMux I__7625 (
            .O(N__36636),
            .I(N__36625));
    LocalMux I__7624 (
            .O(N__36633),
            .I(N__36625));
    LocalMux I__7623 (
            .O(N__36630),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    Odrv4 I__7622 (
            .O(N__36625),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__7621 (
            .O(N__36620),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__7620 (
            .O(N__36617),
            .I(N__36613));
    CascadeMux I__7619 (
            .O(N__36616),
            .I(N__36610));
    InMux I__7618 (
            .O(N__36613),
            .I(N__36604));
    InMux I__7617 (
            .O(N__36610),
            .I(N__36604));
    InMux I__7616 (
            .O(N__36609),
            .I(N__36601));
    LocalMux I__7615 (
            .O(N__36604),
            .I(N__36598));
    LocalMux I__7614 (
            .O(N__36601),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    Odrv4 I__7613 (
            .O(N__36598),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__7612 (
            .O(N__36593),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__7611 (
            .O(N__36590),
            .I(N__36586));
    CascadeMux I__7610 (
            .O(N__36589),
            .I(N__36583));
    InMux I__7609 (
            .O(N__36586),
            .I(N__36577));
    InMux I__7608 (
            .O(N__36583),
            .I(N__36577));
    InMux I__7607 (
            .O(N__36582),
            .I(N__36574));
    LocalMux I__7606 (
            .O(N__36577),
            .I(N__36571));
    LocalMux I__7605 (
            .O(N__36574),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    Odrv4 I__7604 (
            .O(N__36571),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__7603 (
            .O(N__36566),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__7602 (
            .O(N__36563),
            .I(N__36560));
    InMux I__7601 (
            .O(N__36560),
            .I(N__36557));
    LocalMux I__7600 (
            .O(N__36557),
            .I(N__36552));
    InMux I__7599 (
            .O(N__36556),
            .I(N__36549));
    InMux I__7598 (
            .O(N__36555),
            .I(N__36546));
    Span4Mux_v I__7597 (
            .O(N__36552),
            .I(N__36543));
    LocalMux I__7596 (
            .O(N__36549),
            .I(N__36540));
    LocalMux I__7595 (
            .O(N__36546),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__7594 (
            .O(N__36543),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__7593 (
            .O(N__36540),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__7592 (
            .O(N__36533),
            .I(bfn_16_11_0_));
    CascadeMux I__7591 (
            .O(N__36530),
            .I(N__36527));
    InMux I__7590 (
            .O(N__36527),
            .I(N__36524));
    LocalMux I__7589 (
            .O(N__36524),
            .I(N__36519));
    InMux I__7588 (
            .O(N__36523),
            .I(N__36516));
    InMux I__7587 (
            .O(N__36522),
            .I(N__36513));
    Span4Mux_v I__7586 (
            .O(N__36519),
            .I(N__36508));
    LocalMux I__7585 (
            .O(N__36516),
            .I(N__36508));
    LocalMux I__7584 (
            .O(N__36513),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv4 I__7583 (
            .O(N__36508),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__7582 (
            .O(N__36503),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__7581 (
            .O(N__36500),
            .I(N__36493));
    InMux I__7580 (
            .O(N__36499),
            .I(N__36493));
    InMux I__7579 (
            .O(N__36498),
            .I(N__36490));
    LocalMux I__7578 (
            .O(N__36493),
            .I(N__36487));
    LocalMux I__7577 (
            .O(N__36490),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    Odrv4 I__7576 (
            .O(N__36487),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    CascadeMux I__7575 (
            .O(N__36482),
            .I(N__36479));
    InMux I__7574 (
            .O(N__36479),
            .I(N__36476));
    LocalMux I__7573 (
            .O(N__36476),
            .I(N__36472));
    InMux I__7572 (
            .O(N__36475),
            .I(N__36469));
    Span4Mux_h I__7571 (
            .O(N__36472),
            .I(N__36466));
    LocalMux I__7570 (
            .O(N__36469),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    Odrv4 I__7569 (
            .O(N__36466),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__7568 (
            .O(N__36461),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__7567 (
            .O(N__36458),
            .I(N__36451));
    InMux I__7566 (
            .O(N__36457),
            .I(N__36451));
    InMux I__7565 (
            .O(N__36456),
            .I(N__36448));
    LocalMux I__7564 (
            .O(N__36451),
            .I(N__36445));
    LocalMux I__7563 (
            .O(N__36448),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    Odrv4 I__7562 (
            .O(N__36445),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__7561 (
            .O(N__36440),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__7560 (
            .O(N__36437),
            .I(N__36434));
    InMux I__7559 (
            .O(N__36434),
            .I(N__36429));
    InMux I__7558 (
            .O(N__36433),
            .I(N__36426));
    InMux I__7557 (
            .O(N__36432),
            .I(N__36423));
    LocalMux I__7556 (
            .O(N__36429),
            .I(N__36418));
    LocalMux I__7555 (
            .O(N__36426),
            .I(N__36418));
    LocalMux I__7554 (
            .O(N__36423),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    Odrv4 I__7553 (
            .O(N__36418),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__7552 (
            .O(N__36413),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__7551 (
            .O(N__36410),
            .I(N__36406));
    InMux I__7550 (
            .O(N__36409),
            .I(N__36402));
    InMux I__7549 (
            .O(N__36406),
            .I(N__36399));
    InMux I__7548 (
            .O(N__36405),
            .I(N__36396));
    LocalMux I__7547 (
            .O(N__36402),
            .I(N__36391));
    LocalMux I__7546 (
            .O(N__36399),
            .I(N__36391));
    LocalMux I__7545 (
            .O(N__36396),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    Odrv4 I__7544 (
            .O(N__36391),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__7543 (
            .O(N__36386),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__7542 (
            .O(N__36383),
            .I(N__36376));
    InMux I__7541 (
            .O(N__36382),
            .I(N__36376));
    InMux I__7540 (
            .O(N__36381),
            .I(N__36373));
    LocalMux I__7539 (
            .O(N__36376),
            .I(N__36370));
    LocalMux I__7538 (
            .O(N__36373),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    Odrv4 I__7537 (
            .O(N__36370),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__7536 (
            .O(N__36365),
            .I(N__36360));
    InMux I__7535 (
            .O(N__36364),
            .I(N__36355));
    InMux I__7534 (
            .O(N__36363),
            .I(N__36355));
    LocalMux I__7533 (
            .O(N__36360),
            .I(N__36352));
    LocalMux I__7532 (
            .O(N__36355),
            .I(N__36349));
    Odrv4 I__7531 (
            .O(N__36352),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    Odrv4 I__7530 (
            .O(N__36349),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__7529 (
            .O(N__36344),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__7528 (
            .O(N__36341),
            .I(N__36337));
    CascadeMux I__7527 (
            .O(N__36340),
            .I(N__36334));
    InMux I__7526 (
            .O(N__36337),
            .I(N__36328));
    InMux I__7525 (
            .O(N__36334),
            .I(N__36328));
    InMux I__7524 (
            .O(N__36333),
            .I(N__36325));
    LocalMux I__7523 (
            .O(N__36328),
            .I(N__36322));
    LocalMux I__7522 (
            .O(N__36325),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv4 I__7521 (
            .O(N__36322),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    CascadeMux I__7520 (
            .O(N__36317),
            .I(N__36313));
    InMux I__7519 (
            .O(N__36316),
            .I(N__36310));
    InMux I__7518 (
            .O(N__36313),
            .I(N__36306));
    LocalMux I__7517 (
            .O(N__36310),
            .I(N__36303));
    InMux I__7516 (
            .O(N__36309),
            .I(N__36300));
    LocalMux I__7515 (
            .O(N__36306),
            .I(N__36297));
    Span4Mux_h I__7514 (
            .O(N__36303),
            .I(N__36292));
    LocalMux I__7513 (
            .O(N__36300),
            .I(N__36292));
    Odrv12 I__7512 (
            .O(N__36297),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    Odrv4 I__7511 (
            .O(N__36292),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    InMux I__7510 (
            .O(N__36287),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__7509 (
            .O(N__36284),
            .I(N__36280));
    CascadeMux I__7508 (
            .O(N__36283),
            .I(N__36277));
    InMux I__7507 (
            .O(N__36280),
            .I(N__36272));
    InMux I__7506 (
            .O(N__36277),
            .I(N__36272));
    LocalMux I__7505 (
            .O(N__36272),
            .I(N__36268));
    InMux I__7504 (
            .O(N__36271),
            .I(N__36265));
    Span4Mux_v I__7503 (
            .O(N__36268),
            .I(N__36262));
    LocalMux I__7502 (
            .O(N__36265),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    Odrv4 I__7501 (
            .O(N__36262),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__7500 (
            .O(N__36257),
            .I(N__36254));
    LocalMux I__7499 (
            .O(N__36254),
            .I(N__36249));
    InMux I__7498 (
            .O(N__36253),
            .I(N__36244));
    InMux I__7497 (
            .O(N__36252),
            .I(N__36244));
    Span4Mux_h I__7496 (
            .O(N__36249),
            .I(N__36239));
    LocalMux I__7495 (
            .O(N__36244),
            .I(N__36239));
    Odrv4 I__7494 (
            .O(N__36239),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__7493 (
            .O(N__36236),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__7492 (
            .O(N__36233),
            .I(N__36230));
    InMux I__7491 (
            .O(N__36230),
            .I(N__36227));
    LocalMux I__7490 (
            .O(N__36227),
            .I(N__36222));
    InMux I__7489 (
            .O(N__36226),
            .I(N__36219));
    InMux I__7488 (
            .O(N__36225),
            .I(N__36216));
    Span4Mux_v I__7487 (
            .O(N__36222),
            .I(N__36211));
    LocalMux I__7486 (
            .O(N__36219),
            .I(N__36211));
    LocalMux I__7485 (
            .O(N__36216),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv4 I__7484 (
            .O(N__36211),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    CascadeMux I__7483 (
            .O(N__36206),
            .I(N__36203));
    InMux I__7482 (
            .O(N__36203),
            .I(N__36200));
    LocalMux I__7481 (
            .O(N__36200),
            .I(N__36195));
    InMux I__7480 (
            .O(N__36199),
            .I(N__36190));
    InMux I__7479 (
            .O(N__36198),
            .I(N__36190));
    Span4Mux_v I__7478 (
            .O(N__36195),
            .I(N__36187));
    LocalMux I__7477 (
            .O(N__36190),
            .I(N__36184));
    Odrv4 I__7476 (
            .O(N__36187),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv12 I__7475 (
            .O(N__36184),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    InMux I__7474 (
            .O(N__36179),
            .I(bfn_16_10_0_));
    CascadeMux I__7473 (
            .O(N__36176),
            .I(N__36173));
    InMux I__7472 (
            .O(N__36173),
            .I(N__36170));
    LocalMux I__7471 (
            .O(N__36170),
            .I(N__36165));
    InMux I__7470 (
            .O(N__36169),
            .I(N__36162));
    InMux I__7469 (
            .O(N__36168),
            .I(N__36159));
    Span4Mux_v I__7468 (
            .O(N__36165),
            .I(N__36154));
    LocalMux I__7467 (
            .O(N__36162),
            .I(N__36154));
    LocalMux I__7466 (
            .O(N__36159),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__7465 (
            .O(N__36154),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__7464 (
            .O(N__36149),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__7463 (
            .O(N__36146),
            .I(N__36139));
    InMux I__7462 (
            .O(N__36145),
            .I(N__36139));
    InMux I__7461 (
            .O(N__36144),
            .I(N__36136));
    LocalMux I__7460 (
            .O(N__36139),
            .I(N__36133));
    LocalMux I__7459 (
            .O(N__36136),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    Odrv4 I__7458 (
            .O(N__36133),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__7457 (
            .O(N__36128),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__7456 (
            .O(N__36125),
            .I(N__36118));
    InMux I__7455 (
            .O(N__36124),
            .I(N__36118));
    InMux I__7454 (
            .O(N__36123),
            .I(N__36115));
    LocalMux I__7453 (
            .O(N__36118),
            .I(N__36112));
    LocalMux I__7452 (
            .O(N__36115),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    Odrv4 I__7451 (
            .O(N__36112),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__7450 (
            .O(N__36107),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__7449 (
            .O(N__36104),
            .I(N__36100));
    InMux I__7448 (
            .O(N__36103),
            .I(N__36096));
    InMux I__7447 (
            .O(N__36100),
            .I(N__36093));
    InMux I__7446 (
            .O(N__36099),
            .I(N__36090));
    LocalMux I__7445 (
            .O(N__36096),
            .I(N__36085));
    LocalMux I__7444 (
            .O(N__36093),
            .I(N__36085));
    LocalMux I__7443 (
            .O(N__36090),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    Odrv4 I__7442 (
            .O(N__36085),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__7441 (
            .O(N__36080),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__7440 (
            .O(N__36077),
            .I(N__36073));
    InMux I__7439 (
            .O(N__36076),
            .I(N__36069));
    InMux I__7438 (
            .O(N__36073),
            .I(N__36066));
    InMux I__7437 (
            .O(N__36072),
            .I(N__36063));
    LocalMux I__7436 (
            .O(N__36069),
            .I(N__36058));
    LocalMux I__7435 (
            .O(N__36066),
            .I(N__36058));
    LocalMux I__7434 (
            .O(N__36063),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    Odrv4 I__7433 (
            .O(N__36058),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__7432 (
            .O(N__36053),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__7431 (
            .O(N__36050),
            .I(N__36046));
    CascadeMux I__7430 (
            .O(N__36049),
            .I(N__36043));
    InMux I__7429 (
            .O(N__36046),
            .I(N__36037));
    InMux I__7428 (
            .O(N__36043),
            .I(N__36037));
    InMux I__7427 (
            .O(N__36042),
            .I(N__36034));
    LocalMux I__7426 (
            .O(N__36037),
            .I(N__36031));
    LocalMux I__7425 (
            .O(N__36034),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    Odrv4 I__7424 (
            .O(N__36031),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__7423 (
            .O(N__36026),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__7422 (
            .O(N__36023),
            .I(N__36019));
    CascadeMux I__7421 (
            .O(N__36022),
            .I(N__36016));
    InMux I__7420 (
            .O(N__36019),
            .I(N__36010));
    InMux I__7419 (
            .O(N__36016),
            .I(N__36010));
    InMux I__7418 (
            .O(N__36015),
            .I(N__36007));
    LocalMux I__7417 (
            .O(N__36010),
            .I(N__36004));
    LocalMux I__7416 (
            .O(N__36007),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    Odrv4 I__7415 (
            .O(N__36004),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__7414 (
            .O(N__35999),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__7413 (
            .O(N__35996),
            .I(N__35993));
    InMux I__7412 (
            .O(N__35993),
            .I(N__35990));
    LocalMux I__7411 (
            .O(N__35990),
            .I(N__35985));
    InMux I__7410 (
            .O(N__35989),
            .I(N__35982));
    InMux I__7409 (
            .O(N__35988),
            .I(N__35979));
    Span4Mux_v I__7408 (
            .O(N__35985),
            .I(N__35976));
    LocalMux I__7407 (
            .O(N__35982),
            .I(N__35973));
    LocalMux I__7406 (
            .O(N__35979),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    Odrv4 I__7405 (
            .O(N__35976),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    Odrv4 I__7404 (
            .O(N__35973),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__7403 (
            .O(N__35966),
            .I(bfn_16_9_0_));
    CascadeMux I__7402 (
            .O(N__35963),
            .I(N__35960));
    InMux I__7401 (
            .O(N__35960),
            .I(N__35957));
    LocalMux I__7400 (
            .O(N__35957),
            .I(N__35952));
    InMux I__7399 (
            .O(N__35956),
            .I(N__35949));
    InMux I__7398 (
            .O(N__35955),
            .I(N__35946));
    Span4Mux_v I__7397 (
            .O(N__35952),
            .I(N__35941));
    LocalMux I__7396 (
            .O(N__35949),
            .I(N__35941));
    LocalMux I__7395 (
            .O(N__35946),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    Odrv4 I__7394 (
            .O(N__35941),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__7393 (
            .O(N__35936),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__7392 (
            .O(N__35933),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_ ));
    InMux I__7391 (
            .O(N__35930),
            .I(N__35927));
    LocalMux I__7390 (
            .O(N__35927),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ));
    CascadeMux I__7389 (
            .O(N__35924),
            .I(N__35920));
    CascadeMux I__7388 (
            .O(N__35923),
            .I(N__35917));
    InMux I__7387 (
            .O(N__35920),
            .I(N__35914));
    InMux I__7386 (
            .O(N__35917),
            .I(N__35910));
    LocalMux I__7385 (
            .O(N__35914),
            .I(N__35907));
    InMux I__7384 (
            .O(N__35913),
            .I(N__35904));
    LocalMux I__7383 (
            .O(N__35910),
            .I(N__35897));
    Span4Mux_v I__7382 (
            .O(N__35907),
            .I(N__35897));
    LocalMux I__7381 (
            .O(N__35904),
            .I(N__35897));
    Odrv4 I__7380 (
            .O(N__35897),
            .I(elapsed_time_ns_1_RNIAE2591_0_2));
    CascadeMux I__7379 (
            .O(N__35894),
            .I(N__35891));
    InMux I__7378 (
            .O(N__35891),
            .I(N__35887));
    InMux I__7377 (
            .O(N__35890),
            .I(N__35883));
    LocalMux I__7376 (
            .O(N__35887),
            .I(N__35880));
    InMux I__7375 (
            .O(N__35886),
            .I(N__35877));
    LocalMux I__7374 (
            .O(N__35883),
            .I(N__35872));
    Span4Mux_v I__7373 (
            .O(N__35880),
            .I(N__35872));
    LocalMux I__7372 (
            .O(N__35877),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    Odrv4 I__7371 (
            .O(N__35872),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__7370 (
            .O(N__35867),
            .I(N__35864));
    LocalMux I__7369 (
            .O(N__35864),
            .I(N__35861));
    Span4Mux_h I__7368 (
            .O(N__35861),
            .I(N__35857));
    InMux I__7367 (
            .O(N__35860),
            .I(N__35854));
    Odrv4 I__7366 (
            .O(N__35857),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    LocalMux I__7365 (
            .O(N__35854),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__7364 (
            .O(N__35849),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__7363 (
            .O(N__35846),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__7362 (
            .O(N__35843),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__7361 (
            .O(N__35840),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__7360 (
            .O(N__35837),
            .I(N__35834));
    LocalMux I__7359 (
            .O(N__35834),
            .I(N__35831));
    Span4Mux_h I__7358 (
            .O(N__35831),
            .I(N__35828));
    Odrv4 I__7357 (
            .O(N__35828),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__7356 (
            .O(N__35825),
            .I(N__35822));
    LocalMux I__7355 (
            .O(N__35822),
            .I(\phase_controller_inst2.start_timer_hc_RNOZ0Z_0 ));
    InMux I__7354 (
            .O(N__35819),
            .I(N__35814));
    InMux I__7353 (
            .O(N__35818),
            .I(N__35811));
    InMux I__7352 (
            .O(N__35817),
            .I(N__35807));
    LocalMux I__7351 (
            .O(N__35814),
            .I(N__35804));
    LocalMux I__7350 (
            .O(N__35811),
            .I(N__35801));
    InMux I__7349 (
            .O(N__35810),
            .I(N__35798));
    LocalMux I__7348 (
            .O(N__35807),
            .I(N__35791));
    Span12Mux_h I__7347 (
            .O(N__35804),
            .I(N__35791));
    Span12Mux_s5_v I__7346 (
            .O(N__35801),
            .I(N__35791));
    LocalMux I__7345 (
            .O(N__35798),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv12 I__7344 (
            .O(N__35791),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    CEMux I__7343 (
            .O(N__35786),
            .I(N__35781));
    CEMux I__7342 (
            .O(N__35785),
            .I(N__35778));
    CEMux I__7341 (
            .O(N__35784),
            .I(N__35774));
    LocalMux I__7340 (
            .O(N__35781),
            .I(N__35771));
    LocalMux I__7339 (
            .O(N__35778),
            .I(N__35768));
    CEMux I__7338 (
            .O(N__35777),
            .I(N__35765));
    LocalMux I__7337 (
            .O(N__35774),
            .I(N__35762));
    Span4Mux_v I__7336 (
            .O(N__35771),
            .I(N__35757));
    Span4Mux_v I__7335 (
            .O(N__35768),
            .I(N__35757));
    LocalMux I__7334 (
            .O(N__35765),
            .I(N__35754));
    Span4Mux_v I__7333 (
            .O(N__35762),
            .I(N__35747));
    Span4Mux_h I__7332 (
            .O(N__35757),
            .I(N__35747));
    Span4Mux_v I__7331 (
            .O(N__35754),
            .I(N__35747));
    Odrv4 I__7330 (
            .O(N__35747),
            .I(\delay_measurement_inst.delay_tr_timer.N_435_i ));
    InMux I__7329 (
            .O(N__35744),
            .I(N__35738));
    InMux I__7328 (
            .O(N__35743),
            .I(N__35733));
    InMux I__7327 (
            .O(N__35742),
            .I(N__35733));
    InMux I__7326 (
            .O(N__35741),
            .I(N__35730));
    LocalMux I__7325 (
            .O(N__35738),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__7324 (
            .O(N__35733),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__7323 (
            .O(N__35730),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__7322 (
            .O(N__35723),
            .I(N__35709));
    InMux I__7321 (
            .O(N__35722),
            .I(N__35709));
    InMux I__7320 (
            .O(N__35721),
            .I(N__35700));
    InMux I__7319 (
            .O(N__35720),
            .I(N__35700));
    InMux I__7318 (
            .O(N__35719),
            .I(N__35700));
    InMux I__7317 (
            .O(N__35718),
            .I(N__35700));
    InMux I__7316 (
            .O(N__35717),
            .I(N__35687));
    InMux I__7315 (
            .O(N__35716),
            .I(N__35687));
    InMux I__7314 (
            .O(N__35715),
            .I(N__35687));
    InMux I__7313 (
            .O(N__35714),
            .I(N__35687));
    LocalMux I__7312 (
            .O(N__35709),
            .I(N__35666));
    LocalMux I__7311 (
            .O(N__35700),
            .I(N__35666));
    InMux I__7310 (
            .O(N__35699),
            .I(N__35657));
    InMux I__7309 (
            .O(N__35698),
            .I(N__35657));
    InMux I__7308 (
            .O(N__35697),
            .I(N__35657));
    InMux I__7307 (
            .O(N__35696),
            .I(N__35657));
    LocalMux I__7306 (
            .O(N__35687),
            .I(N__35654));
    InMux I__7305 (
            .O(N__35686),
            .I(N__35645));
    InMux I__7304 (
            .O(N__35685),
            .I(N__35645));
    InMux I__7303 (
            .O(N__35684),
            .I(N__35645));
    InMux I__7302 (
            .O(N__35683),
            .I(N__35645));
    InMux I__7301 (
            .O(N__35682),
            .I(N__35636));
    InMux I__7300 (
            .O(N__35681),
            .I(N__35636));
    InMux I__7299 (
            .O(N__35680),
            .I(N__35636));
    InMux I__7298 (
            .O(N__35679),
            .I(N__35636));
    InMux I__7297 (
            .O(N__35678),
            .I(N__35627));
    InMux I__7296 (
            .O(N__35677),
            .I(N__35627));
    InMux I__7295 (
            .O(N__35676),
            .I(N__35627));
    InMux I__7294 (
            .O(N__35675),
            .I(N__35627));
    InMux I__7293 (
            .O(N__35674),
            .I(N__35618));
    InMux I__7292 (
            .O(N__35673),
            .I(N__35618));
    InMux I__7291 (
            .O(N__35672),
            .I(N__35618));
    InMux I__7290 (
            .O(N__35671),
            .I(N__35618));
    Span4Mux_h I__7289 (
            .O(N__35666),
            .I(N__35615));
    LocalMux I__7288 (
            .O(N__35657),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__7287 (
            .O(N__35654),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__7286 (
            .O(N__35645),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__7285 (
            .O(N__35636),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__7284 (
            .O(N__35627),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__7283 (
            .O(N__35618),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__7282 (
            .O(N__35615),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__7281 (
            .O(N__35600),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__7280 (
            .O(N__35597),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__7279 (
            .O(N__35594),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__7278 (
            .O(N__35591),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__7277 (
            .O(N__35588),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__7276 (
            .O(N__35585),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__7275 (
            .O(N__35582),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__7274 (
            .O(N__35579),
            .I(bfn_15_23_0_));
    InMux I__7273 (
            .O(N__35576),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    CascadeMux I__7272 (
            .O(N__35573),
            .I(N__35569));
    InMux I__7271 (
            .O(N__35572),
            .I(N__35565));
    InMux I__7270 (
            .O(N__35569),
            .I(N__35562));
    InMux I__7269 (
            .O(N__35568),
            .I(N__35559));
    LocalMux I__7268 (
            .O(N__35565),
            .I(N__35556));
    LocalMux I__7267 (
            .O(N__35562),
            .I(N__35551));
    LocalMux I__7266 (
            .O(N__35559),
            .I(N__35551));
    Span4Mux_v I__7265 (
            .O(N__35556),
            .I(N__35547));
    Span4Mux_v I__7264 (
            .O(N__35551),
            .I(N__35544));
    InMux I__7263 (
            .O(N__35550),
            .I(N__35541));
    Odrv4 I__7262 (
            .O(N__35547),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__7261 (
            .O(N__35544),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__7260 (
            .O(N__35541),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__7259 (
            .O(N__35534),
            .I(bfn_15_21_0_));
    InMux I__7258 (
            .O(N__35531),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__7257 (
            .O(N__35528),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__7256 (
            .O(N__35525),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__7255 (
            .O(N__35522),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__7254 (
            .O(N__35519),
            .I(N__35516));
    LocalMux I__7253 (
            .O(N__35516),
            .I(N__35512));
    InMux I__7252 (
            .O(N__35515),
            .I(N__35509));
    Span4Mux_h I__7251 (
            .O(N__35512),
            .I(N__35503));
    LocalMux I__7250 (
            .O(N__35509),
            .I(N__35503));
    InMux I__7249 (
            .O(N__35508),
            .I(N__35500));
    Span4Mux_v I__7248 (
            .O(N__35503),
            .I(N__35496));
    LocalMux I__7247 (
            .O(N__35500),
            .I(N__35493));
    InMux I__7246 (
            .O(N__35499),
            .I(N__35490));
    Odrv4 I__7245 (
            .O(N__35496),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__7244 (
            .O(N__35493),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__7243 (
            .O(N__35490),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__7242 (
            .O(N__35483),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__7241 (
            .O(N__35480),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__7240 (
            .O(N__35477),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__7239 (
            .O(N__35474),
            .I(N__35467));
    InMux I__7238 (
            .O(N__35473),
            .I(N__35467));
    CascadeMux I__7237 (
            .O(N__35472),
            .I(N__35464));
    LocalMux I__7236 (
            .O(N__35467),
            .I(N__35461));
    InMux I__7235 (
            .O(N__35464),
            .I(N__35458));
    Span4Mux_h I__7234 (
            .O(N__35461),
            .I(N__35452));
    LocalMux I__7233 (
            .O(N__35458),
            .I(N__35452));
    InMux I__7232 (
            .O(N__35457),
            .I(N__35449));
    Odrv4 I__7231 (
            .O(N__35452),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__7230 (
            .O(N__35449),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__7229 (
            .O(N__35444),
            .I(bfn_15_22_0_));
    CascadeMux I__7228 (
            .O(N__35441),
            .I(N__35438));
    InMux I__7227 (
            .O(N__35438),
            .I(N__35431));
    InMux I__7226 (
            .O(N__35437),
            .I(N__35431));
    InMux I__7225 (
            .O(N__35436),
            .I(N__35428));
    LocalMux I__7224 (
            .O(N__35431),
            .I(N__35424));
    LocalMux I__7223 (
            .O(N__35428),
            .I(N__35421));
    InMux I__7222 (
            .O(N__35427),
            .I(N__35418));
    Span4Mux_v I__7221 (
            .O(N__35424),
            .I(N__35415));
    Span4Mux_h I__7220 (
            .O(N__35421),
            .I(N__35412));
    LocalMux I__7219 (
            .O(N__35418),
            .I(N__35409));
    Odrv4 I__7218 (
            .O(N__35415),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__7217 (
            .O(N__35412),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__7216 (
            .O(N__35409),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__7215 (
            .O(N__35402),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__7214 (
            .O(N__35399),
            .I(N__35396));
    InMux I__7213 (
            .O(N__35396),
            .I(N__35392));
    CascadeMux I__7212 (
            .O(N__35395),
            .I(N__35389));
    LocalMux I__7211 (
            .O(N__35392),
            .I(N__35386));
    InMux I__7210 (
            .O(N__35389),
            .I(N__35383));
    Span4Mux_v I__7209 (
            .O(N__35386),
            .I(N__35376));
    LocalMux I__7208 (
            .O(N__35383),
            .I(N__35376));
    InMux I__7207 (
            .O(N__35382),
            .I(N__35373));
    InMux I__7206 (
            .O(N__35381),
            .I(N__35370));
    Span4Mux_h I__7205 (
            .O(N__35376),
            .I(N__35365));
    LocalMux I__7204 (
            .O(N__35373),
            .I(N__35365));
    LocalMux I__7203 (
            .O(N__35370),
            .I(N__35362));
    Span4Mux_v I__7202 (
            .O(N__35365),
            .I(N__35359));
    Span4Mux_h I__7201 (
            .O(N__35362),
            .I(N__35356));
    Odrv4 I__7200 (
            .O(N__35359),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__7199 (
            .O(N__35356),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__7198 (
            .O(N__35351),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__7197 (
            .O(N__35348),
            .I(N__35345));
    InMux I__7196 (
            .O(N__35345),
            .I(N__35341));
    CascadeMux I__7195 (
            .O(N__35344),
            .I(N__35338));
    LocalMux I__7194 (
            .O(N__35341),
            .I(N__35333));
    InMux I__7193 (
            .O(N__35338),
            .I(N__35328));
    InMux I__7192 (
            .O(N__35337),
            .I(N__35328));
    InMux I__7191 (
            .O(N__35336),
            .I(N__35325));
    Span4Mux_v I__7190 (
            .O(N__35333),
            .I(N__35320));
    LocalMux I__7189 (
            .O(N__35328),
            .I(N__35320));
    LocalMux I__7188 (
            .O(N__35325),
            .I(N__35317));
    Span4Mux_v I__7187 (
            .O(N__35320),
            .I(N__35314));
    Span4Mux_h I__7186 (
            .O(N__35317),
            .I(N__35311));
    Odrv4 I__7185 (
            .O(N__35314),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__7184 (
            .O(N__35311),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__7183 (
            .O(N__35306),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__7182 (
            .O(N__35303),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__7181 (
            .O(N__35300),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__7180 (
            .O(N__35297),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__7179 (
            .O(N__35294),
            .I(N__35290));
    InMux I__7178 (
            .O(N__35293),
            .I(N__35287));
    InMux I__7177 (
            .O(N__35290),
            .I(N__35284));
    LocalMux I__7176 (
            .O(N__35287),
            .I(N__35279));
    LocalMux I__7175 (
            .O(N__35284),
            .I(N__35279));
    Span4Mux_v I__7174 (
            .O(N__35279),
            .I(N__35275));
    InMux I__7173 (
            .O(N__35278),
            .I(N__35271));
    Span4Mux_v I__7172 (
            .O(N__35275),
            .I(N__35268));
    InMux I__7171 (
            .O(N__35274),
            .I(N__35265));
    LocalMux I__7170 (
            .O(N__35271),
            .I(N__35262));
    Odrv4 I__7169 (
            .O(N__35268),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__7168 (
            .O(N__35265),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    Odrv4 I__7167 (
            .O(N__35262),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__7166 (
            .O(N__35255),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__7165 (
            .O(N__35252),
            .I(N__35249));
    LocalMux I__7164 (
            .O(N__35249),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__7163 (
            .O(N__35246),
            .I(N__35241));
    InMux I__7162 (
            .O(N__35245),
            .I(N__35238));
    CascadeMux I__7161 (
            .O(N__35244),
            .I(N__35235));
    LocalMux I__7160 (
            .O(N__35241),
            .I(N__35232));
    LocalMux I__7159 (
            .O(N__35238),
            .I(N__35229));
    InMux I__7158 (
            .O(N__35235),
            .I(N__35226));
    Odrv4 I__7157 (
            .O(N__35232),
            .I(\current_shift_inst.un4_control_input1_10 ));
    Odrv12 I__7156 (
            .O(N__35229),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__7155 (
            .O(N__35226),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__7154 (
            .O(N__35219),
            .I(N__35216));
    LocalMux I__7153 (
            .O(N__35216),
            .I(N__35213));
    Odrv4 I__7152 (
            .O(N__35213),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    InMux I__7151 (
            .O(N__35210),
            .I(N__35207));
    LocalMux I__7150 (
            .O(N__35207),
            .I(N__35204));
    Odrv4 I__7149 (
            .O(N__35204),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    CascadeMux I__7148 (
            .O(N__35201),
            .I(N__35197));
    CascadeMux I__7147 (
            .O(N__35200),
            .I(N__35194));
    InMux I__7146 (
            .O(N__35197),
            .I(N__35188));
    InMux I__7145 (
            .O(N__35194),
            .I(N__35188));
    InMux I__7144 (
            .O(N__35193),
            .I(N__35185));
    LocalMux I__7143 (
            .O(N__35188),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__7142 (
            .O(N__35185),
            .I(\current_shift_inst.un4_control_input1_19 ));
    InMux I__7141 (
            .O(N__35180),
            .I(N__35177));
    LocalMux I__7140 (
            .O(N__35177),
            .I(N__35174));
    Odrv4 I__7139 (
            .O(N__35174),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__7138 (
            .O(N__35171),
            .I(N__35168));
    LocalMux I__7137 (
            .O(N__35168),
            .I(N__35165));
    Span4Mux_h I__7136 (
            .O(N__35165),
            .I(N__35162));
    Odrv4 I__7135 (
            .O(N__35162),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__7134 (
            .O(N__35159),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__7133 (
            .O(N__35156),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__7132 (
            .O(N__35153),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__7131 (
            .O(N__35150),
            .I(N__35147));
    LocalMux I__7130 (
            .O(N__35147),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    CascadeMux I__7129 (
            .O(N__35144),
            .I(N__35141));
    InMux I__7128 (
            .O(N__35141),
            .I(N__35138));
    LocalMux I__7127 (
            .O(N__35138),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__7126 (
            .O(N__35135),
            .I(N__35131));
    InMux I__7125 (
            .O(N__35134),
            .I(N__35128));
    LocalMux I__7124 (
            .O(N__35131),
            .I(N__35122));
    LocalMux I__7123 (
            .O(N__35128),
            .I(N__35122));
    InMux I__7122 (
            .O(N__35127),
            .I(N__35119));
    Odrv12 I__7121 (
            .O(N__35122),
            .I(\current_shift_inst.un4_control_input1_16 ));
    LocalMux I__7120 (
            .O(N__35119),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__7119 (
            .O(N__35114),
            .I(N__35110));
    InMux I__7118 (
            .O(N__35113),
            .I(N__35107));
    LocalMux I__7117 (
            .O(N__35110),
            .I(N__35103));
    LocalMux I__7116 (
            .O(N__35107),
            .I(N__35100));
    InMux I__7115 (
            .O(N__35106),
            .I(N__35097));
    Odrv4 I__7114 (
            .O(N__35103),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv4 I__7113 (
            .O(N__35100),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__7112 (
            .O(N__35097),
            .I(\current_shift_inst.un4_control_input1_11 ));
    CascadeMux I__7111 (
            .O(N__35090),
            .I(N__35087));
    InMux I__7110 (
            .O(N__35087),
            .I(N__35084));
    LocalMux I__7109 (
            .O(N__35084),
            .I(N__35081));
    Span12Mux_v I__7108 (
            .O(N__35081),
            .I(N__35078));
    Odrv12 I__7107 (
            .O(N__35078),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    InMux I__7106 (
            .O(N__35075),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__7105 (
            .O(N__35072),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    CascadeMux I__7104 (
            .O(N__35069),
            .I(N__35066));
    InMux I__7103 (
            .O(N__35066),
            .I(N__35063));
    LocalMux I__7102 (
            .O(N__35063),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    InMux I__7101 (
            .O(N__35060),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__7100 (
            .O(N__35057),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__7099 (
            .O(N__35054),
            .I(bfn_15_17_0_));
    InMux I__7098 (
            .O(N__35051),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    CascadeMux I__7097 (
            .O(N__35048),
            .I(N__35045));
    InMux I__7096 (
            .O(N__35045),
            .I(N__35042));
    LocalMux I__7095 (
            .O(N__35042),
            .I(N__35039));
    Span4Mux_v I__7094 (
            .O(N__35039),
            .I(N__35036));
    Odrv4 I__7093 (
            .O(N__35036),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    InMux I__7092 (
            .O(N__35033),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__7091 (
            .O(N__35030),
            .I(N__35027));
    LocalMux I__7090 (
            .O(N__35027),
            .I(N__35024));
    Span4Mux_h I__7089 (
            .O(N__35024),
            .I(N__35021));
    Odrv4 I__7088 (
            .O(N__35021),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    InMux I__7087 (
            .O(N__35018),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__7086 (
            .O(N__35015),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    CascadeMux I__7085 (
            .O(N__35012),
            .I(N__35009));
    InMux I__7084 (
            .O(N__35009),
            .I(N__35006));
    LocalMux I__7083 (
            .O(N__35006),
            .I(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ));
    InMux I__7082 (
            .O(N__35003),
            .I(N__35000));
    LocalMux I__7081 (
            .O(N__35000),
            .I(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ));
    CascadeMux I__7080 (
            .O(N__34997),
            .I(N__34994));
    InMux I__7079 (
            .O(N__34994),
            .I(N__34991));
    LocalMux I__7078 (
            .O(N__34991),
            .I(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ));
    InMux I__7077 (
            .O(N__34988),
            .I(N__34985));
    LocalMux I__7076 (
            .O(N__34985),
            .I(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ));
    CascadeMux I__7075 (
            .O(N__34982),
            .I(N__34979));
    InMux I__7074 (
            .O(N__34979),
            .I(N__34976));
    LocalMux I__7073 (
            .O(N__34976),
            .I(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ));
    InMux I__7072 (
            .O(N__34973),
            .I(N__34970));
    LocalMux I__7071 (
            .O(N__34970),
            .I(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ));
    CascadeMux I__7070 (
            .O(N__34967),
            .I(N__34964));
    InMux I__7069 (
            .O(N__34964),
            .I(N__34961));
    LocalMux I__7068 (
            .O(N__34961),
            .I(N__34958));
    Span4Mux_v I__7067 (
            .O(N__34958),
            .I(N__34955));
    Odrv4 I__7066 (
            .O(N__34955),
            .I(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ));
    InMux I__7065 (
            .O(N__34952),
            .I(N__34949));
    LocalMux I__7064 (
            .O(N__34949),
            .I(N__34946));
    Span4Mux_h I__7063 (
            .O(N__34946),
            .I(N__34943));
    Odrv4 I__7062 (
            .O(N__34943),
            .I(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ));
    InMux I__7061 (
            .O(N__34940),
            .I(N__34937));
    LocalMux I__7060 (
            .O(N__34937),
            .I(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ));
    CascadeMux I__7059 (
            .O(N__34934),
            .I(N__34931));
    InMux I__7058 (
            .O(N__34931),
            .I(N__34928));
    LocalMux I__7057 (
            .O(N__34928),
            .I(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ));
    InMux I__7056 (
            .O(N__34925),
            .I(N__34922));
    LocalMux I__7055 (
            .O(N__34922),
            .I(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ));
    CascadeMux I__7054 (
            .O(N__34919),
            .I(N__34916));
    InMux I__7053 (
            .O(N__34916),
            .I(N__34913));
    LocalMux I__7052 (
            .O(N__34913),
            .I(N__34910));
    Span12Mux_v I__7051 (
            .O(N__34910),
            .I(N__34907));
    Odrv12 I__7050 (
            .O(N__34907),
            .I(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ));
    InMux I__7049 (
            .O(N__34904),
            .I(N__34901));
    LocalMux I__7048 (
            .O(N__34901),
            .I(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ));
    CascadeMux I__7047 (
            .O(N__34898),
            .I(N__34895));
    InMux I__7046 (
            .O(N__34895),
            .I(N__34892));
    LocalMux I__7045 (
            .O(N__34892),
            .I(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ));
    InMux I__7044 (
            .O(N__34889),
            .I(N__34886));
    LocalMux I__7043 (
            .O(N__34886),
            .I(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ));
    CascadeMux I__7042 (
            .O(N__34883),
            .I(N__34880));
    InMux I__7041 (
            .O(N__34880),
            .I(N__34877));
    LocalMux I__7040 (
            .O(N__34877),
            .I(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ));
    InMux I__7039 (
            .O(N__34874),
            .I(N__34871));
    LocalMux I__7038 (
            .O(N__34871),
            .I(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ));
    InMux I__7037 (
            .O(N__34868),
            .I(N__34865));
    LocalMux I__7036 (
            .O(N__34865),
            .I(N__34862));
    Span4Mux_v I__7035 (
            .O(N__34862),
            .I(N__34859));
    Odrv4 I__7034 (
            .O(N__34859),
            .I(\phase_controller_inst1.stoper_tr.un6_running_17 ));
    InMux I__7033 (
            .O(N__34856),
            .I(N__34852));
    InMux I__7032 (
            .O(N__34855),
            .I(N__34849));
    LocalMux I__7031 (
            .O(N__34852),
            .I(N__34846));
    LocalMux I__7030 (
            .O(N__34849),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__7029 (
            .O(N__34846),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    CascadeMux I__7028 (
            .O(N__34841),
            .I(N__34838));
    InMux I__7027 (
            .O(N__34838),
            .I(N__34835));
    LocalMux I__7026 (
            .O(N__34835),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ));
    CascadeMux I__7025 (
            .O(N__34832),
            .I(N__34829));
    InMux I__7024 (
            .O(N__34829),
            .I(N__34826));
    LocalMux I__7023 (
            .O(N__34826),
            .I(N__34823));
    Odrv12 I__7022 (
            .O(N__34823),
            .I(\phase_controller_inst1.stoper_tr.un6_running_18 ));
    InMux I__7021 (
            .O(N__34820),
            .I(N__34816));
    InMux I__7020 (
            .O(N__34819),
            .I(N__34813));
    LocalMux I__7019 (
            .O(N__34816),
            .I(N__34810));
    LocalMux I__7018 (
            .O(N__34813),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__7017 (
            .O(N__34810),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__7016 (
            .O(N__34805),
            .I(N__34802));
    LocalMux I__7015 (
            .O(N__34802),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ));
    InMux I__7014 (
            .O(N__34799),
            .I(N__34795));
    InMux I__7013 (
            .O(N__34798),
            .I(N__34792));
    LocalMux I__7012 (
            .O(N__34795),
            .I(N__34789));
    LocalMux I__7011 (
            .O(N__34792),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__7010 (
            .O(N__34789),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    CascadeMux I__7009 (
            .O(N__34784),
            .I(N__34781));
    InMux I__7008 (
            .O(N__34781),
            .I(N__34778));
    LocalMux I__7007 (
            .O(N__34778),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ));
    InMux I__7006 (
            .O(N__34775),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_19 ));
    InMux I__7005 (
            .O(N__34772),
            .I(N__34768));
    InMux I__7004 (
            .O(N__34771),
            .I(N__34764));
    LocalMux I__7003 (
            .O(N__34768),
            .I(N__34761));
    InMux I__7002 (
            .O(N__34767),
            .I(N__34758));
    LocalMux I__7001 (
            .O(N__34764),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO ));
    Odrv4 I__7000 (
            .O(N__34761),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO ));
    LocalMux I__6999 (
            .O(N__34758),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO ));
    InMux I__6998 (
            .O(N__34751),
            .I(N__34748));
    LocalMux I__6997 (
            .O(N__34748),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    CascadeMux I__6996 (
            .O(N__34745),
            .I(N__34742));
    InMux I__6995 (
            .O(N__34742),
            .I(N__34739));
    LocalMux I__6994 (
            .O(N__34739),
            .I(N__34736));
    Span4Mux_h I__6993 (
            .O(N__34736),
            .I(N__34733));
    Odrv4 I__6992 (
            .O(N__34733),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    CascadeMux I__6991 (
            .O(N__34730),
            .I(N__34727));
    InMux I__6990 (
            .O(N__34727),
            .I(N__34724));
    LocalMux I__6989 (
            .O(N__34724),
            .I(N__34721));
    Odrv4 I__6988 (
            .O(N__34721),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    InMux I__6987 (
            .O(N__34718),
            .I(N__34715));
    LocalMux I__6986 (
            .O(N__34715),
            .I(N__34712));
    Odrv12 I__6985 (
            .O(N__34712),
            .I(\phase_controller_inst1.stoper_tr.un6_running_10 ));
    InMux I__6984 (
            .O(N__34709),
            .I(N__34705));
    InMux I__6983 (
            .O(N__34708),
            .I(N__34702));
    LocalMux I__6982 (
            .O(N__34705),
            .I(N__34699));
    LocalMux I__6981 (
            .O(N__34702),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__6980 (
            .O(N__34699),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    CascadeMux I__6979 (
            .O(N__34694),
            .I(N__34691));
    InMux I__6978 (
            .O(N__34691),
            .I(N__34688));
    LocalMux I__6977 (
            .O(N__34688),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__6976 (
            .O(N__34685),
            .I(N__34682));
    LocalMux I__6975 (
            .O(N__34682),
            .I(N__34679));
    Odrv4 I__6974 (
            .O(N__34679),
            .I(\phase_controller_inst1.stoper_tr.un6_running_11 ));
    InMux I__6973 (
            .O(N__34676),
            .I(N__34672));
    InMux I__6972 (
            .O(N__34675),
            .I(N__34669));
    LocalMux I__6971 (
            .O(N__34672),
            .I(N__34664));
    LocalMux I__6970 (
            .O(N__34669),
            .I(N__34664));
    Odrv4 I__6969 (
            .O(N__34664),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    CascadeMux I__6968 (
            .O(N__34661),
            .I(N__34658));
    InMux I__6967 (
            .O(N__34658),
            .I(N__34655));
    LocalMux I__6966 (
            .O(N__34655),
            .I(N__34652));
    Odrv4 I__6965 (
            .O(N__34652),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__6964 (
            .O(N__34649),
            .I(N__34646));
    InMux I__6963 (
            .O(N__34646),
            .I(N__34643));
    LocalMux I__6962 (
            .O(N__34643),
            .I(N__34640));
    Sp12to4 I__6961 (
            .O(N__34640),
            .I(N__34637));
    Odrv12 I__6960 (
            .O(N__34637),
            .I(\phase_controller_inst1.stoper_tr.un6_running_12 ));
    InMux I__6959 (
            .O(N__34634),
            .I(N__34630));
    InMux I__6958 (
            .O(N__34633),
            .I(N__34627));
    LocalMux I__6957 (
            .O(N__34630),
            .I(N__34622));
    LocalMux I__6956 (
            .O(N__34627),
            .I(N__34622));
    Odrv4 I__6955 (
            .O(N__34622),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__6954 (
            .O(N__34619),
            .I(N__34616));
    LocalMux I__6953 (
            .O(N__34616),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__6952 (
            .O(N__34613),
            .I(N__34609));
    InMux I__6951 (
            .O(N__34612),
            .I(N__34606));
    LocalMux I__6950 (
            .O(N__34609),
            .I(N__34603));
    LocalMux I__6949 (
            .O(N__34606),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__6948 (
            .O(N__34603),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    CascadeMux I__6947 (
            .O(N__34598),
            .I(N__34595));
    InMux I__6946 (
            .O(N__34595),
            .I(N__34592));
    LocalMux I__6945 (
            .O(N__34592),
            .I(N__34589));
    Odrv4 I__6944 (
            .O(N__34589),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    InMux I__6943 (
            .O(N__34586),
            .I(N__34582));
    InMux I__6942 (
            .O(N__34585),
            .I(N__34579));
    LocalMux I__6941 (
            .O(N__34582),
            .I(N__34576));
    LocalMux I__6940 (
            .O(N__34579),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__6939 (
            .O(N__34576),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__6938 (
            .O(N__34571),
            .I(N__34568));
    InMux I__6937 (
            .O(N__34568),
            .I(N__34565));
    LocalMux I__6936 (
            .O(N__34565),
            .I(N__34562));
    Odrv4 I__6935 (
            .O(N__34562),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    InMux I__6934 (
            .O(N__34559),
            .I(N__34555));
    InMux I__6933 (
            .O(N__34558),
            .I(N__34552));
    LocalMux I__6932 (
            .O(N__34555),
            .I(N__34549));
    LocalMux I__6931 (
            .O(N__34552),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__6930 (
            .O(N__34549),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__6929 (
            .O(N__34544),
            .I(N__34541));
    LocalMux I__6928 (
            .O(N__34541),
            .I(N__34538));
    Span4Mux_v I__6927 (
            .O(N__34538),
            .I(N__34535));
    Odrv4 I__6926 (
            .O(N__34535),
            .I(\phase_controller_inst1.stoper_tr.un6_running_15 ));
    CascadeMux I__6925 (
            .O(N__34532),
            .I(N__34529));
    InMux I__6924 (
            .O(N__34529),
            .I(N__34526));
    LocalMux I__6923 (
            .O(N__34526),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__6922 (
            .O(N__34523),
            .I(N__34519));
    InMux I__6921 (
            .O(N__34522),
            .I(N__34516));
    LocalMux I__6920 (
            .O(N__34519),
            .I(N__34513));
    LocalMux I__6919 (
            .O(N__34516),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__6918 (
            .O(N__34513),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__6917 (
            .O(N__34508),
            .I(N__34505));
    LocalMux I__6916 (
            .O(N__34505),
            .I(N__34502));
    Span4Mux_v I__6915 (
            .O(N__34502),
            .I(N__34499));
    Odrv4 I__6914 (
            .O(N__34499),
            .I(\phase_controller_inst1.stoper_tr.un6_running_16 ));
    CascadeMux I__6913 (
            .O(N__34496),
            .I(N__34493));
    InMux I__6912 (
            .O(N__34493),
            .I(N__34490));
    LocalMux I__6911 (
            .O(N__34490),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ));
    CascadeMux I__6910 (
            .O(N__34487),
            .I(N__34484));
    InMux I__6909 (
            .O(N__34484),
            .I(N__34481));
    LocalMux I__6908 (
            .O(N__34481),
            .I(N__34478));
    Odrv4 I__6907 (
            .O(N__34478),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__6906 (
            .O(N__34475),
            .I(N__34472));
    LocalMux I__6905 (
            .O(N__34472),
            .I(N__34469));
    Span4Mux_v I__6904 (
            .O(N__34469),
            .I(N__34466));
    Odrv4 I__6903 (
            .O(N__34466),
            .I(\phase_controller_inst1.stoper_tr.un6_running_3 ));
    InMux I__6902 (
            .O(N__34463),
            .I(N__34459));
    InMux I__6901 (
            .O(N__34462),
            .I(N__34456));
    LocalMux I__6900 (
            .O(N__34459),
            .I(N__34451));
    LocalMux I__6899 (
            .O(N__34456),
            .I(N__34451));
    Odrv4 I__6898 (
            .O(N__34451),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__6897 (
            .O(N__34448),
            .I(N__34445));
    InMux I__6896 (
            .O(N__34445),
            .I(N__34442));
    LocalMux I__6895 (
            .O(N__34442),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__6894 (
            .O(N__34439),
            .I(N__34436));
    LocalMux I__6893 (
            .O(N__34436),
            .I(N__34433));
    Span4Mux_v I__6892 (
            .O(N__34433),
            .I(N__34430));
    Odrv4 I__6891 (
            .O(N__34430),
            .I(\phase_controller_inst1.stoper_tr.un6_running_4 ));
    InMux I__6890 (
            .O(N__34427),
            .I(N__34423));
    InMux I__6889 (
            .O(N__34426),
            .I(N__34420));
    LocalMux I__6888 (
            .O(N__34423),
            .I(N__34417));
    LocalMux I__6887 (
            .O(N__34420),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__6886 (
            .O(N__34417),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    CascadeMux I__6885 (
            .O(N__34412),
            .I(N__34409));
    InMux I__6884 (
            .O(N__34409),
            .I(N__34406));
    LocalMux I__6883 (
            .O(N__34406),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__6882 (
            .O(N__34403),
            .I(N__34399));
    InMux I__6881 (
            .O(N__34402),
            .I(N__34396));
    LocalMux I__6880 (
            .O(N__34399),
            .I(N__34391));
    LocalMux I__6879 (
            .O(N__34396),
            .I(N__34391));
    Odrv4 I__6878 (
            .O(N__34391),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__6877 (
            .O(N__34388),
            .I(N__34385));
    LocalMux I__6876 (
            .O(N__34385),
            .I(N__34382));
    Span4Mux_v I__6875 (
            .O(N__34382),
            .I(N__34379));
    Odrv4 I__6874 (
            .O(N__34379),
            .I(\phase_controller_inst1.stoper_tr.un6_running_5 ));
    CascadeMux I__6873 (
            .O(N__34376),
            .I(N__34373));
    InMux I__6872 (
            .O(N__34373),
            .I(N__34370));
    LocalMux I__6871 (
            .O(N__34370),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__6870 (
            .O(N__34367),
            .I(N__34363));
    InMux I__6869 (
            .O(N__34366),
            .I(N__34360));
    LocalMux I__6868 (
            .O(N__34363),
            .I(N__34357));
    LocalMux I__6867 (
            .O(N__34360),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__6866 (
            .O(N__34357),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__6865 (
            .O(N__34352),
            .I(N__34349));
    LocalMux I__6864 (
            .O(N__34349),
            .I(N__34346));
    Span4Mux_v I__6863 (
            .O(N__34346),
            .I(N__34343));
    Odrv4 I__6862 (
            .O(N__34343),
            .I(\phase_controller_inst1.stoper_tr.un6_running_6 ));
    CascadeMux I__6861 (
            .O(N__34340),
            .I(N__34337));
    InMux I__6860 (
            .O(N__34337),
            .I(N__34334));
    LocalMux I__6859 (
            .O(N__34334),
            .I(N__34331));
    Odrv4 I__6858 (
            .O(N__34331),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    InMux I__6857 (
            .O(N__34328),
            .I(N__34325));
    LocalMux I__6856 (
            .O(N__34325),
            .I(N__34322));
    Odrv4 I__6855 (
            .O(N__34322),
            .I(\phase_controller_inst1.stoper_tr.un6_running_7 ));
    InMux I__6854 (
            .O(N__34319),
            .I(N__34315));
    InMux I__6853 (
            .O(N__34318),
            .I(N__34312));
    LocalMux I__6852 (
            .O(N__34315),
            .I(N__34309));
    LocalMux I__6851 (
            .O(N__34312),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv12 I__6850 (
            .O(N__34309),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    CascadeMux I__6849 (
            .O(N__34304),
            .I(N__34301));
    InMux I__6848 (
            .O(N__34301),
            .I(N__34298));
    LocalMux I__6847 (
            .O(N__34298),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__6846 (
            .O(N__34295),
            .I(N__34291));
    InMux I__6845 (
            .O(N__34294),
            .I(N__34288));
    LocalMux I__6844 (
            .O(N__34291),
            .I(N__34283));
    LocalMux I__6843 (
            .O(N__34288),
            .I(N__34283));
    Odrv4 I__6842 (
            .O(N__34283),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__6841 (
            .O(N__34280),
            .I(N__34277));
    LocalMux I__6840 (
            .O(N__34277),
            .I(N__34274));
    Odrv12 I__6839 (
            .O(N__34274),
            .I(\phase_controller_inst1.stoper_tr.un6_running_8 ));
    CascadeMux I__6838 (
            .O(N__34271),
            .I(N__34268));
    InMux I__6837 (
            .O(N__34268),
            .I(N__34265));
    LocalMux I__6836 (
            .O(N__34265),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__6835 (
            .O(N__34262),
            .I(N__34259));
    LocalMux I__6834 (
            .O(N__34259),
            .I(N__34256));
    Span4Mux_v I__6833 (
            .O(N__34256),
            .I(N__34253));
    Odrv4 I__6832 (
            .O(N__34253),
            .I(\phase_controller_inst1.stoper_tr.un6_running_9 ));
    InMux I__6831 (
            .O(N__34250),
            .I(N__34246));
    InMux I__6830 (
            .O(N__34249),
            .I(N__34243));
    LocalMux I__6829 (
            .O(N__34246),
            .I(N__34240));
    LocalMux I__6828 (
            .O(N__34243),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__6827 (
            .O(N__34240),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    CascadeMux I__6826 (
            .O(N__34235),
            .I(N__34232));
    InMux I__6825 (
            .O(N__34232),
            .I(N__34229));
    LocalMux I__6824 (
            .O(N__34229),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__6823 (
            .O(N__34226),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14_cascade_ ));
    InMux I__6822 (
            .O(N__34223),
            .I(N__34217));
    InMux I__6821 (
            .O(N__34222),
            .I(N__34214));
    InMux I__6820 (
            .O(N__34221),
            .I(N__34211));
    InMux I__6819 (
            .O(N__34220),
            .I(N__34208));
    LocalMux I__6818 (
            .O(N__34217),
            .I(\phase_controller_inst1.stoper_tr.N_214 ));
    LocalMux I__6817 (
            .O(N__34214),
            .I(\phase_controller_inst1.stoper_tr.N_214 ));
    LocalMux I__6816 (
            .O(N__34211),
            .I(\phase_controller_inst1.stoper_tr.N_214 ));
    LocalMux I__6815 (
            .O(N__34208),
            .I(\phase_controller_inst1.stoper_tr.N_214 ));
    CascadeMux I__6814 (
            .O(N__34199),
            .I(elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_));
    InMux I__6813 (
            .O(N__34196),
            .I(N__34193));
    LocalMux I__6812 (
            .O(N__34193),
            .I(N__34187));
    InMux I__6811 (
            .O(N__34192),
            .I(N__34184));
    CascadeMux I__6810 (
            .O(N__34191),
            .I(N__34181));
    CascadeMux I__6809 (
            .O(N__34190),
            .I(N__34178));
    Span4Mux_v I__6808 (
            .O(N__34187),
            .I(N__34174));
    LocalMux I__6807 (
            .O(N__34184),
            .I(N__34171));
    InMux I__6806 (
            .O(N__34181),
            .I(N__34166));
    InMux I__6805 (
            .O(N__34178),
            .I(N__34163));
    InMux I__6804 (
            .O(N__34177),
            .I(N__34160));
    Sp12to4 I__6803 (
            .O(N__34174),
            .I(N__34157));
    Span4Mux_v I__6802 (
            .O(N__34171),
            .I(N__34154));
    InMux I__6801 (
            .O(N__34170),
            .I(N__34149));
    InMux I__6800 (
            .O(N__34169),
            .I(N__34149));
    LocalMux I__6799 (
            .O(N__34166),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__6798 (
            .O(N__34163),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__6797 (
            .O(N__34160),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    Odrv12 I__6796 (
            .O(N__34157),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    Odrv4 I__6795 (
            .O(N__34154),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__6794 (
            .O(N__34149),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    CascadeMux I__6793 (
            .O(N__34136),
            .I(\phase_controller_inst1.stoper_tr.N_241_cascade_ ));
    InMux I__6792 (
            .O(N__34133),
            .I(N__34130));
    LocalMux I__6791 (
            .O(N__34130),
            .I(N__34127));
    Span4Mux_v I__6790 (
            .O(N__34127),
            .I(N__34124));
    Odrv4 I__6789 (
            .O(N__34124),
            .I(\phase_controller_inst1.stoper_tr.un6_running_1 ));
    CascadeMux I__6788 (
            .O(N__34121),
            .I(N__34117));
    CascadeMux I__6787 (
            .O(N__34120),
            .I(N__34114));
    InMux I__6786 (
            .O(N__34117),
            .I(N__34111));
    InMux I__6785 (
            .O(N__34114),
            .I(N__34107));
    LocalMux I__6784 (
            .O(N__34111),
            .I(N__34104));
    InMux I__6783 (
            .O(N__34110),
            .I(N__34101));
    LocalMux I__6782 (
            .O(N__34107),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__6781 (
            .O(N__34104),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__6780 (
            .O(N__34101),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__6779 (
            .O(N__34094),
            .I(N__34091));
    InMux I__6778 (
            .O(N__34091),
            .I(N__34088));
    LocalMux I__6777 (
            .O(N__34088),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__6776 (
            .O(N__34085),
            .I(N__34082));
    LocalMux I__6775 (
            .O(N__34082),
            .I(N__34079));
    Span4Mux_v I__6774 (
            .O(N__34079),
            .I(N__34076));
    Odrv4 I__6773 (
            .O(N__34076),
            .I(\phase_controller_inst1.stoper_tr.un6_running_2 ));
    InMux I__6772 (
            .O(N__34073),
            .I(N__34069));
    InMux I__6771 (
            .O(N__34072),
            .I(N__34066));
    LocalMux I__6770 (
            .O(N__34069),
            .I(N__34063));
    LocalMux I__6769 (
            .O(N__34066),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__6768 (
            .O(N__34063),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__6767 (
            .O(N__34058),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__6766 (
            .O(N__34055),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    InMux I__6765 (
            .O(N__34052),
            .I(N__34046));
    InMux I__6764 (
            .O(N__34051),
            .I(N__34043));
    InMux I__6763 (
            .O(N__34050),
            .I(N__34040));
    InMux I__6762 (
            .O(N__34049),
            .I(N__34037));
    LocalMux I__6761 (
            .O(N__34046),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    LocalMux I__6760 (
            .O(N__34043),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    LocalMux I__6759 (
            .O(N__34040),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    LocalMux I__6758 (
            .O(N__34037),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    InMux I__6757 (
            .O(N__34028),
            .I(N__34022));
    InMux I__6756 (
            .O(N__34027),
            .I(N__34019));
    InMux I__6755 (
            .O(N__34026),
            .I(N__34014));
    InMux I__6754 (
            .O(N__34025),
            .I(N__34014));
    LocalMux I__6753 (
            .O(N__34022),
            .I(elapsed_time_ns_1_RNIHI4DM1_0_18));
    LocalMux I__6752 (
            .O(N__34019),
            .I(elapsed_time_ns_1_RNIHI4DM1_0_18));
    LocalMux I__6751 (
            .O(N__34014),
            .I(elapsed_time_ns_1_RNIHI4DM1_0_18));
    InMux I__6750 (
            .O(N__34007),
            .I(N__34004));
    LocalMux I__6749 (
            .O(N__34004),
            .I(N__33988));
    InMux I__6748 (
            .O(N__34003),
            .I(N__33983));
    InMux I__6747 (
            .O(N__34002),
            .I(N__33983));
    InMux I__6746 (
            .O(N__34001),
            .I(N__33980));
    InMux I__6745 (
            .O(N__34000),
            .I(N__33973));
    InMux I__6744 (
            .O(N__33999),
            .I(N__33973));
    InMux I__6743 (
            .O(N__33998),
            .I(N__33973));
    InMux I__6742 (
            .O(N__33997),
            .I(N__33966));
    InMux I__6741 (
            .O(N__33996),
            .I(N__33966));
    InMux I__6740 (
            .O(N__33995),
            .I(N__33966));
    InMux I__6739 (
            .O(N__33994),
            .I(N__33957));
    InMux I__6738 (
            .O(N__33993),
            .I(N__33957));
    InMux I__6737 (
            .O(N__33992),
            .I(N__33957));
    InMux I__6736 (
            .O(N__33991),
            .I(N__33957));
    Span4Mux_h I__6735 (
            .O(N__33988),
            .I(N__33954));
    LocalMux I__6734 (
            .O(N__33983),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    LocalMux I__6733 (
            .O(N__33980),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    LocalMux I__6732 (
            .O(N__33973),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    LocalMux I__6731 (
            .O(N__33966),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    LocalMux I__6730 (
            .O(N__33957),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    Odrv4 I__6729 (
            .O(N__33954),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    InMux I__6728 (
            .O(N__33941),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__6727 (
            .O(N__33938),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__6726 (
            .O(N__33935),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__6725 (
            .O(N__33932),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__6724 (
            .O(N__33929),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__6723 (
            .O(N__33926),
            .I(bfn_15_8_0_));
    InMux I__6722 (
            .O(N__33923),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__6721 (
            .O(N__33920),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__6720 (
            .O(N__33917),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__6719 (
            .O(N__33914),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__6718 (
            .O(N__33911),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__6717 (
            .O(N__33908),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__6716 (
            .O(N__33905),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__6715 (
            .O(N__33902),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__6714 (
            .O(N__33899),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__6713 (
            .O(N__33896),
            .I(bfn_15_7_0_));
    InMux I__6712 (
            .O(N__33893),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__6711 (
            .O(N__33890),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__6710 (
            .O(N__33887),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__6709 (
            .O(N__33884),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__6708 (
            .O(N__33881),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__6707 (
            .O(N__33878),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__6706 (
            .O(N__33875),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__6705 (
            .O(N__33872),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__6704 (
            .O(N__33869),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__6703 (
            .O(N__33866),
            .I(bfn_15_6_0_));
    InMux I__6702 (
            .O(N__33863),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__6701 (
            .O(N__33860),
            .I(N__33857));
    LocalMux I__6700 (
            .O(N__33857),
            .I(N__33854));
    Odrv4 I__6699 (
            .O(N__33854),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__6698 (
            .O(N__33851),
            .I(N__33848));
    LocalMux I__6697 (
            .O(N__33848),
            .I(N__33845));
    Odrv4 I__6696 (
            .O(N__33845),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__6695 (
            .O(N__33842),
            .I(N__33839));
    LocalMux I__6694 (
            .O(N__33839),
            .I(N__33836));
    Odrv4 I__6693 (
            .O(N__33836),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__6692 (
            .O(N__33833),
            .I(N__33830));
    LocalMux I__6691 (
            .O(N__33830),
            .I(N__33827));
    Odrv4 I__6690 (
            .O(N__33827),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__6689 (
            .O(N__33824),
            .I(N__33820));
    CascadeMux I__6688 (
            .O(N__33823),
            .I(N__33817));
    LocalMux I__6687 (
            .O(N__33820),
            .I(N__33813));
    InMux I__6686 (
            .O(N__33817),
            .I(N__33810));
    InMux I__6685 (
            .O(N__33816),
            .I(N__33807));
    Odrv4 I__6684 (
            .O(N__33813),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__6683 (
            .O(N__33810),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__6682 (
            .O(N__33807),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__6681 (
            .O(N__33800),
            .I(N__33797));
    LocalMux I__6680 (
            .O(N__33797),
            .I(N__33793));
    InMux I__6679 (
            .O(N__33796),
            .I(N__33790));
    Span4Mux_v I__6678 (
            .O(N__33793),
            .I(N__33787));
    LocalMux I__6677 (
            .O(N__33790),
            .I(N__33784));
    Span4Mux_h I__6676 (
            .O(N__33787),
            .I(N__33781));
    Span4Mux_h I__6675 (
            .O(N__33784),
            .I(N__33778));
    Odrv4 I__6674 (
            .O(N__33781),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    Odrv4 I__6673 (
            .O(N__33778),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    CEMux I__6672 (
            .O(N__33773),
            .I(N__33755));
    CEMux I__6671 (
            .O(N__33772),
            .I(N__33755));
    CEMux I__6670 (
            .O(N__33771),
            .I(N__33755));
    CEMux I__6669 (
            .O(N__33770),
            .I(N__33755));
    CEMux I__6668 (
            .O(N__33769),
            .I(N__33755));
    CEMux I__6667 (
            .O(N__33768),
            .I(N__33755));
    GlobalMux I__6666 (
            .O(N__33755),
            .I(N__33752));
    gio2CtrlBuf I__6665 (
            .O(N__33752),
            .I(\delay_measurement_inst.delay_hc_timer.N_432_i_g ));
    CascadeMux I__6664 (
            .O(N__33749),
            .I(N__33743));
    InMux I__6663 (
            .O(N__33748),
            .I(N__33740));
    InMux I__6662 (
            .O(N__33747),
            .I(N__33735));
    InMux I__6661 (
            .O(N__33746),
            .I(N__33735));
    InMux I__6660 (
            .O(N__33743),
            .I(N__33732));
    LocalMux I__6659 (
            .O(N__33740),
            .I(N__33727));
    LocalMux I__6658 (
            .O(N__33735),
            .I(N__33727));
    LocalMux I__6657 (
            .O(N__33732),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__6656 (
            .O(N__33727),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    InMux I__6655 (
            .O(N__33722),
            .I(N__33719));
    LocalMux I__6654 (
            .O(N__33719),
            .I(N__33716));
    Span4Mux_h I__6653 (
            .O(N__33716),
            .I(N__33711));
    InMux I__6652 (
            .O(N__33715),
            .I(N__33708));
    InMux I__6651 (
            .O(N__33714),
            .I(N__33705));
    Span4Mux_v I__6650 (
            .O(N__33711),
            .I(N__33702));
    LocalMux I__6649 (
            .O(N__33708),
            .I(N__33699));
    LocalMux I__6648 (
            .O(N__33705),
            .I(N__33696));
    Sp12to4 I__6647 (
            .O(N__33702),
            .I(N__33689));
    Sp12to4 I__6646 (
            .O(N__33699),
            .I(N__33689));
    Span12Mux_s9_v I__6645 (
            .O(N__33696),
            .I(N__33689));
    Span12Mux_v I__6644 (
            .O(N__33689),
            .I(N__33686));
    Odrv12 I__6643 (
            .O(N__33686),
            .I(il_max_comp2_D2));
    InMux I__6642 (
            .O(N__33683),
            .I(N__33680));
    LocalMux I__6641 (
            .O(N__33680),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa ));
    IoInMux I__6640 (
            .O(N__33677),
            .I(N__33674));
    LocalMux I__6639 (
            .O(N__33674),
            .I(N__33671));
    Span4Mux_s3_v I__6638 (
            .O(N__33671),
            .I(N__33668));
    Odrv4 I__6637 (
            .O(N__33668),
            .I(\delay_measurement_inst.delay_tr_timer.N_434_i ));
    InMux I__6636 (
            .O(N__33665),
            .I(bfn_15_5_0_));
    InMux I__6635 (
            .O(N__33662),
            .I(N__33659));
    LocalMux I__6634 (
            .O(N__33659),
            .I(N__33656));
    Odrv4 I__6633 (
            .O(N__33656),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__6632 (
            .O(N__33653),
            .I(N__33650));
    LocalMux I__6631 (
            .O(N__33650),
            .I(N__33647));
    Span4Mux_h I__6630 (
            .O(N__33647),
            .I(N__33644));
    Odrv4 I__6629 (
            .O(N__33644),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__6628 (
            .O(N__33641),
            .I(N__33638));
    LocalMux I__6627 (
            .O(N__33638),
            .I(N__33635));
    Odrv12 I__6626 (
            .O(N__33635),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__6625 (
            .O(N__33632),
            .I(N__33629));
    LocalMux I__6624 (
            .O(N__33629),
            .I(N__33626));
    Odrv12 I__6623 (
            .O(N__33626),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__6622 (
            .O(N__33623),
            .I(N__33620));
    LocalMux I__6621 (
            .O(N__33620),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__6620 (
            .O(N__33617),
            .I(N__33614));
    LocalMux I__6619 (
            .O(N__33614),
            .I(N__33611));
    Odrv4 I__6618 (
            .O(N__33611),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__6617 (
            .O(N__33608),
            .I(N__33605));
    LocalMux I__6616 (
            .O(N__33605),
            .I(N__33602));
    Odrv12 I__6615 (
            .O(N__33602),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__6614 (
            .O(N__33599),
            .I(N__33596));
    LocalMux I__6613 (
            .O(N__33596),
            .I(N__33593));
    Odrv12 I__6612 (
            .O(N__33593),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__6611 (
            .O(N__33590),
            .I(N__33587));
    LocalMux I__6610 (
            .O(N__33587),
            .I(N__33584));
    Odrv12 I__6609 (
            .O(N__33584),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__6608 (
            .O(N__33581),
            .I(bfn_14_20_0_));
    InMux I__6607 (
            .O(N__33578),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__6606 (
            .O(N__33575),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__6605 (
            .O(N__33572),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__6604 (
            .O(N__33569),
            .I(N__33566));
    LocalMux I__6603 (
            .O(N__33566),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__6602 (
            .O(N__33563),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__6601 (
            .O(N__33560),
            .I(\current_shift_inst.un4_control_input1_31 ));
    CascadeMux I__6600 (
            .O(N__33557),
            .I(N__33554));
    InMux I__6599 (
            .O(N__33554),
            .I(N__33548));
    InMux I__6598 (
            .O(N__33553),
            .I(N__33548));
    LocalMux I__6597 (
            .O(N__33548),
            .I(N__33545));
    Odrv4 I__6596 (
            .O(N__33545),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    InMux I__6595 (
            .O(N__33542),
            .I(N__33539));
    LocalMux I__6594 (
            .O(N__33539),
            .I(N__33536));
    Odrv12 I__6593 (
            .O(N__33536),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__6592 (
            .O(N__33533),
            .I(N__33530));
    LocalMux I__6591 (
            .O(N__33530),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__6590 (
            .O(N__33527),
            .I(N__33524));
    LocalMux I__6589 (
            .O(N__33524),
            .I(N__33521));
    Odrv4 I__6588 (
            .O(N__33521),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__6587 (
            .O(N__33518),
            .I(N__33515));
    LocalMux I__6586 (
            .O(N__33515),
            .I(N__33512));
    Odrv4 I__6585 (
            .O(N__33512),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__6584 (
            .O(N__33509),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__6583 (
            .O(N__33506),
            .I(bfn_14_19_0_));
    InMux I__6582 (
            .O(N__33503),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__6581 (
            .O(N__33500),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__6580 (
            .O(N__33497),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__6579 (
            .O(N__33494),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__6578 (
            .O(N__33491),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__6577 (
            .O(N__33488),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__6576 (
            .O(N__33485),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__6575 (
            .O(N__33482),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__6574 (
            .O(N__33479),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__6573 (
            .O(N__33476),
            .I(N__33473));
    LocalMux I__6572 (
            .O(N__33473),
            .I(N__33470));
    Span4Mux_v I__6571 (
            .O(N__33470),
            .I(N__33467));
    Span4Mux_h I__6570 (
            .O(N__33467),
            .I(N__33464));
    Odrv4 I__6569 (
            .O(N__33464),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__6568 (
            .O(N__33461),
            .I(bfn_14_18_0_));
    InMux I__6567 (
            .O(N__33458),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__6566 (
            .O(N__33455),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__6565 (
            .O(N__33452),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__6564 (
            .O(N__33449),
            .I(N__33446));
    LocalMux I__6563 (
            .O(N__33446),
            .I(N__33443));
    Odrv4 I__6562 (
            .O(N__33443),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__6561 (
            .O(N__33440),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__6560 (
            .O(N__33437),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__6559 (
            .O(N__33434),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__6558 (
            .O(N__33431),
            .I(N__33428));
    LocalMux I__6557 (
            .O(N__33428),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    CascadeMux I__6556 (
            .O(N__33425),
            .I(N__33422));
    InMux I__6555 (
            .O(N__33422),
            .I(N__33418));
    InMux I__6554 (
            .O(N__33421),
            .I(N__33414));
    LocalMux I__6553 (
            .O(N__33418),
            .I(N__33411));
    CascadeMux I__6552 (
            .O(N__33417),
            .I(N__33407));
    LocalMux I__6551 (
            .O(N__33414),
            .I(N__33404));
    Span4Mux_v I__6550 (
            .O(N__33411),
            .I(N__33401));
    InMux I__6549 (
            .O(N__33410),
            .I(N__33398));
    InMux I__6548 (
            .O(N__33407),
            .I(N__33395));
    Odrv4 I__6547 (
            .O(N__33404),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    Odrv4 I__6546 (
            .O(N__33401),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__6545 (
            .O(N__33398),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__6544 (
            .O(N__33395),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    InMux I__6543 (
            .O(N__33386),
            .I(N__33377));
    InMux I__6542 (
            .O(N__33385),
            .I(N__33377));
    InMux I__6541 (
            .O(N__33384),
            .I(N__33377));
    LocalMux I__6540 (
            .O(N__33377),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__6539 (
            .O(N__33374),
            .I(N__33368));
    InMux I__6538 (
            .O(N__33373),
            .I(N__33368));
    LocalMux I__6537 (
            .O(N__33368),
            .I(N__33364));
    InMux I__6536 (
            .O(N__33367),
            .I(N__33361));
    Odrv4 I__6535 (
            .O(N__33364),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__6534 (
            .O(N__33361),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__6533 (
            .O(N__33356),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__6532 (
            .O(N__33353),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__6531 (
            .O(N__33350),
            .I(N__33347));
    LocalMux I__6530 (
            .O(N__33347),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__6529 (
            .O(N__33344),
            .I(N__33341));
    LocalMux I__6528 (
            .O(N__33341),
            .I(N__33336));
    InMux I__6527 (
            .O(N__33340),
            .I(N__33333));
    InMux I__6526 (
            .O(N__33339),
            .I(N__33330));
    Odrv4 I__6525 (
            .O(N__33336),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__6524 (
            .O(N__33333),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__6523 (
            .O(N__33330),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__6522 (
            .O(N__33323),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__6521 (
            .O(N__33320),
            .I(N__33317));
    LocalMux I__6520 (
            .O(N__33317),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__6519 (
            .O(N__33314),
            .I(N__33311));
    LocalMux I__6518 (
            .O(N__33311),
            .I(N__33306));
    InMux I__6517 (
            .O(N__33310),
            .I(N__33301));
    InMux I__6516 (
            .O(N__33309),
            .I(N__33301));
    Odrv4 I__6515 (
            .O(N__33306),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__6514 (
            .O(N__33301),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__6513 (
            .O(N__33296),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__6512 (
            .O(N__33293),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__6511 (
            .O(N__33290),
            .I(N__33287));
    LocalMux I__6510 (
            .O(N__33287),
            .I(\current_shift_inst.un4_control_input1_1 ));
    CascadeMux I__6509 (
            .O(N__33284),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__6508 (
            .O(N__33281),
            .I(N__33278));
    LocalMux I__6507 (
            .O(N__33278),
            .I(N__33273));
    InMux I__6506 (
            .O(N__33277),
            .I(N__33270));
    InMux I__6505 (
            .O(N__33276),
            .I(N__33267));
    Span4Mux_v I__6504 (
            .O(N__33273),
            .I(N__33264));
    LocalMux I__6503 (
            .O(N__33270),
            .I(N__33258));
    LocalMux I__6502 (
            .O(N__33267),
            .I(N__33258));
    Span4Mux_h I__6501 (
            .O(N__33264),
            .I(N__33255));
    InMux I__6500 (
            .O(N__33263),
            .I(N__33252));
    Odrv4 I__6499 (
            .O(N__33258),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    Odrv4 I__6498 (
            .O(N__33255),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__6497 (
            .O(N__33252),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    InMux I__6496 (
            .O(N__33245),
            .I(N__33241));
    InMux I__6495 (
            .O(N__33244),
            .I(N__33238));
    LocalMux I__6494 (
            .O(N__33241),
            .I(N__33235));
    LocalMux I__6493 (
            .O(N__33238),
            .I(N__33229));
    Span4Mux_v I__6492 (
            .O(N__33235),
            .I(N__33226));
    InMux I__6491 (
            .O(N__33234),
            .I(N__33219));
    InMux I__6490 (
            .O(N__33233),
            .I(N__33219));
    InMux I__6489 (
            .O(N__33232),
            .I(N__33219));
    Odrv4 I__6488 (
            .O(N__33229),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__6487 (
            .O(N__33226),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__6486 (
            .O(N__33219),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    CascadeMux I__6485 (
            .O(N__33212),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__6484 (
            .O(N__33209),
            .I(N__33206));
    LocalMux I__6483 (
            .O(N__33206),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ));
    CascadeMux I__6482 (
            .O(N__33203),
            .I(N__33200));
    InMux I__6481 (
            .O(N__33200),
            .I(N__33194));
    InMux I__6480 (
            .O(N__33199),
            .I(N__33191));
    InMux I__6479 (
            .O(N__33198),
            .I(N__33186));
    InMux I__6478 (
            .O(N__33197),
            .I(N__33186));
    LocalMux I__6477 (
            .O(N__33194),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__6476 (
            .O(N__33191),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__6475 (
            .O(N__33186),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    InMux I__6474 (
            .O(N__33179),
            .I(N__33175));
    InMux I__6473 (
            .O(N__33178),
            .I(N__33172));
    LocalMux I__6472 (
            .O(N__33175),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__6471 (
            .O(N__33172),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    CascadeMux I__6470 (
            .O(N__33167),
            .I(N__33164));
    InMux I__6469 (
            .O(N__33164),
            .I(N__33161));
    LocalMux I__6468 (
            .O(N__33161),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIP6NZ0Z32 ));
    InMux I__6467 (
            .O(N__33158),
            .I(N__33155));
    LocalMux I__6466 (
            .O(N__33155),
            .I(N__33152));
    Span4Mux_h I__6465 (
            .O(N__33152),
            .I(N__33149));
    Span4Mux_h I__6464 (
            .O(N__33149),
            .I(N__33146));
    Odrv4 I__6463 (
            .O(N__33146),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__6462 (
            .O(N__33143),
            .I(N__33140));
    LocalMux I__6461 (
            .O(N__33140),
            .I(N__33137));
    Span4Mux_v I__6460 (
            .O(N__33137),
            .I(N__33122));
    InMux I__6459 (
            .O(N__33136),
            .I(N__33117));
    InMux I__6458 (
            .O(N__33135),
            .I(N__33117));
    CascadeMux I__6457 (
            .O(N__33134),
            .I(N__33113));
    CascadeMux I__6456 (
            .O(N__33133),
            .I(N__33106));
    CascadeMux I__6455 (
            .O(N__33132),
            .I(N__33100));
    CascadeMux I__6454 (
            .O(N__33131),
            .I(N__33097));
    CascadeMux I__6453 (
            .O(N__33130),
            .I(N__33094));
    CascadeMux I__6452 (
            .O(N__33129),
            .I(N__33091));
    CascadeMux I__6451 (
            .O(N__33128),
            .I(N__33085));
    CascadeMux I__6450 (
            .O(N__33127),
            .I(N__33081));
    CascadeMux I__6449 (
            .O(N__33126),
            .I(N__33077));
    CascadeMux I__6448 (
            .O(N__33125),
            .I(N__33070));
    Span4Mux_h I__6447 (
            .O(N__33122),
            .I(N__33060));
    LocalMux I__6446 (
            .O(N__33117),
            .I(N__33060));
    InMux I__6445 (
            .O(N__33116),
            .I(N__33057));
    InMux I__6444 (
            .O(N__33113),
            .I(N__33054));
    InMux I__6443 (
            .O(N__33112),
            .I(N__33051));
    InMux I__6442 (
            .O(N__33111),
            .I(N__33043));
    InMux I__6441 (
            .O(N__33110),
            .I(N__33030));
    InMux I__6440 (
            .O(N__33109),
            .I(N__33030));
    InMux I__6439 (
            .O(N__33106),
            .I(N__33030));
    InMux I__6438 (
            .O(N__33105),
            .I(N__33030));
    InMux I__6437 (
            .O(N__33104),
            .I(N__33030));
    InMux I__6436 (
            .O(N__33103),
            .I(N__33030));
    InMux I__6435 (
            .O(N__33100),
            .I(N__33027));
    InMux I__6434 (
            .O(N__33097),
            .I(N__33024));
    InMux I__6433 (
            .O(N__33094),
            .I(N__33011));
    InMux I__6432 (
            .O(N__33091),
            .I(N__33011));
    InMux I__6431 (
            .O(N__33090),
            .I(N__33011));
    InMux I__6430 (
            .O(N__33089),
            .I(N__33011));
    InMux I__6429 (
            .O(N__33088),
            .I(N__33011));
    InMux I__6428 (
            .O(N__33085),
            .I(N__33011));
    InMux I__6427 (
            .O(N__33084),
            .I(N__33008));
    InMux I__6426 (
            .O(N__33081),
            .I(N__32993));
    InMux I__6425 (
            .O(N__33080),
            .I(N__32993));
    InMux I__6424 (
            .O(N__33077),
            .I(N__32993));
    InMux I__6423 (
            .O(N__33076),
            .I(N__32993));
    InMux I__6422 (
            .O(N__33075),
            .I(N__32993));
    InMux I__6421 (
            .O(N__33074),
            .I(N__32993));
    InMux I__6420 (
            .O(N__33073),
            .I(N__32993));
    InMux I__6419 (
            .O(N__33070),
            .I(N__32986));
    InMux I__6418 (
            .O(N__33069),
            .I(N__32986));
    InMux I__6417 (
            .O(N__33068),
            .I(N__32986));
    CascadeMux I__6416 (
            .O(N__33067),
            .I(N__32983));
    CascadeMux I__6415 (
            .O(N__33066),
            .I(N__32979));
    CascadeMux I__6414 (
            .O(N__33065),
            .I(N__32975));
    Span4Mux_v I__6413 (
            .O(N__33060),
            .I(N__32965));
    LocalMux I__6412 (
            .O(N__33057),
            .I(N__32965));
    LocalMux I__6411 (
            .O(N__33054),
            .I(N__32965));
    LocalMux I__6410 (
            .O(N__33051),
            .I(N__32965));
    InMux I__6409 (
            .O(N__33050),
            .I(N__32960));
    InMux I__6408 (
            .O(N__33049),
            .I(N__32960));
    InMux I__6407 (
            .O(N__33048),
            .I(N__32957));
    InMux I__6406 (
            .O(N__33047),
            .I(N__32954));
    InMux I__6405 (
            .O(N__33046),
            .I(N__32951));
    LocalMux I__6404 (
            .O(N__33043),
            .I(N__32938));
    LocalMux I__6403 (
            .O(N__33030),
            .I(N__32938));
    LocalMux I__6402 (
            .O(N__33027),
            .I(N__32927));
    LocalMux I__6401 (
            .O(N__33024),
            .I(N__32927));
    LocalMux I__6400 (
            .O(N__33011),
            .I(N__32927));
    LocalMux I__6399 (
            .O(N__33008),
            .I(N__32927));
    LocalMux I__6398 (
            .O(N__32993),
            .I(N__32927));
    LocalMux I__6397 (
            .O(N__32986),
            .I(N__32924));
    InMux I__6396 (
            .O(N__32983),
            .I(N__32911));
    InMux I__6395 (
            .O(N__32982),
            .I(N__32911));
    InMux I__6394 (
            .O(N__32979),
            .I(N__32911));
    InMux I__6393 (
            .O(N__32978),
            .I(N__32911));
    InMux I__6392 (
            .O(N__32975),
            .I(N__32911));
    InMux I__6391 (
            .O(N__32974),
            .I(N__32911));
    Span4Mux_v I__6390 (
            .O(N__32965),
            .I(N__32904));
    LocalMux I__6389 (
            .O(N__32960),
            .I(N__32904));
    LocalMux I__6388 (
            .O(N__32957),
            .I(N__32904));
    LocalMux I__6387 (
            .O(N__32954),
            .I(N__32899));
    LocalMux I__6386 (
            .O(N__32951),
            .I(N__32899));
    InMux I__6385 (
            .O(N__32950),
            .I(N__32882));
    InMux I__6384 (
            .O(N__32949),
            .I(N__32882));
    InMux I__6383 (
            .O(N__32948),
            .I(N__32882));
    InMux I__6382 (
            .O(N__32947),
            .I(N__32882));
    InMux I__6381 (
            .O(N__32946),
            .I(N__32882));
    InMux I__6380 (
            .O(N__32945),
            .I(N__32882));
    InMux I__6379 (
            .O(N__32944),
            .I(N__32882));
    InMux I__6378 (
            .O(N__32943),
            .I(N__32882));
    Span4Mux_v I__6377 (
            .O(N__32938),
            .I(N__32877));
    Span4Mux_v I__6376 (
            .O(N__32927),
            .I(N__32877));
    Span12Mux_v I__6375 (
            .O(N__32924),
            .I(N__32872));
    LocalMux I__6374 (
            .O(N__32911),
            .I(N__32872));
    Span4Mux_h I__6373 (
            .O(N__32904),
            .I(N__32869));
    Odrv12 I__6372 (
            .O(N__32899),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    LocalMux I__6371 (
            .O(N__32882),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__6370 (
            .O(N__32877),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv12 I__6369 (
            .O(N__32872),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__6368 (
            .O(N__32869),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    CascadeMux I__6367 (
            .O(N__32858),
            .I(N__32854));
    CascadeMux I__6366 (
            .O(N__32857),
            .I(N__32850));
    InMux I__6365 (
            .O(N__32854),
            .I(N__32843));
    InMux I__6364 (
            .O(N__32853),
            .I(N__32843));
    InMux I__6363 (
            .O(N__32850),
            .I(N__32843));
    LocalMux I__6362 (
            .O(N__32843),
            .I(N__32840));
    Span4Mux_v I__6361 (
            .O(N__32840),
            .I(N__32837));
    Odrv4 I__6360 (
            .O(N__32837),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_0_12 ));
    CascadeMux I__6359 (
            .O(N__32834),
            .I(elapsed_time_ns_1_RNIHI4DM1_0_18_cascade_));
    CascadeMux I__6358 (
            .O(N__32831),
            .I(N__32827));
    CascadeMux I__6357 (
            .O(N__32830),
            .I(N__32824));
    InMux I__6356 (
            .O(N__32827),
            .I(N__32817));
    InMux I__6355 (
            .O(N__32824),
            .I(N__32817));
    InMux I__6354 (
            .O(N__32823),
            .I(N__32814));
    InMux I__6353 (
            .O(N__32822),
            .I(N__32811));
    LocalMux I__6352 (
            .O(N__32817),
            .I(N__32808));
    LocalMux I__6351 (
            .O(N__32814),
            .I(elapsed_time_ns_1_RNIGH4DM1_0_17));
    LocalMux I__6350 (
            .O(N__32811),
            .I(elapsed_time_ns_1_RNIGH4DM1_0_17));
    Odrv4 I__6349 (
            .O(N__32808),
            .I(elapsed_time_ns_1_RNIGH4DM1_0_17));
    InMux I__6348 (
            .O(N__32801),
            .I(N__32798));
    LocalMux I__6347 (
            .O(N__32798),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9 ));
    CascadeMux I__6346 (
            .O(N__32795),
            .I(N__32791));
    InMux I__6345 (
            .O(N__32794),
            .I(N__32788));
    InMux I__6344 (
            .O(N__32791),
            .I(N__32785));
    LocalMux I__6343 (
            .O(N__32788),
            .I(N__32782));
    LocalMux I__6342 (
            .O(N__32785),
            .I(N__32779));
    Odrv4 I__6341 (
            .O(N__32782),
            .I(\phase_controller_inst1.stoper_tr.N_251 ));
    Odrv4 I__6340 (
            .O(N__32779),
            .I(\phase_controller_inst1.stoper_tr.N_251 ));
    CascadeMux I__6339 (
            .O(N__32774),
            .I(elapsed_time_ns_1_RNISCJF91_0_31_cascade_));
    InMux I__6338 (
            .O(N__32771),
            .I(N__32768));
    LocalMux I__6337 (
            .O(N__32768),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9 ));
    InMux I__6336 (
            .O(N__32765),
            .I(N__32760));
    InMux I__6335 (
            .O(N__32764),
            .I(N__32755));
    InMux I__6334 (
            .O(N__32763),
            .I(N__32755));
    LocalMux I__6333 (
            .O(N__32760),
            .I(N__32748));
    LocalMux I__6332 (
            .O(N__32755),
            .I(N__32748));
    InMux I__6331 (
            .O(N__32754),
            .I(N__32743));
    InMux I__6330 (
            .O(N__32753),
            .I(N__32743));
    Odrv4 I__6329 (
            .O(N__32748),
            .I(elapsed_time_ns_1_RNI1OL2M1_0_9));
    LocalMux I__6328 (
            .O(N__32743),
            .I(elapsed_time_ns_1_RNI1OL2M1_0_9));
    CascadeMux I__6327 (
            .O(N__32738),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_ ));
    CascadeMux I__6326 (
            .O(N__32735),
            .I(N__32731));
    InMux I__6325 (
            .O(N__32734),
            .I(N__32727));
    InMux I__6324 (
            .O(N__32731),
            .I(N__32724));
    InMux I__6323 (
            .O(N__32730),
            .I(N__32721));
    LocalMux I__6322 (
            .O(N__32727),
            .I(N__32717));
    LocalMux I__6321 (
            .O(N__32724),
            .I(N__32712));
    LocalMux I__6320 (
            .O(N__32721),
            .I(N__32712));
    InMux I__6319 (
            .O(N__32720),
            .I(N__32709));
    Span4Mux_h I__6318 (
            .O(N__32717),
            .I(N__32706));
    Odrv4 I__6317 (
            .O(N__32712),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__6316 (
            .O(N__32709),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__6315 (
            .O(N__32706),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    CascadeMux I__6314 (
            .O(N__32699),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0_cascade_ ));
    InMux I__6313 (
            .O(N__32696),
            .I(N__32690));
    InMux I__6312 (
            .O(N__32695),
            .I(N__32690));
    LocalMux I__6311 (
            .O(N__32690),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    CascadeMux I__6310 (
            .O(N__32687),
            .I(elapsed_time_ns_1_RNICG2591_0_4_cascade_));
    InMux I__6309 (
            .O(N__32684),
            .I(N__32681));
    LocalMux I__6308 (
            .O(N__32681),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2 ));
    CascadeMux I__6307 (
            .O(N__32678),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16_cascade_ ));
    CascadeMux I__6306 (
            .O(N__32675),
            .I(N__32671));
    InMux I__6305 (
            .O(N__32674),
            .I(N__32665));
    InMux I__6304 (
            .O(N__32671),
            .I(N__32662));
    InMux I__6303 (
            .O(N__32670),
            .I(N__32655));
    InMux I__6302 (
            .O(N__32669),
            .I(N__32655));
    InMux I__6301 (
            .O(N__32668),
            .I(N__32655));
    LocalMux I__6300 (
            .O(N__32665),
            .I(elapsed_time_ns_1_RNIFG4DM1_0_16));
    LocalMux I__6299 (
            .O(N__32662),
            .I(elapsed_time_ns_1_RNIFG4DM1_0_16));
    LocalMux I__6298 (
            .O(N__32655),
            .I(elapsed_time_ns_1_RNIFG4DM1_0_16));
    CascadeMux I__6297 (
            .O(N__32648),
            .I(elapsed_time_ns_1_RNIGH4DM1_0_17_cascade_));
    InMux I__6296 (
            .O(N__32645),
            .I(N__32642));
    LocalMux I__6295 (
            .O(N__32642),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17 ));
    CascadeMux I__6294 (
            .O(N__32639),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18_cascade_ ));
    CascadeMux I__6293 (
            .O(N__32636),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15_cascade_));
    InMux I__6292 (
            .O(N__32633),
            .I(N__32630));
    LocalMux I__6291 (
            .O(N__32630),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9 ));
    CascadeMux I__6290 (
            .O(N__32627),
            .I(elapsed_time_ns_1_RNI1OL2M1_0_9_cascade_));
    CascadeMux I__6289 (
            .O(N__32624),
            .I(\phase_controller_inst1.stoper_tr.N_211_cascade_ ));
    CascadeMux I__6288 (
            .O(N__32621),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6_cascade_ ));
    InMux I__6287 (
            .O(N__32618),
            .I(N__32615));
    LocalMux I__6286 (
            .O(N__32615),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1 ));
    InMux I__6285 (
            .O(N__32612),
            .I(N__32605));
    InMux I__6284 (
            .O(N__32611),
            .I(N__32605));
    InMux I__6283 (
            .O(N__32610),
            .I(N__32602));
    LocalMux I__6282 (
            .O(N__32605),
            .I(elapsed_time_ns_1_RNIPFL2M1_0_1));
    LocalMux I__6281 (
            .O(N__32602),
            .I(elapsed_time_ns_1_RNIPFL2M1_0_1));
    InMux I__6280 (
            .O(N__32597),
            .I(N__32593));
    InMux I__6279 (
            .O(N__32596),
            .I(N__32590));
    LocalMux I__6278 (
            .O(N__32593),
            .I(N__32587));
    LocalMux I__6277 (
            .O(N__32590),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1 ));
    Odrv4 I__6276 (
            .O(N__32587),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1 ));
    CascadeMux I__6275 (
            .O(N__32582),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_ ));
    CascadeMux I__6274 (
            .O(N__32579),
            .I(N__32571));
    CascadeMux I__6273 (
            .O(N__32578),
            .I(N__32568));
    CascadeMux I__6272 (
            .O(N__32577),
            .I(N__32564));
    CascadeMux I__6271 (
            .O(N__32576),
            .I(N__32561));
    CascadeMux I__6270 (
            .O(N__32575),
            .I(N__32555));
    CascadeMux I__6269 (
            .O(N__32574),
            .I(N__32552));
    InMux I__6268 (
            .O(N__32571),
            .I(N__32548));
    InMux I__6267 (
            .O(N__32568),
            .I(N__32545));
    InMux I__6266 (
            .O(N__32567),
            .I(N__32542));
    InMux I__6265 (
            .O(N__32564),
            .I(N__32539));
    InMux I__6264 (
            .O(N__32561),
            .I(N__32534));
    InMux I__6263 (
            .O(N__32560),
            .I(N__32534));
    InMux I__6262 (
            .O(N__32559),
            .I(N__32523));
    InMux I__6261 (
            .O(N__32558),
            .I(N__32523));
    InMux I__6260 (
            .O(N__32555),
            .I(N__32523));
    InMux I__6259 (
            .O(N__32552),
            .I(N__32523));
    InMux I__6258 (
            .O(N__32551),
            .I(N__32523));
    LocalMux I__6257 (
            .O(N__32548),
            .I(N__32518));
    LocalMux I__6256 (
            .O(N__32545),
            .I(N__32518));
    LocalMux I__6255 (
            .O(N__32542),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    LocalMux I__6254 (
            .O(N__32539),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    LocalMux I__6253 (
            .O(N__32534),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    LocalMux I__6252 (
            .O(N__32523),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    Odrv12 I__6251 (
            .O(N__32518),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    InMux I__6250 (
            .O(N__32507),
            .I(N__32498));
    InMux I__6249 (
            .O(N__32506),
            .I(N__32498));
    InMux I__6248 (
            .O(N__32505),
            .I(N__32498));
    LocalMux I__6247 (
            .O(N__32498),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2 ));
    CascadeMux I__6246 (
            .O(N__32495),
            .I(N__32491));
    InMux I__6245 (
            .O(N__32494),
            .I(N__32488));
    InMux I__6244 (
            .O(N__32491),
            .I(N__32485));
    LocalMux I__6243 (
            .O(N__32488),
            .I(N__32479));
    LocalMux I__6242 (
            .O(N__32485),
            .I(N__32479));
    InMux I__6241 (
            .O(N__32484),
            .I(N__32476));
    Odrv4 I__6240 (
            .O(N__32479),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    LocalMux I__6239 (
            .O(N__32476),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    CEMux I__6238 (
            .O(N__32471),
            .I(N__32466));
    CEMux I__6237 (
            .O(N__32470),
            .I(N__32463));
    CEMux I__6236 (
            .O(N__32469),
            .I(N__32459));
    LocalMux I__6235 (
            .O(N__32466),
            .I(N__32454));
    LocalMux I__6234 (
            .O(N__32463),
            .I(N__32454));
    CEMux I__6233 (
            .O(N__32462),
            .I(N__32451));
    LocalMux I__6232 (
            .O(N__32459),
            .I(N__32448));
    Span4Mux_v I__6231 (
            .O(N__32454),
            .I(N__32445));
    LocalMux I__6230 (
            .O(N__32451),
            .I(N__32442));
    Span4Mux_v I__6229 (
            .O(N__32448),
            .I(N__32435));
    Span4Mux_h I__6228 (
            .O(N__32445),
            .I(N__32435));
    Span4Mux_h I__6227 (
            .O(N__32442),
            .I(N__32435));
    Span4Mux_h I__6226 (
            .O(N__32435),
            .I(N__32432));
    Odrv4 I__6225 (
            .O(N__32432),
            .I(\delay_measurement_inst.delay_hc_timer.N_433_i ));
    InMux I__6224 (
            .O(N__32429),
            .I(N__32425));
    InMux I__6223 (
            .O(N__32428),
            .I(N__32420));
    LocalMux I__6222 (
            .O(N__32425),
            .I(N__32417));
    InMux I__6221 (
            .O(N__32424),
            .I(N__32412));
    InMux I__6220 (
            .O(N__32423),
            .I(N__32412));
    LocalMux I__6219 (
            .O(N__32420),
            .I(N__32407));
    Span12Mux_s7_v I__6218 (
            .O(N__32417),
            .I(N__32407));
    LocalMux I__6217 (
            .O(N__32412),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv12 I__6216 (
            .O(N__32407),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    IoInMux I__6215 (
            .O(N__32402),
            .I(N__32399));
    LocalMux I__6214 (
            .O(N__32399),
            .I(N__32396));
    Odrv12 I__6213 (
            .O(N__32396),
            .I(\current_shift_inst.timer_s1.N_166_i ));
    CascadeMux I__6212 (
            .O(N__32393),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_ ));
    CascadeMux I__6211 (
            .O(N__32390),
            .I(elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_));
    CascadeMux I__6210 (
            .O(N__32387),
            .I(N__32383));
    CascadeMux I__6209 (
            .O(N__32386),
            .I(N__32379));
    InMux I__6208 (
            .O(N__32383),
            .I(N__32376));
    InMux I__6207 (
            .O(N__32382),
            .I(N__32373));
    InMux I__6206 (
            .O(N__32379),
            .I(N__32370));
    LocalMux I__6205 (
            .O(N__32376),
            .I(elapsed_time_ns_1_RNIUKL2M1_0_6));
    LocalMux I__6204 (
            .O(N__32373),
            .I(elapsed_time_ns_1_RNIUKL2M1_0_6));
    LocalMux I__6203 (
            .O(N__32370),
            .I(elapsed_time_ns_1_RNIUKL2M1_0_6));
    InMux I__6202 (
            .O(N__32363),
            .I(N__32359));
    InMux I__6201 (
            .O(N__32362),
            .I(N__32356));
    LocalMux I__6200 (
            .O(N__32359),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ));
    LocalMux I__6199 (
            .O(N__32356),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ));
    CascadeMux I__6198 (
            .O(N__32351),
            .I(N__32348));
    InMux I__6197 (
            .O(N__32348),
            .I(N__32343));
    InMux I__6196 (
            .O(N__32347),
            .I(N__32340));
    InMux I__6195 (
            .O(N__32346),
            .I(N__32337));
    LocalMux I__6194 (
            .O(N__32343),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__6193 (
            .O(N__32340),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__6192 (
            .O(N__32337),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__6191 (
            .O(N__32330),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__6190 (
            .O(N__32327),
            .I(N__32322));
    InMux I__6189 (
            .O(N__32326),
            .I(N__32317));
    InMux I__6188 (
            .O(N__32325),
            .I(N__32317));
    LocalMux I__6187 (
            .O(N__32322),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__6186 (
            .O(N__32317),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__6185 (
            .O(N__32312),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__6184 (
            .O(N__32309),
            .I(N__32304));
    InMux I__6183 (
            .O(N__32308),
            .I(N__32299));
    InMux I__6182 (
            .O(N__32307),
            .I(N__32299));
    LocalMux I__6181 (
            .O(N__32304),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__6180 (
            .O(N__32299),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__6179 (
            .O(N__32294),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    CascadeMux I__6178 (
            .O(N__32291),
            .I(N__32287));
    CascadeMux I__6177 (
            .O(N__32290),
            .I(N__32284));
    InMux I__6176 (
            .O(N__32287),
            .I(N__32280));
    InMux I__6175 (
            .O(N__32284),
            .I(N__32277));
    InMux I__6174 (
            .O(N__32283),
            .I(N__32274));
    LocalMux I__6173 (
            .O(N__32280),
            .I(N__32271));
    LocalMux I__6172 (
            .O(N__32277),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__6171 (
            .O(N__32274),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__6170 (
            .O(N__32271),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__6169 (
            .O(N__32264),
            .I(bfn_13_24_0_));
    CascadeMux I__6168 (
            .O(N__32261),
            .I(N__32257));
    CascadeMux I__6167 (
            .O(N__32260),
            .I(N__32254));
    InMux I__6166 (
            .O(N__32257),
            .I(N__32250));
    InMux I__6165 (
            .O(N__32254),
            .I(N__32247));
    InMux I__6164 (
            .O(N__32253),
            .I(N__32244));
    LocalMux I__6163 (
            .O(N__32250),
            .I(N__32241));
    LocalMux I__6162 (
            .O(N__32247),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__6161 (
            .O(N__32244),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__6160 (
            .O(N__32241),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__6159 (
            .O(N__32234),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    CascadeMux I__6158 (
            .O(N__32231),
            .I(N__32228));
    InMux I__6157 (
            .O(N__32228),
            .I(N__32223));
    InMux I__6156 (
            .O(N__32227),
            .I(N__32220));
    InMux I__6155 (
            .O(N__32226),
            .I(N__32217));
    LocalMux I__6154 (
            .O(N__32223),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__6153 (
            .O(N__32220),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__6152 (
            .O(N__32217),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__6151 (
            .O(N__32210),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    CascadeMux I__6150 (
            .O(N__32207),
            .I(N__32204));
    InMux I__6149 (
            .O(N__32204),
            .I(N__32199));
    InMux I__6148 (
            .O(N__32203),
            .I(N__32196));
    InMux I__6147 (
            .O(N__32202),
            .I(N__32193));
    LocalMux I__6146 (
            .O(N__32199),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__6145 (
            .O(N__32196),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__6144 (
            .O(N__32193),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__6143 (
            .O(N__32186),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__6142 (
            .O(N__32183),
            .I(N__32179));
    InMux I__6141 (
            .O(N__32182),
            .I(N__32176));
    LocalMux I__6140 (
            .O(N__32179),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    LocalMux I__6139 (
            .O(N__32176),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__6138 (
            .O(N__32171),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__6137 (
            .O(N__32168),
            .I(N__32130));
    InMux I__6136 (
            .O(N__32167),
            .I(N__32130));
    InMux I__6135 (
            .O(N__32166),
            .I(N__32130));
    InMux I__6134 (
            .O(N__32165),
            .I(N__32130));
    InMux I__6133 (
            .O(N__32164),
            .I(N__32125));
    InMux I__6132 (
            .O(N__32163),
            .I(N__32125));
    InMux I__6131 (
            .O(N__32162),
            .I(N__32116));
    InMux I__6130 (
            .O(N__32161),
            .I(N__32116));
    InMux I__6129 (
            .O(N__32160),
            .I(N__32116));
    InMux I__6128 (
            .O(N__32159),
            .I(N__32116));
    InMux I__6127 (
            .O(N__32158),
            .I(N__32107));
    InMux I__6126 (
            .O(N__32157),
            .I(N__32107));
    InMux I__6125 (
            .O(N__32156),
            .I(N__32107));
    InMux I__6124 (
            .O(N__32155),
            .I(N__32107));
    InMux I__6123 (
            .O(N__32154),
            .I(N__32098));
    InMux I__6122 (
            .O(N__32153),
            .I(N__32098));
    InMux I__6121 (
            .O(N__32152),
            .I(N__32098));
    InMux I__6120 (
            .O(N__32151),
            .I(N__32098));
    InMux I__6119 (
            .O(N__32150),
            .I(N__32089));
    InMux I__6118 (
            .O(N__32149),
            .I(N__32089));
    InMux I__6117 (
            .O(N__32148),
            .I(N__32089));
    InMux I__6116 (
            .O(N__32147),
            .I(N__32089));
    InMux I__6115 (
            .O(N__32146),
            .I(N__32080));
    InMux I__6114 (
            .O(N__32145),
            .I(N__32080));
    InMux I__6113 (
            .O(N__32144),
            .I(N__32080));
    InMux I__6112 (
            .O(N__32143),
            .I(N__32080));
    InMux I__6111 (
            .O(N__32142),
            .I(N__32071));
    InMux I__6110 (
            .O(N__32141),
            .I(N__32071));
    InMux I__6109 (
            .O(N__32140),
            .I(N__32071));
    InMux I__6108 (
            .O(N__32139),
            .I(N__32071));
    LocalMux I__6107 (
            .O(N__32130),
            .I(N__32068));
    LocalMux I__6106 (
            .O(N__32125),
            .I(N__32057));
    LocalMux I__6105 (
            .O(N__32116),
            .I(N__32057));
    LocalMux I__6104 (
            .O(N__32107),
            .I(N__32057));
    LocalMux I__6103 (
            .O(N__32098),
            .I(N__32057));
    LocalMux I__6102 (
            .O(N__32089),
            .I(N__32057));
    LocalMux I__6101 (
            .O(N__32080),
            .I(N__32052));
    LocalMux I__6100 (
            .O(N__32071),
            .I(N__32052));
    Span4Mux_v I__6099 (
            .O(N__32068),
            .I(N__32047));
    Span4Mux_v I__6098 (
            .O(N__32057),
            .I(N__32047));
    Span4Mux_h I__6097 (
            .O(N__32052),
            .I(N__32044));
    Odrv4 I__6096 (
            .O(N__32047),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__6095 (
            .O(N__32044),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__6094 (
            .O(N__32039),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__6093 (
            .O(N__32036),
            .I(N__32032));
    InMux I__6092 (
            .O(N__32035),
            .I(N__32029));
    LocalMux I__6091 (
            .O(N__32032),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    LocalMux I__6090 (
            .O(N__32029),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__6089 (
            .O(N__32024),
            .I(N__32021));
    InMux I__6088 (
            .O(N__32021),
            .I(N__32016));
    InMux I__6087 (
            .O(N__32020),
            .I(N__32013));
    InMux I__6086 (
            .O(N__32019),
            .I(N__32010));
    LocalMux I__6085 (
            .O(N__32016),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__6084 (
            .O(N__32013),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__6083 (
            .O(N__32010),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__6082 (
            .O(N__32003),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__6081 (
            .O(N__32000),
            .I(N__31995));
    InMux I__6080 (
            .O(N__31999),
            .I(N__31990));
    InMux I__6079 (
            .O(N__31998),
            .I(N__31990));
    LocalMux I__6078 (
            .O(N__31995),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__6077 (
            .O(N__31990),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__6076 (
            .O(N__31985),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__6075 (
            .O(N__31982),
            .I(N__31977));
    InMux I__6074 (
            .O(N__31981),
            .I(N__31972));
    InMux I__6073 (
            .O(N__31980),
            .I(N__31972));
    LocalMux I__6072 (
            .O(N__31977),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__6071 (
            .O(N__31972),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__6070 (
            .O(N__31967),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    CascadeMux I__6069 (
            .O(N__31964),
            .I(N__31961));
    InMux I__6068 (
            .O(N__31961),
            .I(N__31957));
    CascadeMux I__6067 (
            .O(N__31960),
            .I(N__31954));
    LocalMux I__6066 (
            .O(N__31957),
            .I(N__31950));
    InMux I__6065 (
            .O(N__31954),
            .I(N__31947));
    InMux I__6064 (
            .O(N__31953),
            .I(N__31944));
    Span4Mux_h I__6063 (
            .O(N__31950),
            .I(N__31941));
    LocalMux I__6062 (
            .O(N__31947),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__6061 (
            .O(N__31944),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__6060 (
            .O(N__31941),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__6059 (
            .O(N__31934),
            .I(bfn_13_23_0_));
    CascadeMux I__6058 (
            .O(N__31931),
            .I(N__31927));
    CascadeMux I__6057 (
            .O(N__31930),
            .I(N__31924));
    InMux I__6056 (
            .O(N__31927),
            .I(N__31920));
    InMux I__6055 (
            .O(N__31924),
            .I(N__31917));
    InMux I__6054 (
            .O(N__31923),
            .I(N__31914));
    LocalMux I__6053 (
            .O(N__31920),
            .I(N__31911));
    LocalMux I__6052 (
            .O(N__31917),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__6051 (
            .O(N__31914),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__6050 (
            .O(N__31911),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__6049 (
            .O(N__31904),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__6048 (
            .O(N__31901),
            .I(N__31897));
    CascadeMux I__6047 (
            .O(N__31900),
            .I(N__31894));
    LocalMux I__6046 (
            .O(N__31897),
            .I(N__31890));
    InMux I__6045 (
            .O(N__31894),
            .I(N__31887));
    InMux I__6044 (
            .O(N__31893),
            .I(N__31884));
    Span4Mux_h I__6043 (
            .O(N__31890),
            .I(N__31881));
    LocalMux I__6042 (
            .O(N__31887),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__6041 (
            .O(N__31884),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv4 I__6040 (
            .O(N__31881),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__6039 (
            .O(N__31874),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    CascadeMux I__6038 (
            .O(N__31871),
            .I(N__31868));
    InMux I__6037 (
            .O(N__31868),
            .I(N__31863));
    InMux I__6036 (
            .O(N__31867),
            .I(N__31860));
    InMux I__6035 (
            .O(N__31866),
            .I(N__31857));
    LocalMux I__6034 (
            .O(N__31863),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__6033 (
            .O(N__31860),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__6032 (
            .O(N__31857),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__6031 (
            .O(N__31850),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    CascadeMux I__6030 (
            .O(N__31847),
            .I(N__31844));
    InMux I__6029 (
            .O(N__31844),
            .I(N__31839));
    InMux I__6028 (
            .O(N__31843),
            .I(N__31836));
    InMux I__6027 (
            .O(N__31842),
            .I(N__31833));
    LocalMux I__6026 (
            .O(N__31839),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__6025 (
            .O(N__31836),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__6024 (
            .O(N__31833),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__6023 (
            .O(N__31826),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__6022 (
            .O(N__31823),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    CascadeMux I__6021 (
            .O(N__31820),
            .I(N__31817));
    InMux I__6020 (
            .O(N__31817),
            .I(N__31812));
    InMux I__6019 (
            .O(N__31816),
            .I(N__31809));
    InMux I__6018 (
            .O(N__31815),
            .I(N__31806));
    LocalMux I__6017 (
            .O(N__31812),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__6016 (
            .O(N__31809),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__6015 (
            .O(N__31806),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__6014 (
            .O(N__31799),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__6013 (
            .O(N__31796),
            .I(N__31791));
    InMux I__6012 (
            .O(N__31795),
            .I(N__31786));
    InMux I__6011 (
            .O(N__31794),
            .I(N__31786));
    LocalMux I__6010 (
            .O(N__31791),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__6009 (
            .O(N__31786),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__6008 (
            .O(N__31781),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__6007 (
            .O(N__31778),
            .I(N__31773));
    InMux I__6006 (
            .O(N__31777),
            .I(N__31768));
    InMux I__6005 (
            .O(N__31776),
            .I(N__31768));
    LocalMux I__6004 (
            .O(N__31773),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__6003 (
            .O(N__31768),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__6002 (
            .O(N__31763),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    CascadeMux I__6001 (
            .O(N__31760),
            .I(N__31756));
    CascadeMux I__6000 (
            .O(N__31759),
            .I(N__31753));
    InMux I__5999 (
            .O(N__31756),
            .I(N__31749));
    InMux I__5998 (
            .O(N__31753),
            .I(N__31746));
    InMux I__5997 (
            .O(N__31752),
            .I(N__31743));
    LocalMux I__5996 (
            .O(N__31749),
            .I(N__31740));
    LocalMux I__5995 (
            .O(N__31746),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__5994 (
            .O(N__31743),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__5993 (
            .O(N__31740),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__5992 (
            .O(N__31733),
            .I(bfn_13_22_0_));
    CascadeMux I__5991 (
            .O(N__31730),
            .I(N__31726));
    CascadeMux I__5990 (
            .O(N__31729),
            .I(N__31723));
    InMux I__5989 (
            .O(N__31726),
            .I(N__31719));
    InMux I__5988 (
            .O(N__31723),
            .I(N__31716));
    InMux I__5987 (
            .O(N__31722),
            .I(N__31713));
    LocalMux I__5986 (
            .O(N__31719),
            .I(N__31710));
    LocalMux I__5985 (
            .O(N__31716),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__5984 (
            .O(N__31713),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__5983 (
            .O(N__31710),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__5982 (
            .O(N__31703),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    CascadeMux I__5981 (
            .O(N__31700),
            .I(N__31697));
    InMux I__5980 (
            .O(N__31697),
            .I(N__31692));
    InMux I__5979 (
            .O(N__31696),
            .I(N__31689));
    InMux I__5978 (
            .O(N__31695),
            .I(N__31686));
    LocalMux I__5977 (
            .O(N__31692),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__5976 (
            .O(N__31689),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__5975 (
            .O(N__31686),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__5974 (
            .O(N__31679),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    CascadeMux I__5973 (
            .O(N__31676),
            .I(N__31673));
    InMux I__5972 (
            .O(N__31673),
            .I(N__31668));
    InMux I__5971 (
            .O(N__31672),
            .I(N__31665));
    InMux I__5970 (
            .O(N__31671),
            .I(N__31662));
    LocalMux I__5969 (
            .O(N__31668),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__5968 (
            .O(N__31665),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__5967 (
            .O(N__31662),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__5966 (
            .O(N__31655),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    CascadeMux I__5965 (
            .O(N__31652),
            .I(N__31649));
    InMux I__5964 (
            .O(N__31649),
            .I(N__31644));
    InMux I__5963 (
            .O(N__31648),
            .I(N__31641));
    InMux I__5962 (
            .O(N__31647),
            .I(N__31638));
    LocalMux I__5961 (
            .O(N__31644),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__5960 (
            .O(N__31641),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__5959 (
            .O(N__31638),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__5958 (
            .O(N__31631),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__5957 (
            .O(N__31628),
            .I(N__31625));
    LocalMux I__5956 (
            .O(N__31625),
            .I(N__31622));
    Span4Mux_h I__5955 (
            .O(N__31622),
            .I(N__31619));
    Span4Mux_h I__5954 (
            .O(N__31619),
            .I(N__31616));
    Odrv4 I__5953 (
            .O(N__31616),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__5952 (
            .O(N__31613),
            .I(bfn_13_21_0_));
    InMux I__5951 (
            .O(N__31610),
            .I(N__31607));
    LocalMux I__5950 (
            .O(N__31607),
            .I(N__31604));
    Span4Mux_h I__5949 (
            .O(N__31604),
            .I(N__31600));
    CascadeMux I__5948 (
            .O(N__31603),
            .I(N__31597));
    Span4Mux_h I__5947 (
            .O(N__31600),
            .I(N__31593));
    InMux I__5946 (
            .O(N__31597),
            .I(N__31590));
    InMux I__5945 (
            .O(N__31596),
            .I(N__31587));
    Odrv4 I__5944 (
            .O(N__31593),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__5943 (
            .O(N__31590),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__5942 (
            .O(N__31587),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__5941 (
            .O(N__31580),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    CascadeMux I__5940 (
            .O(N__31577),
            .I(N__31574));
    InMux I__5939 (
            .O(N__31574),
            .I(N__31569));
    InMux I__5938 (
            .O(N__31573),
            .I(N__31566));
    InMux I__5937 (
            .O(N__31572),
            .I(N__31563));
    LocalMux I__5936 (
            .O(N__31569),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__5935 (
            .O(N__31566),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__5934 (
            .O(N__31563),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__5933 (
            .O(N__31556),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    CascadeMux I__5932 (
            .O(N__31553),
            .I(N__31550));
    InMux I__5931 (
            .O(N__31550),
            .I(N__31545));
    InMux I__5930 (
            .O(N__31549),
            .I(N__31542));
    InMux I__5929 (
            .O(N__31548),
            .I(N__31539));
    LocalMux I__5928 (
            .O(N__31545),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__5927 (
            .O(N__31542),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__5926 (
            .O(N__31539),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__5925 (
            .O(N__31532),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    CascadeMux I__5924 (
            .O(N__31529),
            .I(N__31526));
    InMux I__5923 (
            .O(N__31526),
            .I(N__31521));
    InMux I__5922 (
            .O(N__31525),
            .I(N__31518));
    InMux I__5921 (
            .O(N__31524),
            .I(N__31515));
    LocalMux I__5920 (
            .O(N__31521),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__5919 (
            .O(N__31518),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__5918 (
            .O(N__31515),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__5917 (
            .O(N__31508),
            .I(N__31504));
    CascadeMux I__5916 (
            .O(N__31507),
            .I(N__31499));
    LocalMux I__5915 (
            .O(N__31504),
            .I(N__31496));
    InMux I__5914 (
            .O(N__31503),
            .I(N__31489));
    InMux I__5913 (
            .O(N__31502),
            .I(N__31489));
    InMux I__5912 (
            .O(N__31499),
            .I(N__31489));
    Span4Mux_v I__5911 (
            .O(N__31496),
            .I(N__31486));
    LocalMux I__5910 (
            .O(N__31489),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv4 I__5909 (
            .O(N__31486),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    CascadeMux I__5908 (
            .O(N__31481),
            .I(N__31477));
    InMux I__5907 (
            .O(N__31480),
            .I(N__31466));
    InMux I__5906 (
            .O(N__31477),
            .I(N__31466));
    InMux I__5905 (
            .O(N__31476),
            .I(N__31466));
    InMux I__5904 (
            .O(N__31475),
            .I(N__31466));
    LocalMux I__5903 (
            .O(N__31466),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    CascadeMux I__5902 (
            .O(N__31463),
            .I(N__31460));
    InMux I__5901 (
            .O(N__31460),
            .I(N__31456));
    InMux I__5900 (
            .O(N__31459),
            .I(N__31452));
    LocalMux I__5899 (
            .O(N__31456),
            .I(N__31449));
    InMux I__5898 (
            .O(N__31455),
            .I(N__31445));
    LocalMux I__5897 (
            .O(N__31452),
            .I(N__31442));
    Span4Mux_h I__5896 (
            .O(N__31449),
            .I(N__31439));
    InMux I__5895 (
            .O(N__31448),
            .I(N__31436));
    LocalMux I__5894 (
            .O(N__31445),
            .I(N__31431));
    Span4Mux_h I__5893 (
            .O(N__31442),
            .I(N__31431));
    Span4Mux_h I__5892 (
            .O(N__31439),
            .I(N__31428));
    LocalMux I__5891 (
            .O(N__31436),
            .I(N__31423));
    Span4Mux_v I__5890 (
            .O(N__31431),
            .I(N__31423));
    Odrv4 I__5889 (
            .O(N__31428),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__5888 (
            .O(N__31423),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__5887 (
            .O(N__31418),
            .I(N__31415));
    LocalMux I__5886 (
            .O(N__31415),
            .I(N__31412));
    Odrv12 I__5885 (
            .O(N__31412),
            .I(\current_shift_inst.PI_CTRL.integrator_i_30 ));
    InMux I__5884 (
            .O(N__31409),
            .I(N__31405));
    InMux I__5883 (
            .O(N__31408),
            .I(N__31402));
    LocalMux I__5882 (
            .O(N__31405),
            .I(N__31398));
    LocalMux I__5881 (
            .O(N__31402),
            .I(N__31395));
    InMux I__5880 (
            .O(N__31401),
            .I(N__31392));
    Span4Mux_v I__5879 (
            .O(N__31398),
            .I(N__31387));
    Span4Mux_v I__5878 (
            .O(N__31395),
            .I(N__31384));
    LocalMux I__5877 (
            .O(N__31392),
            .I(N__31381));
    InMux I__5876 (
            .O(N__31391),
            .I(N__31376));
    InMux I__5875 (
            .O(N__31390),
            .I(N__31376));
    Span4Mux_v I__5874 (
            .O(N__31387),
            .I(N__31369));
    Span4Mux_h I__5873 (
            .O(N__31384),
            .I(N__31369));
    Span4Mux_v I__5872 (
            .O(N__31381),
            .I(N__31369));
    LocalMux I__5871 (
            .O(N__31376),
            .I(N__31366));
    Odrv4 I__5870 (
            .O(N__31369),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv12 I__5869 (
            .O(N__31366),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__5868 (
            .O(N__31361),
            .I(N__31358));
    LocalMux I__5867 (
            .O(N__31358),
            .I(N__31355));
    Odrv12 I__5866 (
            .O(N__31355),
            .I(\current_shift_inst.PI_CTRL.integrator_i_27 ));
    CascadeMux I__5865 (
            .O(N__31352),
            .I(N__31349));
    InMux I__5864 (
            .O(N__31349),
            .I(N__31346));
    LocalMux I__5863 (
            .O(N__31346),
            .I(N__31342));
    CascadeMux I__5862 (
            .O(N__31345),
            .I(N__31339));
    Span4Mux_v I__5861 (
            .O(N__31342),
            .I(N__31335));
    InMux I__5860 (
            .O(N__31339),
            .I(N__31329));
    InMux I__5859 (
            .O(N__31338),
            .I(N__31329));
    Span4Mux_h I__5858 (
            .O(N__31335),
            .I(N__31326));
    InMux I__5857 (
            .O(N__31334),
            .I(N__31323));
    LocalMux I__5856 (
            .O(N__31329),
            .I(N__31320));
    Span4Mux_h I__5855 (
            .O(N__31326),
            .I(N__31315));
    LocalMux I__5854 (
            .O(N__31323),
            .I(N__31315));
    Span4Mux_h I__5853 (
            .O(N__31320),
            .I(N__31312));
    Odrv4 I__5852 (
            .O(N__31315),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__5851 (
            .O(N__31312),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__5850 (
            .O(N__31307),
            .I(N__31304));
    LocalMux I__5849 (
            .O(N__31304),
            .I(N__31301));
    Odrv12 I__5848 (
            .O(N__31301),
            .I(\current_shift_inst.PI_CTRL.integrator_i_28 ));
    CascadeMux I__5847 (
            .O(N__31298),
            .I(N__31295));
    InMux I__5846 (
            .O(N__31295),
            .I(N__31291));
    InMux I__5845 (
            .O(N__31294),
            .I(N__31288));
    LocalMux I__5844 (
            .O(N__31291),
            .I(N__31282));
    LocalMux I__5843 (
            .O(N__31288),
            .I(N__31282));
    InMux I__5842 (
            .O(N__31287),
            .I(N__31279));
    Span4Mux_h I__5841 (
            .O(N__31282),
            .I(N__31276));
    LocalMux I__5840 (
            .O(N__31279),
            .I(\phase_controller_inst1.tr_time_passed ));
    Odrv4 I__5839 (
            .O(N__31276),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__5838 (
            .O(N__31271),
            .I(N__31262));
    InMux I__5837 (
            .O(N__31270),
            .I(N__31262));
    InMux I__5836 (
            .O(N__31269),
            .I(N__31262));
    LocalMux I__5835 (
            .O(N__31262),
            .I(\phase_controller_inst2.tr_time_passed ));
    CascadeMux I__5834 (
            .O(N__31259),
            .I(\phase_controller_inst2.time_passed_RNI9M3O_cascade_ ));
    CascadeMux I__5833 (
            .O(N__31256),
            .I(N__31249));
    InMux I__5832 (
            .O(N__31255),
            .I(N__31242));
    InMux I__5831 (
            .O(N__31254),
            .I(N__31242));
    InMux I__5830 (
            .O(N__31253),
            .I(N__31242));
    CascadeMux I__5829 (
            .O(N__31252),
            .I(N__31239));
    InMux I__5828 (
            .O(N__31249),
            .I(N__31235));
    LocalMux I__5827 (
            .O(N__31242),
            .I(N__31232));
    InMux I__5826 (
            .O(N__31239),
            .I(N__31229));
    InMux I__5825 (
            .O(N__31238),
            .I(N__31226));
    LocalMux I__5824 (
            .O(N__31235),
            .I(N__31221));
    Span4Mux_v I__5823 (
            .O(N__31232),
            .I(N__31221));
    LocalMux I__5822 (
            .O(N__31229),
            .I(N__31216));
    LocalMux I__5821 (
            .O(N__31226),
            .I(N__31216));
    Odrv4 I__5820 (
            .O(N__31221),
            .I(state_3));
    Odrv4 I__5819 (
            .O(N__31216),
            .I(state_3));
    IoInMux I__5818 (
            .O(N__31211),
            .I(N__31208));
    LocalMux I__5817 (
            .O(N__31208),
            .I(N__31205));
    Span4Mux_s3_v I__5816 (
            .O(N__31205),
            .I(N__31202));
    Sp12to4 I__5815 (
            .O(N__31202),
            .I(N__31199));
    Span12Mux_h I__5814 (
            .O(N__31199),
            .I(N__31196));
    Span12Mux_v I__5813 (
            .O(N__31196),
            .I(N__31191));
    InMux I__5812 (
            .O(N__31195),
            .I(N__31186));
    InMux I__5811 (
            .O(N__31194),
            .I(N__31186));
    Odrv12 I__5810 (
            .O(N__31191),
            .I(s1_phy_c));
    LocalMux I__5809 (
            .O(N__31186),
            .I(s1_phy_c));
    InMux I__5808 (
            .O(N__31181),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__5807 (
            .O(N__31178),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__5806 (
            .O(N__31175),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__5805 (
            .O(N__31172),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__5804 (
            .O(N__31169),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__5803 (
            .O(N__31166),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__5802 (
            .O(N__31163),
            .I(bfn_13_13_0_));
    InMux I__5801 (
            .O(N__31160),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__5800 (
            .O(N__31157),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__5799 (
            .O(N__31154),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ));
    InMux I__5798 (
            .O(N__31151),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__5797 (
            .O(N__31148),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__5796 (
            .O(N__31145),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__5795 (
            .O(N__31142),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__5794 (
            .O(N__31139),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__5793 (
            .O(N__31136),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__5792 (
            .O(N__31133),
            .I(bfn_13_12_0_));
    InMux I__5791 (
            .O(N__31130),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ));
    CascadeMux I__5790 (
            .O(N__31127),
            .I(N__31123));
    InMux I__5789 (
            .O(N__31126),
            .I(N__31120));
    InMux I__5788 (
            .O(N__31123),
            .I(N__31117));
    LocalMux I__5787 (
            .O(N__31120),
            .I(N__31114));
    LocalMux I__5786 (
            .O(N__31117),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ));
    Odrv4 I__5785 (
            .O(N__31114),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ));
    CascadeMux I__5784 (
            .O(N__31109),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6_cascade_ ));
    CascadeMux I__5783 (
            .O(N__31106),
            .I(elapsed_time_ns_1_RNIUKL2M1_0_6_cascade_));
    InMux I__5782 (
            .O(N__31103),
            .I(N__31094));
    InMux I__5781 (
            .O(N__31102),
            .I(N__31094));
    InMux I__5780 (
            .O(N__31101),
            .I(N__31094));
    LocalMux I__5779 (
            .O(N__31094),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2 ));
    CascadeMux I__5778 (
            .O(N__31091),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_ ));
    CascadeMux I__5777 (
            .O(N__31088),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_ ));
    CascadeMux I__5776 (
            .O(N__31085),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19_cascade_ ));
    CascadeMux I__5775 (
            .O(N__31082),
            .I(elapsed_time_ns_1_RNIIJ4DM1_0_19_cascade_));
    InMux I__5774 (
            .O(N__31079),
            .I(N__31075));
    InMux I__5773 (
            .O(N__31078),
            .I(N__31070));
    LocalMux I__5772 (
            .O(N__31075),
            .I(N__31067));
    InMux I__5771 (
            .O(N__31074),
            .I(N__31064));
    InMux I__5770 (
            .O(N__31073),
            .I(N__31061));
    LocalMux I__5769 (
            .O(N__31070),
            .I(N__31056));
    Span12Mux_s9_v I__5768 (
            .O(N__31067),
            .I(N__31056));
    LocalMux I__5767 (
            .O(N__31064),
            .I(N__31053));
    LocalMux I__5766 (
            .O(N__31061),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv12 I__5765 (
            .O(N__31056),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__5764 (
            .O(N__31053),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__5763 (
            .O(N__31046),
            .I(N__31043));
    LocalMux I__5762 (
            .O(N__31043),
            .I(N__31040));
    Span4Mux_s1_v I__5761 (
            .O(N__31040),
            .I(N__31037));
    Odrv4 I__5760 (
            .O(N__31037),
            .I(s2_phy_c));
    IoInMux I__5759 (
            .O(N__31034),
            .I(N__31031));
    LocalMux I__5758 (
            .O(N__31031),
            .I(N__31028));
    Span4Mux_s0_v I__5757 (
            .O(N__31028),
            .I(N__31025));
    Odrv4 I__5756 (
            .O(N__31025),
            .I(\pll_inst.red_c_i ));
    InMux I__5755 (
            .O(N__31022),
            .I(N__31019));
    LocalMux I__5754 (
            .O(N__31019),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1 ));
    InMux I__5753 (
            .O(N__31016),
            .I(N__31012));
    CascadeMux I__5752 (
            .O(N__31015),
            .I(N__31009));
    LocalMux I__5751 (
            .O(N__31012),
            .I(N__31006));
    InMux I__5750 (
            .O(N__31009),
            .I(N__31003));
    Odrv4 I__5749 (
            .O(N__31006),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    LocalMux I__5748 (
            .O(N__31003),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__5747 (
            .O(N__30998),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__5746 (
            .O(N__30995),
            .I(N__30992));
    InMux I__5745 (
            .O(N__30992),
            .I(N__30989));
    LocalMux I__5744 (
            .O(N__30989),
            .I(N__30986));
    Span4Mux_v I__5743 (
            .O(N__30986),
            .I(N__30982));
    InMux I__5742 (
            .O(N__30985),
            .I(N__30979));
    Odrv4 I__5741 (
            .O(N__30982),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    LocalMux I__5740 (
            .O(N__30979),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__5739 (
            .O(N__30974),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__5738 (
            .O(N__30971),
            .I(N__30968));
    InMux I__5737 (
            .O(N__30968),
            .I(N__30965));
    LocalMux I__5736 (
            .O(N__30965),
            .I(N__30962));
    Span4Mux_v I__5735 (
            .O(N__30962),
            .I(N__30958));
    InMux I__5734 (
            .O(N__30961),
            .I(N__30955));
    Odrv4 I__5733 (
            .O(N__30958),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    LocalMux I__5732 (
            .O(N__30955),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__5731 (
            .O(N__30950),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__5730 (
            .O(N__30947),
            .I(N__30944));
    LocalMux I__5729 (
            .O(N__30944),
            .I(N__30941));
    Span4Mux_h I__5728 (
            .O(N__30941),
            .I(N__30937));
    InMux I__5727 (
            .O(N__30940),
            .I(N__30934));
    Odrv4 I__5726 (
            .O(N__30937),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    LocalMux I__5725 (
            .O(N__30934),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__5724 (
            .O(N__30929),
            .I(bfn_12_23_0_));
    InMux I__5723 (
            .O(N__30926),
            .I(N__30923));
    LocalMux I__5722 (
            .O(N__30923),
            .I(N__30920));
    Span4Mux_h I__5721 (
            .O(N__30920),
            .I(N__30916));
    InMux I__5720 (
            .O(N__30919),
            .I(N__30913));
    Odrv4 I__5719 (
            .O(N__30916),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    LocalMux I__5718 (
            .O(N__30913),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__5717 (
            .O(N__30908),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    CascadeMux I__5716 (
            .O(N__30905),
            .I(N__30902));
    InMux I__5715 (
            .O(N__30902),
            .I(N__30899));
    LocalMux I__5714 (
            .O(N__30899),
            .I(N__30896));
    Span4Mux_v I__5713 (
            .O(N__30896),
            .I(N__30892));
    InMux I__5712 (
            .O(N__30895),
            .I(N__30889));
    Odrv4 I__5711 (
            .O(N__30892),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    LocalMux I__5710 (
            .O(N__30889),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__5709 (
            .O(N__30884),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__5708 (
            .O(N__30881),
            .I(N__30878));
    LocalMux I__5707 (
            .O(N__30878),
            .I(N__30875));
    Span4Mux_h I__5706 (
            .O(N__30875),
            .I(N__30871));
    InMux I__5705 (
            .O(N__30874),
            .I(N__30868));
    Odrv4 I__5704 (
            .O(N__30871),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    LocalMux I__5703 (
            .O(N__30868),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__5702 (
            .O(N__30863),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__5701 (
            .O(N__30860),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__5700 (
            .O(N__30857),
            .I(N__30851));
    InMux I__5699 (
            .O(N__30856),
            .I(N__30845));
    InMux I__5698 (
            .O(N__30855),
            .I(N__30845));
    InMux I__5697 (
            .O(N__30854),
            .I(N__30842));
    InMux I__5696 (
            .O(N__30851),
            .I(N__30838));
    InMux I__5695 (
            .O(N__30850),
            .I(N__30835));
    LocalMux I__5694 (
            .O(N__30845),
            .I(N__30830));
    LocalMux I__5693 (
            .O(N__30842),
            .I(N__30830));
    InMux I__5692 (
            .O(N__30841),
            .I(N__30827));
    LocalMux I__5691 (
            .O(N__30838),
            .I(N__30824));
    LocalMux I__5690 (
            .O(N__30835),
            .I(N__30821));
    Span4Mux_h I__5689 (
            .O(N__30830),
            .I(N__30816));
    LocalMux I__5688 (
            .O(N__30827),
            .I(N__30816));
    Span4Mux_v I__5687 (
            .O(N__30824),
            .I(N__30813));
    Span4Mux_v I__5686 (
            .O(N__30821),
            .I(N__30810));
    Span4Mux_v I__5685 (
            .O(N__30816),
            .I(N__30807));
    Odrv4 I__5684 (
            .O(N__30813),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__5683 (
            .O(N__30810),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__5682 (
            .O(N__30807),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__5681 (
            .O(N__30800),
            .I(N__30796));
    CascadeMux I__5680 (
            .O(N__30799),
            .I(N__30792));
    LocalMux I__5679 (
            .O(N__30796),
            .I(N__30787));
    InMux I__5678 (
            .O(N__30795),
            .I(N__30782));
    InMux I__5677 (
            .O(N__30792),
            .I(N__30782));
    InMux I__5676 (
            .O(N__30791),
            .I(N__30777));
    InMux I__5675 (
            .O(N__30790),
            .I(N__30777));
    Span4Mux_v I__5674 (
            .O(N__30787),
            .I(N__30774));
    LocalMux I__5673 (
            .O(N__30782),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__5672 (
            .O(N__30777),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__5671 (
            .O(N__30774),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    CascadeMux I__5670 (
            .O(N__30767),
            .I(N__30764));
    InMux I__5669 (
            .O(N__30764),
            .I(N__30760));
    CascadeMux I__5668 (
            .O(N__30763),
            .I(N__30757));
    LocalMux I__5667 (
            .O(N__30760),
            .I(N__30754));
    InMux I__5666 (
            .O(N__30757),
            .I(N__30751));
    Span4Mux_h I__5665 (
            .O(N__30754),
            .I(N__30747));
    LocalMux I__5664 (
            .O(N__30751),
            .I(N__30744));
    InMux I__5663 (
            .O(N__30750),
            .I(N__30741));
    Odrv4 I__5662 (
            .O(N__30747),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    Odrv4 I__5661 (
            .O(N__30744),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    LocalMux I__5660 (
            .O(N__30741),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    InMux I__5659 (
            .O(N__30734),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__5658 (
            .O(N__30731),
            .I(N__30728));
    LocalMux I__5657 (
            .O(N__30728),
            .I(N__30724));
    InMux I__5656 (
            .O(N__30727),
            .I(N__30721));
    Span4Mux_h I__5655 (
            .O(N__30724),
            .I(N__30717));
    LocalMux I__5654 (
            .O(N__30721),
            .I(N__30714));
    InMux I__5653 (
            .O(N__30720),
            .I(N__30711));
    Odrv4 I__5652 (
            .O(N__30717),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    Odrv4 I__5651 (
            .O(N__30714),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    LocalMux I__5650 (
            .O(N__30711),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    InMux I__5649 (
            .O(N__30704),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__5648 (
            .O(N__30701),
            .I(N__30698));
    InMux I__5647 (
            .O(N__30698),
            .I(N__30695));
    LocalMux I__5646 (
            .O(N__30695),
            .I(N__30692));
    Span4Mux_h I__5645 (
            .O(N__30692),
            .I(N__30688));
    InMux I__5644 (
            .O(N__30691),
            .I(N__30685));
    Span4Mux_h I__5643 (
            .O(N__30688),
            .I(N__30681));
    LocalMux I__5642 (
            .O(N__30685),
            .I(N__30678));
    InMux I__5641 (
            .O(N__30684),
            .I(N__30675));
    Odrv4 I__5640 (
            .O(N__30681),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    Odrv4 I__5639 (
            .O(N__30678),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    LocalMux I__5638 (
            .O(N__30675),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__5637 (
            .O(N__30668),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__5636 (
            .O(N__30665),
            .I(N__30662));
    InMux I__5635 (
            .O(N__30662),
            .I(N__30658));
    CascadeMux I__5634 (
            .O(N__30661),
            .I(N__30654));
    LocalMux I__5633 (
            .O(N__30658),
            .I(N__30651));
    InMux I__5632 (
            .O(N__30657),
            .I(N__30648));
    InMux I__5631 (
            .O(N__30654),
            .I(N__30645));
    Span4Mux_h I__5630 (
            .O(N__30651),
            .I(N__30642));
    LocalMux I__5629 (
            .O(N__30648),
            .I(N__30637));
    LocalMux I__5628 (
            .O(N__30645),
            .I(N__30637));
    Odrv4 I__5627 (
            .O(N__30642),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    Odrv4 I__5626 (
            .O(N__30637),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    InMux I__5625 (
            .O(N__30632),
            .I(bfn_12_22_0_));
    InMux I__5624 (
            .O(N__30629),
            .I(N__30626));
    LocalMux I__5623 (
            .O(N__30626),
            .I(N__30623));
    Span4Mux_h I__5622 (
            .O(N__30623),
            .I(N__30619));
    InMux I__5621 (
            .O(N__30622),
            .I(N__30616));
    Odrv4 I__5620 (
            .O(N__30619),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    LocalMux I__5619 (
            .O(N__30616),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__5618 (
            .O(N__30611),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__5617 (
            .O(N__30608),
            .I(N__30605));
    InMux I__5616 (
            .O(N__30605),
            .I(N__30602));
    LocalMux I__5615 (
            .O(N__30602),
            .I(N__30599));
    Span4Mux_h I__5614 (
            .O(N__30599),
            .I(N__30595));
    InMux I__5613 (
            .O(N__30598),
            .I(N__30592));
    Odrv4 I__5612 (
            .O(N__30595),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    LocalMux I__5611 (
            .O(N__30592),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__5610 (
            .O(N__30587),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__5609 (
            .O(N__30584),
            .I(N__30581));
    LocalMux I__5608 (
            .O(N__30581),
            .I(N__30577));
    InMux I__5607 (
            .O(N__30580),
            .I(N__30574));
    Odrv4 I__5606 (
            .O(N__30577),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    LocalMux I__5605 (
            .O(N__30574),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__5604 (
            .O(N__30569),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__5603 (
            .O(N__30566),
            .I(N__30563));
    InMux I__5602 (
            .O(N__30563),
            .I(N__30560));
    LocalMux I__5601 (
            .O(N__30560),
            .I(N__30556));
    CascadeMux I__5600 (
            .O(N__30559),
            .I(N__30553));
    Span4Mux_h I__5599 (
            .O(N__30556),
            .I(N__30550));
    InMux I__5598 (
            .O(N__30553),
            .I(N__30547));
    Odrv4 I__5597 (
            .O(N__30550),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    LocalMux I__5596 (
            .O(N__30547),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__5595 (
            .O(N__30542),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__5594 (
            .O(N__30539),
            .I(N__30536));
    InMux I__5593 (
            .O(N__30536),
            .I(N__30533));
    LocalMux I__5592 (
            .O(N__30533),
            .I(N__30530));
    Span4Mux_v I__5591 (
            .O(N__30530),
            .I(N__30525));
    InMux I__5590 (
            .O(N__30529),
            .I(N__30520));
    InMux I__5589 (
            .O(N__30528),
            .I(N__30520));
    Odrv4 I__5588 (
            .O(N__30525),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    LocalMux I__5587 (
            .O(N__30520),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__5586 (
            .O(N__30515),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__5585 (
            .O(N__30512),
            .I(N__30509));
    InMux I__5584 (
            .O(N__30509),
            .I(N__30506));
    LocalMux I__5583 (
            .O(N__30506),
            .I(N__30503));
    Span4Mux_v I__5582 (
            .O(N__30503),
            .I(N__30498));
    InMux I__5581 (
            .O(N__30502),
            .I(N__30493));
    InMux I__5580 (
            .O(N__30501),
            .I(N__30493));
    Odrv4 I__5579 (
            .O(N__30498),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    LocalMux I__5578 (
            .O(N__30493),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__5577 (
            .O(N__30488),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__5576 (
            .O(N__30485),
            .I(N__30482));
    InMux I__5575 (
            .O(N__30482),
            .I(N__30479));
    LocalMux I__5574 (
            .O(N__30479),
            .I(N__30476));
    Span4Mux_v I__5573 (
            .O(N__30476),
            .I(N__30473));
    Span4Mux_h I__5572 (
            .O(N__30473),
            .I(N__30467));
    InMux I__5571 (
            .O(N__30472),
            .I(N__30464));
    InMux I__5570 (
            .O(N__30471),
            .I(N__30461));
    InMux I__5569 (
            .O(N__30470),
            .I(N__30458));
    Odrv4 I__5568 (
            .O(N__30467),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ));
    LocalMux I__5567 (
            .O(N__30464),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ));
    LocalMux I__5566 (
            .O(N__30461),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ));
    LocalMux I__5565 (
            .O(N__30458),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ));
    InMux I__5564 (
            .O(N__30449),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__5563 (
            .O(N__30446),
            .I(N__30443));
    InMux I__5562 (
            .O(N__30443),
            .I(N__30440));
    LocalMux I__5561 (
            .O(N__30440),
            .I(N__30436));
    CascadeMux I__5560 (
            .O(N__30439),
            .I(N__30433));
    Span4Mux_v I__5559 (
            .O(N__30436),
            .I(N__30430));
    InMux I__5558 (
            .O(N__30433),
            .I(N__30427));
    Odrv4 I__5557 (
            .O(N__30430),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    LocalMux I__5556 (
            .O(N__30427),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__5555 (
            .O(N__30422),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__5554 (
            .O(N__30419),
            .I(N__30416));
    InMux I__5553 (
            .O(N__30416),
            .I(N__30413));
    LocalMux I__5552 (
            .O(N__30413),
            .I(N__30410));
    Span4Mux_h I__5551 (
            .O(N__30410),
            .I(N__30406));
    InMux I__5550 (
            .O(N__30409),
            .I(N__30403));
    Odrv4 I__5549 (
            .O(N__30406),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    LocalMux I__5548 (
            .O(N__30403),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__5547 (
            .O(N__30398),
            .I(bfn_12_21_0_));
    CascadeMux I__5546 (
            .O(N__30395),
            .I(N__30392));
    InMux I__5545 (
            .O(N__30392),
            .I(N__30389));
    LocalMux I__5544 (
            .O(N__30389),
            .I(N__30386));
    Span4Mux_v I__5543 (
            .O(N__30386),
            .I(N__30382));
    InMux I__5542 (
            .O(N__30385),
            .I(N__30379));
    Odrv4 I__5541 (
            .O(N__30382),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    LocalMux I__5540 (
            .O(N__30379),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__5539 (
            .O(N__30374),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__5538 (
            .O(N__30371),
            .I(N__30368));
    InMux I__5537 (
            .O(N__30368),
            .I(N__30365));
    LocalMux I__5536 (
            .O(N__30365),
            .I(N__30362));
    Span4Mux_h I__5535 (
            .O(N__30362),
            .I(N__30358));
    InMux I__5534 (
            .O(N__30361),
            .I(N__30355));
    Odrv4 I__5533 (
            .O(N__30358),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__5532 (
            .O(N__30355),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__5531 (
            .O(N__30350),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__5530 (
            .O(N__30347),
            .I(N__30344));
    InMux I__5529 (
            .O(N__30344),
            .I(N__30341));
    LocalMux I__5528 (
            .O(N__30341),
            .I(N__30337));
    InMux I__5527 (
            .O(N__30340),
            .I(N__30332));
    Span4Mux_v I__5526 (
            .O(N__30337),
            .I(N__30329));
    InMux I__5525 (
            .O(N__30336),
            .I(N__30326));
    InMux I__5524 (
            .O(N__30335),
            .I(N__30323));
    LocalMux I__5523 (
            .O(N__30332),
            .I(N__30320));
    Span4Mux_h I__5522 (
            .O(N__30329),
            .I(N__30315));
    LocalMux I__5521 (
            .O(N__30326),
            .I(N__30315));
    LocalMux I__5520 (
            .O(N__30323),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto14 ));
    Odrv4 I__5519 (
            .O(N__30320),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto14 ));
    Odrv4 I__5518 (
            .O(N__30315),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto14 ));
    InMux I__5517 (
            .O(N__30308),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__5516 (
            .O(N__30305),
            .I(N__30302));
    InMux I__5515 (
            .O(N__30302),
            .I(N__30297));
    InMux I__5514 (
            .O(N__30301),
            .I(N__30294));
    InMux I__5513 (
            .O(N__30300),
            .I(N__30291));
    LocalMux I__5512 (
            .O(N__30297),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto15 ));
    LocalMux I__5511 (
            .O(N__30294),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto15 ));
    LocalMux I__5510 (
            .O(N__30291),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto15 ));
    InMux I__5509 (
            .O(N__30284),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__5508 (
            .O(N__30281),
            .I(N__30277));
    InMux I__5507 (
            .O(N__30280),
            .I(N__30274));
    LocalMux I__5506 (
            .O(N__30277),
            .I(N__30271));
    LocalMux I__5505 (
            .O(N__30274),
            .I(N__30267));
    Span4Mux_h I__5504 (
            .O(N__30271),
            .I(N__30260));
    InMux I__5503 (
            .O(N__30270),
            .I(N__30257));
    Span4Mux_h I__5502 (
            .O(N__30267),
            .I(N__30254));
    InMux I__5501 (
            .O(N__30266),
            .I(N__30247));
    InMux I__5500 (
            .O(N__30265),
            .I(N__30247));
    InMux I__5499 (
            .O(N__30264),
            .I(N__30247));
    InMux I__5498 (
            .O(N__30263),
            .I(N__30244));
    Odrv4 I__5497 (
            .O(N__30260),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    LocalMux I__5496 (
            .O(N__30257),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    Odrv4 I__5495 (
            .O(N__30254),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    LocalMux I__5494 (
            .O(N__30247),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    LocalMux I__5493 (
            .O(N__30244),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ));
    InMux I__5492 (
            .O(N__30233),
            .I(N__30228));
    InMux I__5491 (
            .O(N__30232),
            .I(N__30225));
    CascadeMux I__5490 (
            .O(N__30231),
            .I(N__30222));
    LocalMux I__5489 (
            .O(N__30228),
            .I(N__30217));
    LocalMux I__5488 (
            .O(N__30225),
            .I(N__30217));
    InMux I__5487 (
            .O(N__30222),
            .I(N__30214));
    Span4Mux_h I__5486 (
            .O(N__30217),
            .I(N__30211));
    LocalMux I__5485 (
            .O(N__30214),
            .I(elapsed_time_ns_1_RNIIU2KD1_0_6));
    Odrv4 I__5484 (
            .O(N__30211),
            .I(elapsed_time_ns_1_RNIIU2KD1_0_6));
    InMux I__5483 (
            .O(N__30206),
            .I(N__30197));
    InMux I__5482 (
            .O(N__30205),
            .I(N__30194));
    InMux I__5481 (
            .O(N__30204),
            .I(N__30187));
    InMux I__5480 (
            .O(N__30203),
            .I(N__30187));
    InMux I__5479 (
            .O(N__30202),
            .I(N__30187));
    InMux I__5478 (
            .O(N__30201),
            .I(N__30182));
    InMux I__5477 (
            .O(N__30200),
            .I(N__30179));
    LocalMux I__5476 (
            .O(N__30197),
            .I(N__30174));
    LocalMux I__5475 (
            .O(N__30194),
            .I(N__30174));
    LocalMux I__5474 (
            .O(N__30187),
            .I(N__30171));
    InMux I__5473 (
            .O(N__30186),
            .I(N__30168));
    InMux I__5472 (
            .O(N__30185),
            .I(N__30165));
    LocalMux I__5471 (
            .O(N__30182),
            .I(N__30162));
    LocalMux I__5470 (
            .O(N__30179),
            .I(N__30157));
    Span4Mux_v I__5469 (
            .O(N__30174),
            .I(N__30157));
    Odrv12 I__5468 (
            .O(N__30171),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5 ));
    LocalMux I__5467 (
            .O(N__30168),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5 ));
    LocalMux I__5466 (
            .O(N__30165),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5 ));
    Odrv4 I__5465 (
            .O(N__30162),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5 ));
    Odrv4 I__5464 (
            .O(N__30157),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5 ));
    CascadeMux I__5463 (
            .O(N__30146),
            .I(elapsed_time_ns_1_RNIIU2KD1_0_6_cascade_));
    InMux I__5462 (
            .O(N__30143),
            .I(N__30140));
    LocalMux I__5461 (
            .O(N__30140),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6 ));
    InMux I__5460 (
            .O(N__30137),
            .I(N__30134));
    LocalMux I__5459 (
            .O(N__30134),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6 ));
    InMux I__5458 (
            .O(N__30131),
            .I(N__30125));
    InMux I__5457 (
            .O(N__30130),
            .I(N__30125));
    LocalMux I__5456 (
            .O(N__30125),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4 ));
    InMux I__5455 (
            .O(N__30122),
            .I(N__30117));
    InMux I__5454 (
            .O(N__30121),
            .I(N__30112));
    InMux I__5453 (
            .O(N__30120),
            .I(N__30112));
    LocalMux I__5452 (
            .O(N__30117),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    LocalMux I__5451 (
            .O(N__30112),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    CascadeMux I__5450 (
            .O(N__30107),
            .I(N__30104));
    InMux I__5449 (
            .O(N__30104),
            .I(N__30101));
    LocalMux I__5448 (
            .O(N__30101),
            .I(N__30098));
    Span4Mux_v I__5447 (
            .O(N__30098),
            .I(N__30094));
    InMux I__5446 (
            .O(N__30097),
            .I(N__30091));
    Odrv4 I__5445 (
            .O(N__30094),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    LocalMux I__5444 (
            .O(N__30091),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__5443 (
            .O(N__30086),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__5442 (
            .O(N__30083),
            .I(N__30080));
    InMux I__5441 (
            .O(N__30080),
            .I(N__30077));
    LocalMux I__5440 (
            .O(N__30077),
            .I(N__30074));
    Span4Mux_h I__5439 (
            .O(N__30074),
            .I(N__30070));
    InMux I__5438 (
            .O(N__30073),
            .I(N__30067));
    Odrv4 I__5437 (
            .O(N__30070),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    LocalMux I__5436 (
            .O(N__30067),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__5435 (
            .O(N__30062),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__5434 (
            .O(N__30059),
            .I(N__30052));
    InMux I__5433 (
            .O(N__30058),
            .I(N__30052));
    InMux I__5432 (
            .O(N__30057),
            .I(N__30049));
    LocalMux I__5431 (
            .O(N__30052),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto6 ));
    LocalMux I__5430 (
            .O(N__30049),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lto6 ));
    InMux I__5429 (
            .O(N__30044),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__5428 (
            .O(N__30041),
            .I(N__30038));
    LocalMux I__5427 (
            .O(N__30038),
            .I(N__30035));
    Span4Mux_h I__5426 (
            .O(N__30035),
            .I(N__30032));
    Odrv4 I__5425 (
            .O(N__30032),
            .I(\phase_controller_inst1.stoper_hc.un6_running_17 ));
    InMux I__5424 (
            .O(N__30029),
            .I(N__30025));
    InMux I__5423 (
            .O(N__30028),
            .I(N__30022));
    LocalMux I__5422 (
            .O(N__30025),
            .I(N__30019));
    LocalMux I__5421 (
            .O(N__30022),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv12 I__5420 (
            .O(N__30019),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__5419 (
            .O(N__30014),
            .I(N__30011));
    InMux I__5418 (
            .O(N__30011),
            .I(N__30008));
    LocalMux I__5417 (
            .O(N__30008),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ));
    InMux I__5416 (
            .O(N__30005),
            .I(N__30002));
    LocalMux I__5415 (
            .O(N__30002),
            .I(N__29999));
    Span4Mux_v I__5414 (
            .O(N__29999),
            .I(N__29996));
    Odrv4 I__5413 (
            .O(N__29996),
            .I(\phase_controller_inst1.stoper_hc.un6_running_18 ));
    InMux I__5412 (
            .O(N__29993),
            .I(N__29989));
    InMux I__5411 (
            .O(N__29992),
            .I(N__29986));
    LocalMux I__5410 (
            .O(N__29989),
            .I(N__29983));
    LocalMux I__5409 (
            .O(N__29986),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv12 I__5408 (
            .O(N__29983),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__5407 (
            .O(N__29978),
            .I(N__29975));
    InMux I__5406 (
            .O(N__29975),
            .I(N__29972));
    LocalMux I__5405 (
            .O(N__29972),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ));
    InMux I__5404 (
            .O(N__29969),
            .I(N__29966));
    LocalMux I__5403 (
            .O(N__29966),
            .I(N__29963));
    Span4Mux_v I__5402 (
            .O(N__29963),
            .I(N__29960));
    Odrv4 I__5401 (
            .O(N__29960),
            .I(\phase_controller_inst1.stoper_hc.un6_running_19 ));
    InMux I__5400 (
            .O(N__29957),
            .I(N__29953));
    InMux I__5399 (
            .O(N__29956),
            .I(N__29950));
    LocalMux I__5398 (
            .O(N__29953),
            .I(N__29947));
    LocalMux I__5397 (
            .O(N__29950),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__5396 (
            .O(N__29947),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    CascadeMux I__5395 (
            .O(N__29942),
            .I(N__29939));
    InMux I__5394 (
            .O(N__29939),
            .I(N__29936));
    LocalMux I__5393 (
            .O(N__29936),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ));
    InMux I__5392 (
            .O(N__29933),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_19 ));
    InMux I__5391 (
            .O(N__29930),
            .I(N__29926));
    InMux I__5390 (
            .O(N__29929),
            .I(N__29922));
    LocalMux I__5389 (
            .O(N__29926),
            .I(N__29919));
    InMux I__5388 (
            .O(N__29925),
            .I(N__29916));
    LocalMux I__5387 (
            .O(N__29922),
            .I(N__29913));
    Span4Mux_h I__5386 (
            .O(N__29919),
            .I(N__29910));
    LocalMux I__5385 (
            .O(N__29916),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1 ));
    Odrv4 I__5384 (
            .O(N__29913),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1 ));
    Odrv4 I__5383 (
            .O(N__29910),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1 ));
    CascadeMux I__5382 (
            .O(N__29903),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2_cascade_ ));
    InMux I__5381 (
            .O(N__29900),
            .I(N__29897));
    LocalMux I__5380 (
            .O(N__29897),
            .I(N__29893));
    InMux I__5379 (
            .O(N__29896),
            .I(N__29890));
    Span4Mux_v I__5378 (
            .O(N__29893),
            .I(N__29887));
    LocalMux I__5377 (
            .O(N__29890),
            .I(N__29884));
    Odrv4 I__5376 (
            .O(N__29887),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15 ));
    Odrv4 I__5375 (
            .O(N__29884),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15 ));
    CascadeMux I__5374 (
            .O(N__29879),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5_cascade_ ));
    InMux I__5373 (
            .O(N__29876),
            .I(N__29871));
    InMux I__5372 (
            .O(N__29875),
            .I(N__29865));
    InMux I__5371 (
            .O(N__29874),
            .I(N__29865));
    LocalMux I__5370 (
            .O(N__29871),
            .I(N__29862));
    InMux I__5369 (
            .O(N__29870),
            .I(N__29859));
    LocalMux I__5368 (
            .O(N__29865),
            .I(N__29856));
    Span4Mux_h I__5367 (
            .O(N__29862),
            .I(N__29853));
    LocalMux I__5366 (
            .O(N__29859),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17 ));
    Odrv4 I__5365 (
            .O(N__29856),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17 ));
    Odrv4 I__5364 (
            .O(N__29853),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17 ));
    InMux I__5363 (
            .O(N__29846),
            .I(N__29843));
    LocalMux I__5362 (
            .O(N__29843),
            .I(N__29840));
    Span4Mux_h I__5361 (
            .O(N__29840),
            .I(N__29837));
    Odrv4 I__5360 (
            .O(N__29837),
            .I(\phase_controller_inst1.stoper_hc.un6_running_9 ));
    InMux I__5359 (
            .O(N__29834),
            .I(N__29830));
    InMux I__5358 (
            .O(N__29833),
            .I(N__29827));
    LocalMux I__5357 (
            .O(N__29830),
            .I(N__29824));
    LocalMux I__5356 (
            .O(N__29827),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv12 I__5355 (
            .O(N__29824),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__5354 (
            .O(N__29819),
            .I(N__29816));
    InMux I__5353 (
            .O(N__29816),
            .I(N__29813));
    LocalMux I__5352 (
            .O(N__29813),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__5351 (
            .O(N__29810),
            .I(N__29807));
    InMux I__5350 (
            .O(N__29807),
            .I(N__29804));
    LocalMux I__5349 (
            .O(N__29804),
            .I(N__29801));
    Span4Mux_h I__5348 (
            .O(N__29801),
            .I(N__29798));
    Odrv4 I__5347 (
            .O(N__29798),
            .I(\phase_controller_inst1.stoper_hc.un6_running_10 ));
    InMux I__5346 (
            .O(N__29795),
            .I(N__29791));
    InMux I__5345 (
            .O(N__29794),
            .I(N__29788));
    LocalMux I__5344 (
            .O(N__29791),
            .I(N__29785));
    LocalMux I__5343 (
            .O(N__29788),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv12 I__5342 (
            .O(N__29785),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__5341 (
            .O(N__29780),
            .I(N__29777));
    LocalMux I__5340 (
            .O(N__29777),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__5339 (
            .O(N__29774),
            .I(N__29771));
    InMux I__5338 (
            .O(N__29771),
            .I(N__29768));
    LocalMux I__5337 (
            .O(N__29768),
            .I(\phase_controller_inst1.stoper_hc.un6_running_11 ));
    InMux I__5336 (
            .O(N__29765),
            .I(N__29761));
    InMux I__5335 (
            .O(N__29764),
            .I(N__29758));
    LocalMux I__5334 (
            .O(N__29761),
            .I(N__29755));
    LocalMux I__5333 (
            .O(N__29758),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__5332 (
            .O(N__29755),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__5331 (
            .O(N__29750),
            .I(N__29747));
    LocalMux I__5330 (
            .O(N__29747),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__5329 (
            .O(N__29744),
            .I(N__29741));
    InMux I__5328 (
            .O(N__29741),
            .I(N__29738));
    LocalMux I__5327 (
            .O(N__29738),
            .I(\phase_controller_inst1.stoper_hc.un6_running_12 ));
    InMux I__5326 (
            .O(N__29735),
            .I(N__29731));
    InMux I__5325 (
            .O(N__29734),
            .I(N__29728));
    LocalMux I__5324 (
            .O(N__29731),
            .I(N__29725));
    LocalMux I__5323 (
            .O(N__29728),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__5322 (
            .O(N__29725),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__5321 (
            .O(N__29720),
            .I(N__29717));
    LocalMux I__5320 (
            .O(N__29717),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__5319 (
            .O(N__29714),
            .I(N__29711));
    InMux I__5318 (
            .O(N__29711),
            .I(N__29708));
    LocalMux I__5317 (
            .O(N__29708),
            .I(\phase_controller_inst1.stoper_hc.un6_running_13 ));
    InMux I__5316 (
            .O(N__29705),
            .I(N__29701));
    InMux I__5315 (
            .O(N__29704),
            .I(N__29698));
    LocalMux I__5314 (
            .O(N__29701),
            .I(N__29695));
    LocalMux I__5313 (
            .O(N__29698),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__5312 (
            .O(N__29695),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__5311 (
            .O(N__29690),
            .I(N__29687));
    LocalMux I__5310 (
            .O(N__29687),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__5309 (
            .O(N__29684),
            .I(N__29681));
    LocalMux I__5308 (
            .O(N__29681),
            .I(N__29678));
    Span12Mux_h I__5307 (
            .O(N__29678),
            .I(N__29675));
    Odrv12 I__5306 (
            .O(N__29675),
            .I(\phase_controller_inst1.stoper_hc.un6_running_14 ));
    InMux I__5305 (
            .O(N__29672),
            .I(N__29668));
    InMux I__5304 (
            .O(N__29671),
            .I(N__29665));
    LocalMux I__5303 (
            .O(N__29668),
            .I(N__29662));
    LocalMux I__5302 (
            .O(N__29665),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__5301 (
            .O(N__29662),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__5300 (
            .O(N__29657),
            .I(N__29654));
    InMux I__5299 (
            .O(N__29654),
            .I(N__29651));
    LocalMux I__5298 (
            .O(N__29651),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__5297 (
            .O(N__29648),
            .I(N__29644));
    InMux I__5296 (
            .O(N__29647),
            .I(N__29641));
    LocalMux I__5295 (
            .O(N__29644),
            .I(N__29638));
    LocalMux I__5294 (
            .O(N__29641),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__5293 (
            .O(N__29638),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__5292 (
            .O(N__29633),
            .I(N__29630));
    LocalMux I__5291 (
            .O(N__29630),
            .I(\phase_controller_inst1.stoper_hc.un6_running_15 ));
    CascadeMux I__5290 (
            .O(N__29627),
            .I(N__29624));
    InMux I__5289 (
            .O(N__29624),
            .I(N__29621));
    LocalMux I__5288 (
            .O(N__29621),
            .I(N__29618));
    Odrv4 I__5287 (
            .O(N__29618),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__5286 (
            .O(N__29615),
            .I(N__29612));
    LocalMux I__5285 (
            .O(N__29612),
            .I(N__29609));
    Span12Mux_v I__5284 (
            .O(N__29609),
            .I(N__29606));
    Odrv12 I__5283 (
            .O(N__29606),
            .I(\phase_controller_inst1.stoper_hc.un6_running_16 ));
    InMux I__5282 (
            .O(N__29603),
            .I(N__29599));
    InMux I__5281 (
            .O(N__29602),
            .I(N__29596));
    LocalMux I__5280 (
            .O(N__29599),
            .I(N__29593));
    LocalMux I__5279 (
            .O(N__29596),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__5278 (
            .O(N__29593),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__5277 (
            .O(N__29588),
            .I(N__29585));
    InMux I__5276 (
            .O(N__29585),
            .I(N__29582));
    LocalMux I__5275 (
            .O(N__29582),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ));
    InMux I__5274 (
            .O(N__29579),
            .I(N__29576));
    LocalMux I__5273 (
            .O(N__29576),
            .I(N__29573));
    Odrv4 I__5272 (
            .O(N__29573),
            .I(\phase_controller_inst1.stoper_hc.un6_running_2 ));
    InMux I__5271 (
            .O(N__29570),
            .I(N__29567));
    LocalMux I__5270 (
            .O(N__29567),
            .I(N__29563));
    InMux I__5269 (
            .O(N__29566),
            .I(N__29560));
    Span4Mux_v I__5268 (
            .O(N__29563),
            .I(N__29557));
    LocalMux I__5267 (
            .O(N__29560),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__5266 (
            .O(N__29557),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__5265 (
            .O(N__29552),
            .I(N__29549));
    InMux I__5264 (
            .O(N__29549),
            .I(N__29546));
    LocalMux I__5263 (
            .O(N__29546),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__5262 (
            .O(N__29543),
            .I(N__29540));
    LocalMux I__5261 (
            .O(N__29540),
            .I(\phase_controller_inst1.stoper_hc.un6_running_3 ));
    CascadeMux I__5260 (
            .O(N__29537),
            .I(N__29533));
    InMux I__5259 (
            .O(N__29536),
            .I(N__29530));
    InMux I__5258 (
            .O(N__29533),
            .I(N__29527));
    LocalMux I__5257 (
            .O(N__29530),
            .I(N__29524));
    LocalMux I__5256 (
            .O(N__29527),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__5255 (
            .O(N__29524),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__5254 (
            .O(N__29519),
            .I(N__29516));
    InMux I__5253 (
            .O(N__29516),
            .I(N__29513));
    LocalMux I__5252 (
            .O(N__29513),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__5251 (
            .O(N__29510),
            .I(N__29506));
    InMux I__5250 (
            .O(N__29509),
            .I(N__29503));
    LocalMux I__5249 (
            .O(N__29506),
            .I(N__29500));
    LocalMux I__5248 (
            .O(N__29503),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv4 I__5247 (
            .O(N__29500),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__5246 (
            .O(N__29495),
            .I(N__29492));
    LocalMux I__5245 (
            .O(N__29492),
            .I(N__29489));
    Odrv4 I__5244 (
            .O(N__29489),
            .I(\phase_controller_inst1.stoper_hc.un6_running_4 ));
    CascadeMux I__5243 (
            .O(N__29486),
            .I(N__29483));
    InMux I__5242 (
            .O(N__29483),
            .I(N__29480));
    LocalMux I__5241 (
            .O(N__29480),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__5240 (
            .O(N__29477),
            .I(N__29474));
    LocalMux I__5239 (
            .O(N__29474),
            .I(N__29471));
    Odrv4 I__5238 (
            .O(N__29471),
            .I(\phase_controller_inst1.stoper_hc.un6_running_5 ));
    InMux I__5237 (
            .O(N__29468),
            .I(N__29464));
    InMux I__5236 (
            .O(N__29467),
            .I(N__29461));
    LocalMux I__5235 (
            .O(N__29464),
            .I(N__29458));
    LocalMux I__5234 (
            .O(N__29461),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv4 I__5233 (
            .O(N__29458),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__5232 (
            .O(N__29453),
            .I(N__29450));
    InMux I__5231 (
            .O(N__29450),
            .I(N__29447));
    LocalMux I__5230 (
            .O(N__29447),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__5229 (
            .O(N__29444),
            .I(N__29441));
    LocalMux I__5228 (
            .O(N__29441),
            .I(N__29438));
    Odrv4 I__5227 (
            .O(N__29438),
            .I(\phase_controller_inst1.stoper_hc.un6_running_6 ));
    InMux I__5226 (
            .O(N__29435),
            .I(N__29431));
    InMux I__5225 (
            .O(N__29434),
            .I(N__29428));
    LocalMux I__5224 (
            .O(N__29431),
            .I(N__29425));
    LocalMux I__5223 (
            .O(N__29428),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv4 I__5222 (
            .O(N__29425),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__5221 (
            .O(N__29420),
            .I(N__29417));
    InMux I__5220 (
            .O(N__29417),
            .I(N__29414));
    LocalMux I__5219 (
            .O(N__29414),
            .I(N__29411));
    Odrv4 I__5218 (
            .O(N__29411),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__5217 (
            .O(N__29408),
            .I(N__29404));
    InMux I__5216 (
            .O(N__29407),
            .I(N__29401));
    LocalMux I__5215 (
            .O(N__29404),
            .I(N__29398));
    LocalMux I__5214 (
            .O(N__29401),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv4 I__5213 (
            .O(N__29398),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__5212 (
            .O(N__29393),
            .I(N__29390));
    InMux I__5211 (
            .O(N__29390),
            .I(N__29387));
    LocalMux I__5210 (
            .O(N__29387),
            .I(\phase_controller_inst1.stoper_hc.un6_running_7 ));
    InMux I__5209 (
            .O(N__29384),
            .I(N__29381));
    LocalMux I__5208 (
            .O(N__29381),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    CascadeMux I__5207 (
            .O(N__29378),
            .I(N__29375));
    InMux I__5206 (
            .O(N__29375),
            .I(N__29372));
    LocalMux I__5205 (
            .O(N__29372),
            .I(\phase_controller_inst1.stoper_hc.un6_running_8 ));
    InMux I__5204 (
            .O(N__29369),
            .I(N__29365));
    InMux I__5203 (
            .O(N__29368),
            .I(N__29362));
    LocalMux I__5202 (
            .O(N__29365),
            .I(N__29359));
    LocalMux I__5201 (
            .O(N__29362),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__5200 (
            .O(N__29359),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__5199 (
            .O(N__29354),
            .I(N__29351));
    LocalMux I__5198 (
            .O(N__29351),
            .I(N__29348));
    Odrv4 I__5197 (
            .O(N__29348),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__5196 (
            .O(N__29345),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__5195 (
            .O(N__29342),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__5194 (
            .O(N__29339),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__5193 (
            .O(N__29336),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__5192 (
            .O(N__29333),
            .I(bfn_12_15_0_));
    InMux I__5191 (
            .O(N__29330),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__5190 (
            .O(N__29327),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__5189 (
            .O(N__29324),
            .I(N__29321));
    LocalMux I__5188 (
            .O(N__29321),
            .I(N__29317));
    InMux I__5187 (
            .O(N__29320),
            .I(N__29314));
    Odrv4 I__5186 (
            .O(N__29317),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__5185 (
            .O(N__29314),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    CEMux I__5184 (
            .O(N__29309),
            .I(N__29305));
    CEMux I__5183 (
            .O(N__29308),
            .I(N__29301));
    LocalMux I__5182 (
            .O(N__29305),
            .I(N__29294));
    CEMux I__5181 (
            .O(N__29304),
            .I(N__29291));
    LocalMux I__5180 (
            .O(N__29301),
            .I(N__29288));
    InMux I__5179 (
            .O(N__29300),
            .I(N__29268));
    InMux I__5178 (
            .O(N__29299),
            .I(N__29268));
    InMux I__5177 (
            .O(N__29298),
            .I(N__29263));
    InMux I__5176 (
            .O(N__29297),
            .I(N__29263));
    Span4Mux_v I__5175 (
            .O(N__29294),
            .I(N__29258));
    LocalMux I__5174 (
            .O(N__29291),
            .I(N__29258));
    Span4Mux_v I__5173 (
            .O(N__29288),
            .I(N__29255));
    InMux I__5172 (
            .O(N__29287),
            .I(N__29246));
    InMux I__5171 (
            .O(N__29286),
            .I(N__29246));
    InMux I__5170 (
            .O(N__29285),
            .I(N__29246));
    InMux I__5169 (
            .O(N__29284),
            .I(N__29246));
    InMux I__5168 (
            .O(N__29283),
            .I(N__29237));
    InMux I__5167 (
            .O(N__29282),
            .I(N__29237));
    InMux I__5166 (
            .O(N__29281),
            .I(N__29237));
    InMux I__5165 (
            .O(N__29280),
            .I(N__29237));
    InMux I__5164 (
            .O(N__29279),
            .I(N__29230));
    InMux I__5163 (
            .O(N__29278),
            .I(N__29230));
    InMux I__5162 (
            .O(N__29277),
            .I(N__29230));
    InMux I__5161 (
            .O(N__29276),
            .I(N__29221));
    InMux I__5160 (
            .O(N__29275),
            .I(N__29221));
    InMux I__5159 (
            .O(N__29274),
            .I(N__29221));
    InMux I__5158 (
            .O(N__29273),
            .I(N__29221));
    LocalMux I__5157 (
            .O(N__29268),
            .I(N__29214));
    LocalMux I__5156 (
            .O(N__29263),
            .I(N__29214));
    Span4Mux_h I__5155 (
            .O(N__29258),
            .I(N__29214));
    Span4Mux_h I__5154 (
            .O(N__29255),
            .I(N__29211));
    LocalMux I__5153 (
            .O(N__29246),
            .I(N__29208));
    LocalMux I__5152 (
            .O(N__29237),
            .I(N__29199));
    LocalMux I__5151 (
            .O(N__29230),
            .I(N__29199));
    LocalMux I__5150 (
            .O(N__29221),
            .I(N__29199));
    Span4Mux_v I__5149 (
            .O(N__29214),
            .I(N__29199));
    Span4Mux_v I__5148 (
            .O(N__29211),
            .I(N__29196));
    Span4Mux_v I__5147 (
            .O(N__29208),
            .I(N__29191));
    Span4Mux_v I__5146 (
            .O(N__29199),
            .I(N__29191));
    Span4Mux_v I__5145 (
            .O(N__29196),
            .I(N__29188));
    Odrv4 I__5144 (
            .O(N__29191),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__5143 (
            .O(N__29188),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    InMux I__5142 (
            .O(N__29183),
            .I(N__29180));
    LocalMux I__5141 (
            .O(N__29180),
            .I(N__29177));
    Span4Mux_v I__5140 (
            .O(N__29177),
            .I(N__29174));
    Span4Mux_h I__5139 (
            .O(N__29174),
            .I(N__29171));
    Odrv4 I__5138 (
            .O(N__29171),
            .I(\phase_controller_inst1.stoper_hc.un6_running_1 ));
    CascadeMux I__5137 (
            .O(N__29168),
            .I(N__29164));
    InMux I__5136 (
            .O(N__29167),
            .I(N__29161));
    InMux I__5135 (
            .O(N__29164),
            .I(N__29157));
    LocalMux I__5134 (
            .O(N__29161),
            .I(N__29154));
    InMux I__5133 (
            .O(N__29160),
            .I(N__29151));
    LocalMux I__5132 (
            .O(N__29157),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__5131 (
            .O(N__29154),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__5130 (
            .O(N__29151),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    CascadeMux I__5129 (
            .O(N__29144),
            .I(N__29141));
    InMux I__5128 (
            .O(N__29141),
            .I(N__29138));
    LocalMux I__5127 (
            .O(N__29138),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__5126 (
            .O(N__29135),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__5125 (
            .O(N__29132),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__5124 (
            .O(N__29129),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__5123 (
            .O(N__29126),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__5122 (
            .O(N__29123),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__5121 (
            .O(N__29120),
            .I(bfn_12_14_0_));
    InMux I__5120 (
            .O(N__29117),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__5119 (
            .O(N__29114),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__5118 (
            .O(N__29111),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__5117 (
            .O(N__29108),
            .I(N__29105));
    LocalMux I__5116 (
            .O(N__29105),
            .I(N__29101));
    InMux I__5115 (
            .O(N__29104),
            .I(N__29098));
    Span4Mux_v I__5114 (
            .O(N__29101),
            .I(N__29092));
    LocalMux I__5113 (
            .O(N__29098),
            .I(N__29092));
    InMux I__5112 (
            .O(N__29097),
            .I(N__29089));
    Odrv4 I__5111 (
            .O(N__29092),
            .I(il_min_comp1_D2));
    LocalMux I__5110 (
            .O(N__29089),
            .I(il_min_comp1_D2));
    InMux I__5109 (
            .O(N__29084),
            .I(N__29080));
    InMux I__5108 (
            .O(N__29083),
            .I(N__29077));
    LocalMux I__5107 (
            .O(N__29080),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__5106 (
            .O(N__29077),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__5105 (
            .O(N__29072),
            .I(N__29068));
    InMux I__5104 (
            .O(N__29071),
            .I(N__29065));
    LocalMux I__5103 (
            .O(N__29068),
            .I(N__29059));
    LocalMux I__5102 (
            .O(N__29065),
            .I(N__29059));
    InMux I__5101 (
            .O(N__29064),
            .I(N__29056));
    Odrv4 I__5100 (
            .O(N__29059),
            .I(il_max_comp1_D2));
    LocalMux I__5099 (
            .O(N__29056),
            .I(il_max_comp1_D2));
    InMux I__5098 (
            .O(N__29051),
            .I(N__29045));
    InMux I__5097 (
            .O(N__29050),
            .I(N__29045));
    LocalMux I__5096 (
            .O(N__29045),
            .I(\phase_controller_inst1.N_56 ));
    CascadeMux I__5095 (
            .O(N__29042),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    CascadeMux I__5094 (
            .O(N__29039),
            .I(N__29036));
    InMux I__5093 (
            .O(N__29036),
            .I(N__29033));
    LocalMux I__5092 (
            .O(N__29033),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ));
    InMux I__5091 (
            .O(N__29030),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ));
    InMux I__5090 (
            .O(N__29027),
            .I(N__29024));
    LocalMux I__5089 (
            .O(N__29024),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNII3DZ0Z41 ));
    InMux I__5088 (
            .O(N__29021),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__5087 (
            .O(N__29018),
            .I(N__29015));
    LocalMux I__5086 (
            .O(N__29015),
            .I(N__29012));
    Span4Mux_v I__5085 (
            .O(N__29012),
            .I(N__29009));
    Odrv4 I__5084 (
            .O(N__29009),
            .I(il_max_comp1_D1));
    InMux I__5083 (
            .O(N__29006),
            .I(N__29003));
    LocalMux I__5082 (
            .O(N__29003),
            .I(N__29000));
    Odrv12 I__5081 (
            .O(N__29000),
            .I(il_min_comp2_D1));
    InMux I__5080 (
            .O(N__28997),
            .I(N__28994));
    LocalMux I__5079 (
            .O(N__28994),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    InMux I__5078 (
            .O(N__28991),
            .I(N__28988));
    LocalMux I__5077 (
            .O(N__28988),
            .I(\phase_controller_inst1.N_55 ));
    InMux I__5076 (
            .O(N__28985),
            .I(N__28978));
    InMux I__5075 (
            .O(N__28984),
            .I(N__28978));
    InMux I__5074 (
            .O(N__28983),
            .I(N__28975));
    LocalMux I__5073 (
            .O(N__28978),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__5072 (
            .O(N__28975),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    CascadeMux I__5071 (
            .O(N__28970),
            .I(N__28966));
    InMux I__5070 (
            .O(N__28969),
            .I(N__28959));
    InMux I__5069 (
            .O(N__28966),
            .I(N__28959));
    InMux I__5068 (
            .O(N__28965),
            .I(N__28956));
    InMux I__5067 (
            .O(N__28964),
            .I(N__28953));
    LocalMux I__5066 (
            .O(N__28959),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__5065 (
            .O(N__28956),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__5064 (
            .O(N__28953),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__5063 (
            .O(N__28946),
            .I(N__28943));
    LocalMux I__5062 (
            .O(N__28943),
            .I(N__28940));
    Span4Mux_h I__5061 (
            .O(N__28940),
            .I(N__28937));
    Odrv4 I__5060 (
            .O(N__28937),
            .I(\phase_controller_inst1.start_timer_tr_0_sqmuxa ));
    InMux I__5059 (
            .O(N__28934),
            .I(N__28931));
    LocalMux I__5058 (
            .O(N__28931),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5 ));
    InMux I__5057 (
            .O(N__28928),
            .I(N__28921));
    InMux I__5056 (
            .O(N__28927),
            .I(N__28921));
    InMux I__5055 (
            .O(N__28926),
            .I(N__28918));
    LocalMux I__5054 (
            .O(N__28921),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO ));
    LocalMux I__5053 (
            .O(N__28918),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO ));
    InMux I__5052 (
            .O(N__28913),
            .I(N__28909));
    InMux I__5051 (
            .O(N__28912),
            .I(N__28906));
    LocalMux I__5050 (
            .O(N__28909),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__5049 (
            .O(N__28906),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__5048 (
            .O(N__28901),
            .I(N__28898));
    InMux I__5047 (
            .O(N__28898),
            .I(N__28893));
    InMux I__5046 (
            .O(N__28897),
            .I(N__28890));
    InMux I__5045 (
            .O(N__28896),
            .I(N__28887));
    LocalMux I__5044 (
            .O(N__28893),
            .I(N__28884));
    LocalMux I__5043 (
            .O(N__28890),
            .I(N__28881));
    LocalMux I__5042 (
            .O(N__28887),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__5041 (
            .O(N__28884),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__5040 (
            .O(N__28881),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    CEMux I__5039 (
            .O(N__28874),
            .I(N__28863));
    CEMux I__5038 (
            .O(N__28873),
            .I(N__28859));
    CEMux I__5037 (
            .O(N__28872),
            .I(N__28856));
    CEMux I__5036 (
            .O(N__28871),
            .I(N__28853));
    InMux I__5035 (
            .O(N__28870),
            .I(N__28844));
    InMux I__5034 (
            .O(N__28869),
            .I(N__28844));
    InMux I__5033 (
            .O(N__28868),
            .I(N__28844));
    InMux I__5032 (
            .O(N__28867),
            .I(N__28844));
    InMux I__5031 (
            .O(N__28866),
            .I(N__28841));
    LocalMux I__5030 (
            .O(N__28863),
            .I(N__28838));
    CEMux I__5029 (
            .O(N__28862),
            .I(N__28835));
    LocalMux I__5028 (
            .O(N__28859),
            .I(N__28830));
    LocalMux I__5027 (
            .O(N__28856),
            .I(N__28830));
    LocalMux I__5026 (
            .O(N__28853),
            .I(N__28825));
    LocalMux I__5025 (
            .O(N__28844),
            .I(N__28808));
    LocalMux I__5024 (
            .O(N__28841),
            .I(N__28808));
    Sp12to4 I__5023 (
            .O(N__28838),
            .I(N__28805));
    LocalMux I__5022 (
            .O(N__28835),
            .I(N__28802));
    Span4Mux_h I__5021 (
            .O(N__28830),
            .I(N__28799));
    InMux I__5020 (
            .O(N__28829),
            .I(N__28794));
    InMux I__5019 (
            .O(N__28828),
            .I(N__28794));
    Span4Mux_h I__5018 (
            .O(N__28825),
            .I(N__28791));
    InMux I__5017 (
            .O(N__28824),
            .I(N__28784));
    InMux I__5016 (
            .O(N__28823),
            .I(N__28784));
    InMux I__5015 (
            .O(N__28822),
            .I(N__28784));
    InMux I__5014 (
            .O(N__28821),
            .I(N__28781));
    InMux I__5013 (
            .O(N__28820),
            .I(N__28772));
    InMux I__5012 (
            .O(N__28819),
            .I(N__28772));
    InMux I__5011 (
            .O(N__28818),
            .I(N__28772));
    InMux I__5010 (
            .O(N__28817),
            .I(N__28772));
    InMux I__5009 (
            .O(N__28816),
            .I(N__28763));
    InMux I__5008 (
            .O(N__28815),
            .I(N__28763));
    InMux I__5007 (
            .O(N__28814),
            .I(N__28763));
    InMux I__5006 (
            .O(N__28813),
            .I(N__28763));
    Span12Mux_s6_v I__5005 (
            .O(N__28808),
            .I(N__28758));
    Span12Mux_v I__5004 (
            .O(N__28805),
            .I(N__28758));
    Span4Mux_h I__5003 (
            .O(N__28802),
            .I(N__28753));
    Span4Mux_v I__5002 (
            .O(N__28799),
            .I(N__28753));
    LocalMux I__5001 (
            .O(N__28794),
            .I(N__28748));
    Span4Mux_v I__5000 (
            .O(N__28791),
            .I(N__28748));
    LocalMux I__4999 (
            .O(N__28784),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    LocalMux I__4998 (
            .O(N__28781),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    LocalMux I__4997 (
            .O(N__28772),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    LocalMux I__4996 (
            .O(N__28763),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv12 I__4995 (
            .O(N__28758),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__4994 (
            .O(N__28753),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__4993 (
            .O(N__28748),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    InMux I__4992 (
            .O(N__28733),
            .I(N__28729));
    InMux I__4991 (
            .O(N__28732),
            .I(N__28726));
    LocalMux I__4990 (
            .O(N__28729),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    LocalMux I__4989 (
            .O(N__28726),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    CascadeMux I__4988 (
            .O(N__28721),
            .I(N__28717));
    CascadeMux I__4987 (
            .O(N__28720),
            .I(N__28714));
    InMux I__4986 (
            .O(N__28717),
            .I(N__28708));
    InMux I__4985 (
            .O(N__28714),
            .I(N__28703));
    InMux I__4984 (
            .O(N__28713),
            .I(N__28703));
    InMux I__4983 (
            .O(N__28712),
            .I(N__28698));
    InMux I__4982 (
            .O(N__28711),
            .I(N__28698));
    LocalMux I__4981 (
            .O(N__28708),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    LocalMux I__4980 (
            .O(N__28703),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    LocalMux I__4979 (
            .O(N__28698),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    InMux I__4978 (
            .O(N__28691),
            .I(N__28686));
    InMux I__4977 (
            .O(N__28690),
            .I(N__28682));
    InMux I__4976 (
            .O(N__28689),
            .I(N__28679));
    LocalMux I__4975 (
            .O(N__28686),
            .I(N__28676));
    InMux I__4974 (
            .O(N__28685),
            .I(N__28673));
    LocalMux I__4973 (
            .O(N__28682),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__4972 (
            .O(N__28679),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__4971 (
            .O(N__28676),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__4970 (
            .O(N__28673),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    IoInMux I__4969 (
            .O(N__28664),
            .I(N__28661));
    LocalMux I__4968 (
            .O(N__28661),
            .I(N__28658));
    Span4Mux_s1_v I__4967 (
            .O(N__28658),
            .I(N__28655));
    Odrv4 I__4966 (
            .O(N__28655),
            .I(s4_phy_c));
    CascadeMux I__4965 (
            .O(N__28652),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_ ));
    InMux I__4964 (
            .O(N__28649),
            .I(N__28646));
    LocalMux I__4963 (
            .O(N__28646),
            .I(N__28640));
    InMux I__4962 (
            .O(N__28645),
            .I(N__28637));
    InMux I__4961 (
            .O(N__28644),
            .I(N__28634));
    InMux I__4960 (
            .O(N__28643),
            .I(N__28631));
    Span4Mux_h I__4959 (
            .O(N__28640),
            .I(N__28628));
    LocalMux I__4958 (
            .O(N__28637),
            .I(N__28623));
    LocalMux I__4957 (
            .O(N__28634),
            .I(N__28623));
    LocalMux I__4956 (
            .O(N__28631),
            .I(elapsed_time_ns_1_RNIQURR91_0_3));
    Odrv4 I__4955 (
            .O(N__28628),
            .I(elapsed_time_ns_1_RNIQURR91_0_3));
    Odrv4 I__4954 (
            .O(N__28623),
            .I(elapsed_time_ns_1_RNIQURR91_0_3));
    CascadeMux I__4953 (
            .O(N__28616),
            .I(elapsed_time_ns_1_RNIQURR91_0_3_cascade_));
    InMux I__4952 (
            .O(N__28613),
            .I(N__28610));
    LocalMux I__4951 (
            .O(N__28610),
            .I(N__28607));
    Odrv4 I__4950 (
            .O(N__28607),
            .I(\phase_controller_inst1.stoper_hc.N_283 ));
    InMux I__4949 (
            .O(N__28604),
            .I(N__28598));
    InMux I__4948 (
            .O(N__28603),
            .I(N__28598));
    LocalMux I__4947 (
            .O(N__28598),
            .I(N__28595));
    Span4Mux_v I__4946 (
            .O(N__28595),
            .I(N__28591));
    InMux I__4945 (
            .O(N__28594),
            .I(N__28588));
    Odrv4 I__4944 (
            .O(N__28591),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24 ));
    LocalMux I__4943 (
            .O(N__28588),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24 ));
    CascadeMux I__4942 (
            .O(N__28583),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_ ));
    InMux I__4941 (
            .O(N__28580),
            .I(N__28577));
    LocalMux I__4940 (
            .O(N__28577),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15 ));
    InMux I__4939 (
            .O(N__28574),
            .I(N__28571));
    LocalMux I__4938 (
            .O(N__28571),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10 ));
    CascadeMux I__4937 (
            .O(N__28568),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10_cascade_ ));
    CascadeMux I__4936 (
            .O(N__28565),
            .I(N__28561));
    CascadeMux I__4935 (
            .O(N__28564),
            .I(N__28558));
    InMux I__4934 (
            .O(N__28561),
            .I(N__28553));
    InMux I__4933 (
            .O(N__28558),
            .I(N__28553));
    LocalMux I__4932 (
            .O(N__28553),
            .I(N__28549));
    InMux I__4931 (
            .O(N__28552),
            .I(N__28546));
    Span4Mux_h I__4930 (
            .O(N__28549),
            .I(N__28543));
    LocalMux I__4929 (
            .O(N__28546),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2 ));
    Odrv4 I__4928 (
            .O(N__28543),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2 ));
    InMux I__4927 (
            .O(N__28538),
            .I(N__28535));
    LocalMux I__4926 (
            .O(N__28535),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4 ));
    CascadeMux I__4925 (
            .O(N__28532),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_ ));
    InMux I__4924 (
            .O(N__28529),
            .I(N__28526));
    LocalMux I__4923 (
            .O(N__28526),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31 ));
    CascadeMux I__4922 (
            .O(N__28523),
            .I(\delay_measurement_inst.delay_hc_timer.N_382_i_cascade_ ));
    InMux I__4921 (
            .O(N__28520),
            .I(N__28516));
    InMux I__4920 (
            .O(N__28519),
            .I(N__28513));
    LocalMux I__4919 (
            .O(N__28516),
            .I(elapsed_time_ns_1_RNIS5ND11_0_24));
    LocalMux I__4918 (
            .O(N__28513),
            .I(elapsed_time_ns_1_RNIS5ND11_0_24));
    InMux I__4917 (
            .O(N__28508),
            .I(N__28504));
    InMux I__4916 (
            .O(N__28507),
            .I(N__28501));
    LocalMux I__4915 (
            .O(N__28504),
            .I(elapsed_time_ns_1_RNIT6ND11_0_25));
    LocalMux I__4914 (
            .O(N__28501),
            .I(elapsed_time_ns_1_RNIT6ND11_0_25));
    CascadeMux I__4913 (
            .O(N__28496),
            .I(N__28491));
    CascadeMux I__4912 (
            .O(N__28495),
            .I(N__28486));
    CascadeMux I__4911 (
            .O(N__28494),
            .I(N__28482));
    InMux I__4910 (
            .O(N__28491),
            .I(N__28477));
    InMux I__4909 (
            .O(N__28490),
            .I(N__28474));
    InMux I__4908 (
            .O(N__28489),
            .I(N__28471));
    InMux I__4907 (
            .O(N__28486),
            .I(N__28468));
    InMux I__4906 (
            .O(N__28485),
            .I(N__28465));
    InMux I__4905 (
            .O(N__28482),
            .I(N__28462));
    InMux I__4904 (
            .O(N__28481),
            .I(N__28458));
    InMux I__4903 (
            .O(N__28480),
            .I(N__28455));
    LocalMux I__4902 (
            .O(N__28477),
            .I(N__28452));
    LocalMux I__4901 (
            .O(N__28474),
            .I(N__28447));
    LocalMux I__4900 (
            .O(N__28471),
            .I(N__28447));
    LocalMux I__4899 (
            .O(N__28468),
            .I(N__28444));
    LocalMux I__4898 (
            .O(N__28465),
            .I(N__28439));
    LocalMux I__4897 (
            .O(N__28462),
            .I(N__28439));
    InMux I__4896 (
            .O(N__28461),
            .I(N__28436));
    LocalMux I__4895 (
            .O(N__28458),
            .I(N__28433));
    LocalMux I__4894 (
            .O(N__28455),
            .I(N__28426));
    Span4Mux_h I__4893 (
            .O(N__28452),
            .I(N__28426));
    Span4Mux_h I__4892 (
            .O(N__28447),
            .I(N__28426));
    Span4Mux_v I__4891 (
            .O(N__28444),
            .I(N__28421));
    Span4Mux_h I__4890 (
            .O(N__28439),
            .I(N__28421));
    LocalMux I__4889 (
            .O(N__28436),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    Odrv12 I__4888 (
            .O(N__28433),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    Odrv4 I__4887 (
            .O(N__28426),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    Odrv4 I__4886 (
            .O(N__28421),
            .I(elapsed_time_ns_1_RNIS4MD11_0_15));
    CascadeMux I__4885 (
            .O(N__28412),
            .I(N__28408));
    CascadeMux I__4884 (
            .O(N__28411),
            .I(N__28405));
    InMux I__4883 (
            .O(N__28408),
            .I(N__28402));
    InMux I__4882 (
            .O(N__28405),
            .I(N__28399));
    LocalMux I__4881 (
            .O(N__28402),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16 ));
    LocalMux I__4880 (
            .O(N__28399),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16 ));
    InMux I__4879 (
            .O(N__28394),
            .I(N__28390));
    InMux I__4878 (
            .O(N__28393),
            .I(N__28387));
    LocalMux I__4877 (
            .O(N__28390),
            .I(elapsed_time_ns_1_RNIQ3ND11_0_22));
    LocalMux I__4876 (
            .O(N__28387),
            .I(elapsed_time_ns_1_RNIQ3ND11_0_22));
    CascadeMux I__4875 (
            .O(N__28382),
            .I(N__28379));
    InMux I__4874 (
            .O(N__28379),
            .I(N__28375));
    InMux I__4873 (
            .O(N__28378),
            .I(N__28372));
    LocalMux I__4872 (
            .O(N__28375),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31 ));
    LocalMux I__4871 (
            .O(N__28372),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31 ));
    CascadeMux I__4870 (
            .O(N__28367),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31_cascade_ ));
    CascadeMux I__4869 (
            .O(N__28364),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_));
    CascadeMux I__4868 (
            .O(N__28361),
            .I(N__28358));
    InMux I__4867 (
            .O(N__28358),
            .I(N__28355));
    LocalMux I__4866 (
            .O(N__28355),
            .I(N__28351));
    InMux I__4865 (
            .O(N__28354),
            .I(N__28348));
    Odrv4 I__4864 (
            .O(N__28351),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ));
    LocalMux I__4863 (
            .O(N__28348),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ));
    CascadeMux I__4862 (
            .O(N__28343),
            .I(N__28340));
    InMux I__4861 (
            .O(N__28340),
            .I(N__28334));
    InMux I__4860 (
            .O(N__28339),
            .I(N__28331));
    InMux I__4859 (
            .O(N__28338),
            .I(N__28328));
    InMux I__4858 (
            .O(N__28337),
            .I(N__28325));
    LocalMux I__4857 (
            .O(N__28334),
            .I(N__28320));
    LocalMux I__4856 (
            .O(N__28331),
            .I(N__28320));
    LocalMux I__4855 (
            .O(N__28328),
            .I(elapsed_time_ns_1_RNIA3DJ11_0_4));
    LocalMux I__4854 (
            .O(N__28325),
            .I(elapsed_time_ns_1_RNIA3DJ11_0_4));
    Odrv4 I__4853 (
            .O(N__28320),
            .I(elapsed_time_ns_1_RNIA3DJ11_0_4));
    InMux I__4852 (
            .O(N__28313),
            .I(N__28299));
    InMux I__4851 (
            .O(N__28312),
            .I(N__28299));
    InMux I__4850 (
            .O(N__28311),
            .I(N__28299));
    CascadeMux I__4849 (
            .O(N__28310),
            .I(N__28295));
    InMux I__4848 (
            .O(N__28309),
            .I(N__28281));
    InMux I__4847 (
            .O(N__28308),
            .I(N__28281));
    InMux I__4846 (
            .O(N__28307),
            .I(N__28281));
    InMux I__4845 (
            .O(N__28306),
            .I(N__28281));
    LocalMux I__4844 (
            .O(N__28299),
            .I(N__28278));
    InMux I__4843 (
            .O(N__28298),
            .I(N__28273));
    InMux I__4842 (
            .O(N__28295),
            .I(N__28273));
    InMux I__4841 (
            .O(N__28294),
            .I(N__28262));
    InMux I__4840 (
            .O(N__28293),
            .I(N__28262));
    InMux I__4839 (
            .O(N__28292),
            .I(N__28262));
    InMux I__4838 (
            .O(N__28291),
            .I(N__28262));
    InMux I__4837 (
            .O(N__28290),
            .I(N__28262));
    LocalMux I__4836 (
            .O(N__28281),
            .I(N__28259));
    Span4Mux_h I__4835 (
            .O(N__28278),
            .I(N__28256));
    LocalMux I__4834 (
            .O(N__28273),
            .I(\phase_controller_inst1.stoper_hc.N_325 ));
    LocalMux I__4833 (
            .O(N__28262),
            .I(\phase_controller_inst1.stoper_hc.N_325 ));
    Odrv4 I__4832 (
            .O(N__28259),
            .I(\phase_controller_inst1.stoper_hc.N_325 ));
    Odrv4 I__4831 (
            .O(N__28256),
            .I(\phase_controller_inst1.stoper_hc.N_325 ));
    InMux I__4830 (
            .O(N__28247),
            .I(N__28215));
    InMux I__4829 (
            .O(N__28246),
            .I(N__28215));
    InMux I__4828 (
            .O(N__28245),
            .I(N__28215));
    InMux I__4827 (
            .O(N__28244),
            .I(N__28215));
    InMux I__4826 (
            .O(N__28243),
            .I(N__28215));
    InMux I__4825 (
            .O(N__28242),
            .I(N__28212));
    InMux I__4824 (
            .O(N__28241),
            .I(N__28201));
    InMux I__4823 (
            .O(N__28240),
            .I(N__28201));
    InMux I__4822 (
            .O(N__28239),
            .I(N__28201));
    InMux I__4821 (
            .O(N__28238),
            .I(N__28201));
    InMux I__4820 (
            .O(N__28237),
            .I(N__28201));
    InMux I__4819 (
            .O(N__28236),
            .I(N__28186));
    InMux I__4818 (
            .O(N__28235),
            .I(N__28186));
    InMux I__4817 (
            .O(N__28234),
            .I(N__28186));
    InMux I__4816 (
            .O(N__28233),
            .I(N__28186));
    InMux I__4815 (
            .O(N__28232),
            .I(N__28186));
    InMux I__4814 (
            .O(N__28231),
            .I(N__28186));
    InMux I__4813 (
            .O(N__28230),
            .I(N__28186));
    InMux I__4812 (
            .O(N__28229),
            .I(N__28177));
    InMux I__4811 (
            .O(N__28228),
            .I(N__28177));
    InMux I__4810 (
            .O(N__28227),
            .I(N__28177));
    InMux I__4809 (
            .O(N__28226),
            .I(N__28177));
    LocalMux I__4808 (
            .O(N__28215),
            .I(N__28160));
    LocalMux I__4807 (
            .O(N__28212),
            .I(N__28157));
    LocalMux I__4806 (
            .O(N__28201),
            .I(N__28150));
    LocalMux I__4805 (
            .O(N__28186),
            .I(N__28150));
    LocalMux I__4804 (
            .O(N__28177),
            .I(N__28150));
    InMux I__4803 (
            .O(N__28176),
            .I(N__28147));
    InMux I__4802 (
            .O(N__28175),
            .I(N__28140));
    InMux I__4801 (
            .O(N__28174),
            .I(N__28140));
    InMux I__4800 (
            .O(N__28173),
            .I(N__28140));
    InMux I__4799 (
            .O(N__28172),
            .I(N__28127));
    InMux I__4798 (
            .O(N__28171),
            .I(N__28127));
    InMux I__4797 (
            .O(N__28170),
            .I(N__28127));
    InMux I__4796 (
            .O(N__28169),
            .I(N__28127));
    InMux I__4795 (
            .O(N__28168),
            .I(N__28127));
    InMux I__4794 (
            .O(N__28167),
            .I(N__28127));
    InMux I__4793 (
            .O(N__28166),
            .I(N__28118));
    InMux I__4792 (
            .O(N__28165),
            .I(N__28118));
    InMux I__4791 (
            .O(N__28164),
            .I(N__28118));
    InMux I__4790 (
            .O(N__28163),
            .I(N__28118));
    Span4Mux_h I__4789 (
            .O(N__28160),
            .I(N__28115));
    Span4Mux_h I__4788 (
            .O(N__28157),
            .I(N__28106));
    Span4Mux_v I__4787 (
            .O(N__28150),
            .I(N__28106));
    LocalMux I__4786 (
            .O(N__28147),
            .I(N__28106));
    LocalMux I__4785 (
            .O(N__28140),
            .I(N__28106));
    LocalMux I__4784 (
            .O(N__28127),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    LocalMux I__4783 (
            .O(N__28118),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    Odrv4 I__4782 (
            .O(N__28115),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    Odrv4 I__4781 (
            .O(N__28106),
            .I(elapsed_time_ns_1_RNIQ4OD11_0_31));
    CascadeMux I__4780 (
            .O(N__28097),
            .I(N__28094));
    InMux I__4779 (
            .O(N__28094),
            .I(N__28091));
    LocalMux I__4778 (
            .O(N__28091),
            .I(N__28087));
    InMux I__4777 (
            .O(N__28090),
            .I(N__28083));
    Span4Mux_v I__4776 (
            .O(N__28087),
            .I(N__28080));
    InMux I__4775 (
            .O(N__28086),
            .I(N__28077));
    LocalMux I__4774 (
            .O(N__28083),
            .I(elapsed_time_ns_1_RNIB4DJ11_0_5));
    Odrv4 I__4773 (
            .O(N__28080),
            .I(elapsed_time_ns_1_RNIB4DJ11_0_5));
    LocalMux I__4772 (
            .O(N__28077),
            .I(elapsed_time_ns_1_RNIB4DJ11_0_5));
    CascadeMux I__4771 (
            .O(N__28070),
            .I(N__28057));
    InMux I__4770 (
            .O(N__28069),
            .I(N__28049));
    InMux I__4769 (
            .O(N__28068),
            .I(N__28049));
    InMux I__4768 (
            .O(N__28067),
            .I(N__28049));
    InMux I__4767 (
            .O(N__28066),
            .I(N__28046));
    InMux I__4766 (
            .O(N__28065),
            .I(N__28039));
    InMux I__4765 (
            .O(N__28064),
            .I(N__28039));
    InMux I__4764 (
            .O(N__28063),
            .I(N__28039));
    InMux I__4763 (
            .O(N__28062),
            .I(N__28028));
    InMux I__4762 (
            .O(N__28061),
            .I(N__28028));
    InMux I__4761 (
            .O(N__28060),
            .I(N__28028));
    InMux I__4760 (
            .O(N__28057),
            .I(N__28028));
    InMux I__4759 (
            .O(N__28056),
            .I(N__28028));
    LocalMux I__4758 (
            .O(N__28049),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    LocalMux I__4757 (
            .O(N__28046),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    LocalMux I__4756 (
            .O(N__28039),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    LocalMux I__4755 (
            .O(N__28028),
            .I(\phase_controller_inst1.stoper_hc.N_327 ));
    InMux I__4754 (
            .O(N__28019),
            .I(N__28015));
    InMux I__4753 (
            .O(N__28018),
            .I(N__28012));
    LocalMux I__4752 (
            .O(N__28015),
            .I(elapsed_time_ns_1_RNIP3OD11_0_30));
    LocalMux I__4751 (
            .O(N__28012),
            .I(elapsed_time_ns_1_RNIP3OD11_0_30));
    InMux I__4750 (
            .O(N__28007),
            .I(N__28003));
    InMux I__4749 (
            .O(N__28006),
            .I(N__28000));
    LocalMux I__4748 (
            .O(N__28003),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15 ));
    LocalMux I__4747 (
            .O(N__28000),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15 ));
    CascadeMux I__4746 (
            .O(N__27995),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31_cascade_ ));
    InMux I__4745 (
            .O(N__27992),
            .I(N__27988));
    CascadeMux I__4744 (
            .O(N__27991),
            .I(N__27985));
    LocalMux I__4743 (
            .O(N__27988),
            .I(N__27981));
    InMux I__4742 (
            .O(N__27985),
            .I(N__27978));
    InMux I__4741 (
            .O(N__27984),
            .I(N__27975));
    Span4Mux_h I__4740 (
            .O(N__27981),
            .I(N__27972));
    LocalMux I__4739 (
            .O(N__27978),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ));
    LocalMux I__4738 (
            .O(N__27975),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ));
    Odrv4 I__4737 (
            .O(N__27972),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ));
    CascadeMux I__4736 (
            .O(N__27965),
            .I(N__27961));
    CascadeMux I__4735 (
            .O(N__27964),
            .I(N__27954));
    InMux I__4734 (
            .O(N__27961),
            .I(N__27947));
    InMux I__4733 (
            .O(N__27960),
            .I(N__27947));
    InMux I__4732 (
            .O(N__27959),
            .I(N__27947));
    CascadeMux I__4731 (
            .O(N__27958),
            .I(N__27943));
    CascadeMux I__4730 (
            .O(N__27957),
            .I(N__27940));
    InMux I__4729 (
            .O(N__27954),
            .I(N__27936));
    LocalMux I__4728 (
            .O(N__27947),
            .I(N__27933));
    InMux I__4727 (
            .O(N__27946),
            .I(N__27928));
    InMux I__4726 (
            .O(N__27943),
            .I(N__27928));
    InMux I__4725 (
            .O(N__27940),
            .I(N__27925));
    InMux I__4724 (
            .O(N__27939),
            .I(N__27922));
    LocalMux I__4723 (
            .O(N__27936),
            .I(N__27917));
    Span4Mux_h I__4722 (
            .O(N__27933),
            .I(N__27917));
    LocalMux I__4721 (
            .O(N__27928),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2Z0Z_10 ));
    LocalMux I__4720 (
            .O(N__27925),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2Z0Z_10 ));
    LocalMux I__4719 (
            .O(N__27922),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2Z0Z_10 ));
    Odrv4 I__4718 (
            .O(N__27917),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2Z0Z_10 ));
    InMux I__4717 (
            .O(N__27908),
            .I(N__27904));
    CascadeMux I__4716 (
            .O(N__27907),
            .I(N__27901));
    LocalMux I__4715 (
            .O(N__27904),
            .I(N__27898));
    InMux I__4714 (
            .O(N__27901),
            .I(N__27893));
    Span4Mux_v I__4713 (
            .O(N__27898),
            .I(N__27890));
    InMux I__4712 (
            .O(N__27897),
            .I(N__27885));
    InMux I__4711 (
            .O(N__27896),
            .I(N__27885));
    LocalMux I__4710 (
            .O(N__27893),
            .I(elapsed_time_ns_1_RNIQ2MD11_0_13));
    Odrv4 I__4709 (
            .O(N__27890),
            .I(elapsed_time_ns_1_RNIQ2MD11_0_13));
    LocalMux I__4708 (
            .O(N__27885),
            .I(elapsed_time_ns_1_RNIQ2MD11_0_13));
    CascadeMux I__4707 (
            .O(N__27878),
            .I(N__27875));
    InMux I__4706 (
            .O(N__27875),
            .I(N__27858));
    InMux I__4705 (
            .O(N__27874),
            .I(N__27841));
    InMux I__4704 (
            .O(N__27873),
            .I(N__27841));
    InMux I__4703 (
            .O(N__27872),
            .I(N__27841));
    InMux I__4702 (
            .O(N__27871),
            .I(N__27841));
    InMux I__4701 (
            .O(N__27870),
            .I(N__27830));
    InMux I__4700 (
            .O(N__27869),
            .I(N__27830));
    InMux I__4699 (
            .O(N__27868),
            .I(N__27830));
    InMux I__4698 (
            .O(N__27867),
            .I(N__27830));
    InMux I__4697 (
            .O(N__27866),
            .I(N__27830));
    InMux I__4696 (
            .O(N__27865),
            .I(N__27819));
    InMux I__4695 (
            .O(N__27864),
            .I(N__27819));
    InMux I__4694 (
            .O(N__27863),
            .I(N__27819));
    InMux I__4693 (
            .O(N__27862),
            .I(N__27819));
    InMux I__4692 (
            .O(N__27861),
            .I(N__27819));
    LocalMux I__4691 (
            .O(N__27858),
            .I(N__27816));
    CascadeMux I__4690 (
            .O(N__27857),
            .I(N__27812));
    InMux I__4689 (
            .O(N__27856),
            .I(N__27807));
    InMux I__4688 (
            .O(N__27855),
            .I(N__27794));
    InMux I__4687 (
            .O(N__27854),
            .I(N__27794));
    InMux I__4686 (
            .O(N__27853),
            .I(N__27794));
    InMux I__4685 (
            .O(N__27852),
            .I(N__27794));
    InMux I__4684 (
            .O(N__27851),
            .I(N__27794));
    InMux I__4683 (
            .O(N__27850),
            .I(N__27794));
    LocalMux I__4682 (
            .O(N__27841),
            .I(N__27791));
    LocalMux I__4681 (
            .O(N__27830),
            .I(N__27784));
    LocalMux I__4680 (
            .O(N__27819),
            .I(N__27784));
    Span4Mux_h I__4679 (
            .O(N__27816),
            .I(N__27784));
    InMux I__4678 (
            .O(N__27815),
            .I(N__27777));
    InMux I__4677 (
            .O(N__27812),
            .I(N__27777));
    InMux I__4676 (
            .O(N__27811),
            .I(N__27777));
    InMux I__4675 (
            .O(N__27810),
            .I(N__27774));
    LocalMux I__4674 (
            .O(N__27807),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    LocalMux I__4673 (
            .O(N__27794),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    Odrv4 I__4672 (
            .O(N__27791),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    Odrv4 I__4671 (
            .O(N__27784),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    LocalMux I__4670 (
            .O(N__27777),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    LocalMux I__4669 (
            .O(N__27774),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    CascadeMux I__4668 (
            .O(N__27761),
            .I(N__27757));
    InMux I__4667 (
            .O(N__27760),
            .I(N__27754));
    InMux I__4666 (
            .O(N__27757),
            .I(N__27748));
    LocalMux I__4665 (
            .O(N__27754),
            .I(N__27745));
    InMux I__4664 (
            .O(N__27753),
            .I(N__27741));
    InMux I__4663 (
            .O(N__27752),
            .I(N__27738));
    InMux I__4662 (
            .O(N__27751),
            .I(N__27735));
    LocalMux I__4661 (
            .O(N__27748),
            .I(N__27732));
    Span4Mux_h I__4660 (
            .O(N__27745),
            .I(N__27729));
    InMux I__4659 (
            .O(N__27744),
            .I(N__27726));
    LocalMux I__4658 (
            .O(N__27741),
            .I(N__27723));
    LocalMux I__4657 (
            .O(N__27738),
            .I(N__27718));
    LocalMux I__4656 (
            .O(N__27735),
            .I(N__27718));
    Odrv4 I__4655 (
            .O(N__27732),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ));
    Odrv4 I__4654 (
            .O(N__27729),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ));
    LocalMux I__4653 (
            .O(N__27726),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ));
    Odrv4 I__4652 (
            .O(N__27723),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ));
    Odrv4 I__4651 (
            .O(N__27718),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ));
    InMux I__4650 (
            .O(N__27707),
            .I(N__27703));
    InMux I__4649 (
            .O(N__27706),
            .I(N__27698));
    LocalMux I__4648 (
            .O(N__27703),
            .I(N__27695));
    InMux I__4647 (
            .O(N__27702),
            .I(N__27692));
    InMux I__4646 (
            .O(N__27701),
            .I(N__27689));
    LocalMux I__4645 (
            .O(N__27698),
            .I(elapsed_time_ns_1_RNID6DJ11_0_7));
    Odrv4 I__4644 (
            .O(N__27695),
            .I(elapsed_time_ns_1_RNID6DJ11_0_7));
    LocalMux I__4643 (
            .O(N__27692),
            .I(elapsed_time_ns_1_RNID6DJ11_0_7));
    LocalMux I__4642 (
            .O(N__27689),
            .I(elapsed_time_ns_1_RNID6DJ11_0_7));
    InMux I__4641 (
            .O(N__27680),
            .I(N__27674));
    CascadeMux I__4640 (
            .O(N__27679),
            .I(N__27671));
    InMux I__4639 (
            .O(N__27678),
            .I(N__27668));
    InMux I__4638 (
            .O(N__27677),
            .I(N__27665));
    LocalMux I__4637 (
            .O(N__27674),
            .I(N__27662));
    InMux I__4636 (
            .O(N__27671),
            .I(N__27659));
    LocalMux I__4635 (
            .O(N__27668),
            .I(elapsed_time_ns_1_RNIE7DJ11_0_8));
    LocalMux I__4634 (
            .O(N__27665),
            .I(elapsed_time_ns_1_RNIE7DJ11_0_8));
    Odrv4 I__4633 (
            .O(N__27662),
            .I(elapsed_time_ns_1_RNIE7DJ11_0_8));
    LocalMux I__4632 (
            .O(N__27659),
            .I(elapsed_time_ns_1_RNIE7DJ11_0_8));
    CascadeMux I__4631 (
            .O(N__27650),
            .I(N__27646));
    CascadeMux I__4630 (
            .O(N__27649),
            .I(N__27643));
    InMux I__4629 (
            .O(N__27646),
            .I(N__27640));
    InMux I__4628 (
            .O(N__27643),
            .I(N__27637));
    LocalMux I__4627 (
            .O(N__27640),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ));
    LocalMux I__4626 (
            .O(N__27637),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ));
    CascadeMux I__4625 (
            .O(N__27632),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ));
    InMux I__4624 (
            .O(N__27629),
            .I(N__27623));
    InMux I__4623 (
            .O(N__27628),
            .I(N__27623));
    LocalMux I__4622 (
            .O(N__27623),
            .I(N__27619));
    InMux I__4621 (
            .O(N__27622),
            .I(N__27616));
    Odrv12 I__4620 (
            .O(N__27619),
            .I(elapsed_time_ns_1_RNIDP2KD1_0_1));
    LocalMux I__4619 (
            .O(N__27616),
            .I(elapsed_time_ns_1_RNIDP2KD1_0_1));
    InMux I__4618 (
            .O(N__27611),
            .I(N__27608));
    LocalMux I__4617 (
            .O(N__27608),
            .I(N__27605));
    Odrv4 I__4616 (
            .O(N__27605),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ));
    CascadeMux I__4615 (
            .O(N__27602),
            .I(elapsed_time_ns_1_RNIDP2KD1_0_1_cascade_));
    InMux I__4614 (
            .O(N__27599),
            .I(N__27595));
    InMux I__4613 (
            .O(N__27598),
            .I(N__27592));
    LocalMux I__4612 (
            .O(N__27595),
            .I(\phase_controller_inst1.stoper_hc.N_307 ));
    LocalMux I__4611 (
            .O(N__27592),
            .I(\phase_controller_inst1.stoper_hc.N_307 ));
    InMux I__4610 (
            .O(N__27587),
            .I(N__27583));
    InMux I__4609 (
            .O(N__27586),
            .I(N__27580));
    LocalMux I__4608 (
            .O(N__27583),
            .I(N__27576));
    LocalMux I__4607 (
            .O(N__27580),
            .I(N__27573));
    InMux I__4606 (
            .O(N__27579),
            .I(N__27570));
    Odrv12 I__4605 (
            .O(N__27576),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv12 I__4604 (
            .O(N__27573),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    LocalMux I__4603 (
            .O(N__27570),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__4602 (
            .O(N__27563),
            .I(N__27560));
    LocalMux I__4601 (
            .O(N__27560),
            .I(N__27557));
    Odrv4 I__4600 (
            .O(N__27557),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_10 ));
    CascadeMux I__4599 (
            .O(N__27554),
            .I(N__27551));
    InMux I__4598 (
            .O(N__27551),
            .I(N__27548));
    LocalMux I__4597 (
            .O(N__27548),
            .I(N__27545));
    Span4Mux_h I__4596 (
            .O(N__27545),
            .I(N__27542));
    Odrv4 I__4595 (
            .O(N__27542),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10 ));
    InMux I__4594 (
            .O(N__27539),
            .I(N__27536));
    LocalMux I__4593 (
            .O(N__27536),
            .I(N__27533));
    Odrv4 I__4592 (
            .O(N__27533),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    CascadeMux I__4591 (
            .O(N__27530),
            .I(N__27525));
    CascadeMux I__4590 (
            .O(N__27529),
            .I(N__27522));
    CascadeMux I__4589 (
            .O(N__27528),
            .I(N__27519));
    InMux I__4588 (
            .O(N__27525),
            .I(N__27516));
    InMux I__4587 (
            .O(N__27522),
            .I(N__27511));
    InMux I__4586 (
            .O(N__27519),
            .I(N__27511));
    LocalMux I__4585 (
            .O(N__27516),
            .I(N__27506));
    LocalMux I__4584 (
            .O(N__27511),
            .I(N__27503));
    InMux I__4583 (
            .O(N__27510),
            .I(N__27500));
    InMux I__4582 (
            .O(N__27509),
            .I(N__27497));
    Span12Mux_v I__4581 (
            .O(N__27506),
            .I(N__27494));
    Span4Mux_h I__4580 (
            .O(N__27503),
            .I(N__27491));
    LocalMux I__4579 (
            .O(N__27500),
            .I(N__27488));
    LocalMux I__4578 (
            .O(N__27497),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv12 I__4577 (
            .O(N__27494),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__4576 (
            .O(N__27491),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv12 I__4575 (
            .O(N__27488),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    CascadeMux I__4574 (
            .O(N__27479),
            .I(N__27476));
    InMux I__4573 (
            .O(N__27476),
            .I(N__27473));
    LocalMux I__4572 (
            .O(N__27473),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__4571 (
            .O(N__27470),
            .I(N__27467));
    LocalMux I__4570 (
            .O(N__27467),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__4569 (
            .O(N__27464),
            .I(N__27461));
    LocalMux I__4568 (
            .O(N__27461),
            .I(N__27455));
    InMux I__4567 (
            .O(N__27460),
            .I(N__27452));
    InMux I__4566 (
            .O(N__27459),
            .I(N__27449));
    InMux I__4565 (
            .O(N__27458),
            .I(N__27446));
    Span4Mux_v I__4564 (
            .O(N__27455),
            .I(N__27443));
    LocalMux I__4563 (
            .O(N__27452),
            .I(N__27440));
    LocalMux I__4562 (
            .O(N__27449),
            .I(N__27435));
    LocalMux I__4561 (
            .O(N__27446),
            .I(N__27435));
    Span4Mux_h I__4560 (
            .O(N__27443),
            .I(N__27432));
    Span4Mux_h I__4559 (
            .O(N__27440),
            .I(N__27429));
    Span4Mux_h I__4558 (
            .O(N__27435),
            .I(N__27426));
    Odrv4 I__4557 (
            .O(N__27432),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__4556 (
            .O(N__27429),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__4555 (
            .O(N__27426),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    CascadeMux I__4554 (
            .O(N__27419),
            .I(N__27416));
    InMux I__4553 (
            .O(N__27416),
            .I(N__27413));
    LocalMux I__4552 (
            .O(N__27413),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__4551 (
            .O(N__27410),
            .I(N__27407));
    LocalMux I__4550 (
            .O(N__27407),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    InMux I__4549 (
            .O(N__27404),
            .I(N__27392));
    InMux I__4548 (
            .O(N__27403),
            .I(N__27380));
    InMux I__4547 (
            .O(N__27402),
            .I(N__27380));
    InMux I__4546 (
            .O(N__27401),
            .I(N__27380));
    InMux I__4545 (
            .O(N__27400),
            .I(N__27359));
    InMux I__4544 (
            .O(N__27399),
            .I(N__27359));
    InMux I__4543 (
            .O(N__27398),
            .I(N__27359));
    InMux I__4542 (
            .O(N__27397),
            .I(N__27359));
    InMux I__4541 (
            .O(N__27396),
            .I(N__27359));
    InMux I__4540 (
            .O(N__27395),
            .I(N__27356));
    LocalMux I__4539 (
            .O(N__27392),
            .I(N__27353));
    InMux I__4538 (
            .O(N__27391),
            .I(N__27342));
    InMux I__4537 (
            .O(N__27390),
            .I(N__27342));
    InMux I__4536 (
            .O(N__27389),
            .I(N__27342));
    InMux I__4535 (
            .O(N__27388),
            .I(N__27342));
    InMux I__4534 (
            .O(N__27387),
            .I(N__27342));
    LocalMux I__4533 (
            .O(N__27380),
            .I(N__27339));
    InMux I__4532 (
            .O(N__27379),
            .I(N__27328));
    InMux I__4531 (
            .O(N__27378),
            .I(N__27328));
    InMux I__4530 (
            .O(N__27377),
            .I(N__27328));
    InMux I__4529 (
            .O(N__27376),
            .I(N__27328));
    InMux I__4528 (
            .O(N__27375),
            .I(N__27328));
    InMux I__4527 (
            .O(N__27374),
            .I(N__27311));
    InMux I__4526 (
            .O(N__27373),
            .I(N__27311));
    InMux I__4525 (
            .O(N__27372),
            .I(N__27311));
    InMux I__4524 (
            .O(N__27371),
            .I(N__27311));
    InMux I__4523 (
            .O(N__27370),
            .I(N__27311));
    LocalMux I__4522 (
            .O(N__27359),
            .I(N__27305));
    LocalMux I__4521 (
            .O(N__27356),
            .I(N__27305));
    Span4Mux_v I__4520 (
            .O(N__27353),
            .I(N__27302));
    LocalMux I__4519 (
            .O(N__27342),
            .I(N__27295));
    Span4Mux_h I__4518 (
            .O(N__27339),
            .I(N__27295));
    LocalMux I__4517 (
            .O(N__27328),
            .I(N__27295));
    InMux I__4516 (
            .O(N__27327),
            .I(N__27282));
    InMux I__4515 (
            .O(N__27326),
            .I(N__27282));
    InMux I__4514 (
            .O(N__27325),
            .I(N__27282));
    InMux I__4513 (
            .O(N__27324),
            .I(N__27282));
    InMux I__4512 (
            .O(N__27323),
            .I(N__27282));
    InMux I__4511 (
            .O(N__27322),
            .I(N__27282));
    LocalMux I__4510 (
            .O(N__27311),
            .I(N__27279));
    InMux I__4509 (
            .O(N__27310),
            .I(N__27276));
    Span4Mux_v I__4508 (
            .O(N__27305),
            .I(N__27273));
    Span4Mux_h I__4507 (
            .O(N__27302),
            .I(N__27268));
    Span4Mux_v I__4506 (
            .O(N__27295),
            .I(N__27268));
    LocalMux I__4505 (
            .O(N__27282),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__4504 (
            .O(N__27279),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__4503 (
            .O(N__27276),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__4502 (
            .O(N__27273),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__4501 (
            .O(N__27268),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    CascadeMux I__4500 (
            .O(N__27257),
            .I(N__27244));
    CascadeMux I__4499 (
            .O(N__27256),
            .I(N__27241));
    InMux I__4498 (
            .O(N__27255),
            .I(N__27225));
    InMux I__4497 (
            .O(N__27254),
            .I(N__27225));
    InMux I__4496 (
            .O(N__27253),
            .I(N__27225));
    InMux I__4495 (
            .O(N__27252),
            .I(N__27225));
    InMux I__4494 (
            .O(N__27251),
            .I(N__27225));
    InMux I__4493 (
            .O(N__27250),
            .I(N__27225));
    InMux I__4492 (
            .O(N__27249),
            .I(N__27210));
    InMux I__4491 (
            .O(N__27248),
            .I(N__27210));
    InMux I__4490 (
            .O(N__27247),
            .I(N__27210));
    InMux I__4489 (
            .O(N__27244),
            .I(N__27210));
    InMux I__4488 (
            .O(N__27241),
            .I(N__27210));
    InMux I__4487 (
            .O(N__27240),
            .I(N__27203));
    InMux I__4486 (
            .O(N__27239),
            .I(N__27203));
    InMux I__4485 (
            .O(N__27238),
            .I(N__27203));
    LocalMux I__4484 (
            .O(N__27225),
            .I(N__27190));
    InMux I__4483 (
            .O(N__27224),
            .I(N__27181));
    InMux I__4482 (
            .O(N__27223),
            .I(N__27181));
    InMux I__4481 (
            .O(N__27222),
            .I(N__27181));
    InMux I__4480 (
            .O(N__27221),
            .I(N__27181));
    LocalMux I__4479 (
            .O(N__27210),
            .I(N__27178));
    LocalMux I__4478 (
            .O(N__27203),
            .I(N__27175));
    InMux I__4477 (
            .O(N__27202),
            .I(N__27164));
    InMux I__4476 (
            .O(N__27201),
            .I(N__27164));
    InMux I__4475 (
            .O(N__27200),
            .I(N__27164));
    InMux I__4474 (
            .O(N__27199),
            .I(N__27164));
    InMux I__4473 (
            .O(N__27198),
            .I(N__27164));
    InMux I__4472 (
            .O(N__27197),
            .I(N__27153));
    InMux I__4471 (
            .O(N__27196),
            .I(N__27153));
    InMux I__4470 (
            .O(N__27195),
            .I(N__27153));
    InMux I__4469 (
            .O(N__27194),
            .I(N__27153));
    InMux I__4468 (
            .O(N__27193),
            .I(N__27153));
    Span4Mux_v I__4467 (
            .O(N__27190),
            .I(N__27150));
    LocalMux I__4466 (
            .O(N__27181),
            .I(N__27143));
    Span4Mux_h I__4465 (
            .O(N__27178),
            .I(N__27143));
    Span4Mux_v I__4464 (
            .O(N__27175),
            .I(N__27143));
    LocalMux I__4463 (
            .O(N__27164),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    LocalMux I__4462 (
            .O(N__27153),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    Odrv4 I__4461 (
            .O(N__27150),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    Odrv4 I__4460 (
            .O(N__27143),
            .I(\current_shift_inst.PI_CTRL.N_103 ));
    CascadeMux I__4459 (
            .O(N__27134),
            .I(N__27131));
    InMux I__4458 (
            .O(N__27131),
            .I(N__27128));
    LocalMux I__4457 (
            .O(N__27128),
            .I(N__27125));
    Span4Mux_v I__4456 (
            .O(N__27125),
            .I(N__27122));
    Odrv4 I__4455 (
            .O(N__27122),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    CascadeMux I__4454 (
            .O(N__27119),
            .I(N__27106));
    CascadeMux I__4453 (
            .O(N__27118),
            .I(N__27103));
    CascadeMux I__4452 (
            .O(N__27117),
            .I(N__27100));
    CascadeMux I__4451 (
            .O(N__27116),
            .I(N__27095));
    CascadeMux I__4450 (
            .O(N__27115),
            .I(N__27085));
    CascadeMux I__4449 (
            .O(N__27114),
            .I(N__27077));
    CascadeMux I__4448 (
            .O(N__27113),
            .I(N__27074));
    CascadeMux I__4447 (
            .O(N__27112),
            .I(N__27071));
    InMux I__4446 (
            .O(N__27111),
            .I(N__27056));
    InMux I__4445 (
            .O(N__27110),
            .I(N__27056));
    InMux I__4444 (
            .O(N__27109),
            .I(N__27056));
    InMux I__4443 (
            .O(N__27106),
            .I(N__27056));
    InMux I__4442 (
            .O(N__27103),
            .I(N__27056));
    InMux I__4441 (
            .O(N__27100),
            .I(N__27056));
    InMux I__4440 (
            .O(N__27099),
            .I(N__27049));
    InMux I__4439 (
            .O(N__27098),
            .I(N__27049));
    InMux I__4438 (
            .O(N__27095),
            .I(N__27049));
    CascadeMux I__4437 (
            .O(N__27094),
            .I(N__27044));
    CascadeMux I__4436 (
            .O(N__27093),
            .I(N__27041));
    CascadeMux I__4435 (
            .O(N__27092),
            .I(N__27038));
    CascadeMux I__4434 (
            .O(N__27091),
            .I(N__27032));
    CascadeMux I__4433 (
            .O(N__27090),
            .I(N__27029));
    InMux I__4432 (
            .O(N__27089),
            .I(N__27024));
    InMux I__4431 (
            .O(N__27088),
            .I(N__27024));
    InMux I__4430 (
            .O(N__27085),
            .I(N__27021));
    InMux I__4429 (
            .O(N__27084),
            .I(N__27010));
    InMux I__4428 (
            .O(N__27083),
            .I(N__27010));
    InMux I__4427 (
            .O(N__27082),
            .I(N__27010));
    InMux I__4426 (
            .O(N__27081),
            .I(N__27010));
    InMux I__4425 (
            .O(N__27080),
            .I(N__27010));
    InMux I__4424 (
            .O(N__27077),
            .I(N__27003));
    InMux I__4423 (
            .O(N__27074),
            .I(N__27003));
    InMux I__4422 (
            .O(N__27071),
            .I(N__27003));
    InMux I__4421 (
            .O(N__27070),
            .I(N__26998));
    InMux I__4420 (
            .O(N__27069),
            .I(N__26998));
    LocalMux I__4419 (
            .O(N__27056),
            .I(N__26995));
    LocalMux I__4418 (
            .O(N__27049),
            .I(N__26992));
    InMux I__4417 (
            .O(N__27048),
            .I(N__26981));
    InMux I__4416 (
            .O(N__27047),
            .I(N__26981));
    InMux I__4415 (
            .O(N__27044),
            .I(N__26981));
    InMux I__4414 (
            .O(N__27041),
            .I(N__26981));
    InMux I__4413 (
            .O(N__27038),
            .I(N__26981));
    InMux I__4412 (
            .O(N__27037),
            .I(N__26970));
    InMux I__4411 (
            .O(N__27036),
            .I(N__26970));
    InMux I__4410 (
            .O(N__27035),
            .I(N__26970));
    InMux I__4409 (
            .O(N__27032),
            .I(N__26970));
    InMux I__4408 (
            .O(N__27029),
            .I(N__26970));
    LocalMux I__4407 (
            .O(N__27024),
            .I(N__26959));
    LocalMux I__4406 (
            .O(N__27021),
            .I(N__26959));
    LocalMux I__4405 (
            .O(N__27010),
            .I(N__26959));
    LocalMux I__4404 (
            .O(N__27003),
            .I(N__26959));
    LocalMux I__4403 (
            .O(N__26998),
            .I(N__26959));
    Span4Mux_h I__4402 (
            .O(N__26995),
            .I(N__26956));
    Span4Mux_h I__4401 (
            .O(N__26992),
            .I(N__26953));
    LocalMux I__4400 (
            .O(N__26981),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    LocalMux I__4399 (
            .O(N__26970),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv12 I__4398 (
            .O(N__26959),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__4397 (
            .O(N__26956),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__4396 (
            .O(N__26953),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    CascadeMux I__4395 (
            .O(N__26942),
            .I(N__26939));
    InMux I__4394 (
            .O(N__26939),
            .I(N__26934));
    CascadeMux I__4393 (
            .O(N__26938),
            .I(N__26931));
    InMux I__4392 (
            .O(N__26937),
            .I(N__26927));
    LocalMux I__4391 (
            .O(N__26934),
            .I(N__26924));
    InMux I__4390 (
            .O(N__26931),
            .I(N__26921));
    InMux I__4389 (
            .O(N__26930),
            .I(N__26918));
    LocalMux I__4388 (
            .O(N__26927),
            .I(N__26915));
    Span4Mux_v I__4387 (
            .O(N__26924),
            .I(N__26910));
    LocalMux I__4386 (
            .O(N__26921),
            .I(N__26910));
    LocalMux I__4385 (
            .O(N__26918),
            .I(N__26903));
    Span4Mux_h I__4384 (
            .O(N__26915),
            .I(N__26903));
    Span4Mux_h I__4383 (
            .O(N__26910),
            .I(N__26903));
    Span4Mux_v I__4382 (
            .O(N__26903),
            .I(N__26899));
    InMux I__4381 (
            .O(N__26902),
            .I(N__26896));
    Odrv4 I__4380 (
            .O(N__26899),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__4379 (
            .O(N__26896),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    CascadeMux I__4378 (
            .O(N__26891),
            .I(N__26887));
    InMux I__4377 (
            .O(N__26890),
            .I(N__26884));
    InMux I__4376 (
            .O(N__26887),
            .I(N__26879));
    LocalMux I__4375 (
            .O(N__26884),
            .I(N__26876));
    InMux I__4374 (
            .O(N__26883),
            .I(N__26871));
    InMux I__4373 (
            .O(N__26882),
            .I(N__26871));
    LocalMux I__4372 (
            .O(N__26879),
            .I(elapsed_time_ns_1_RNIO0MD11_0_11));
    Odrv4 I__4371 (
            .O(N__26876),
            .I(elapsed_time_ns_1_RNIO0MD11_0_11));
    LocalMux I__4370 (
            .O(N__26871),
            .I(elapsed_time_ns_1_RNIO0MD11_0_11));
    CascadeMux I__4369 (
            .O(N__26864),
            .I(N__26860));
    InMux I__4368 (
            .O(N__26863),
            .I(N__26857));
    InMux I__4367 (
            .O(N__26860),
            .I(N__26854));
    LocalMux I__4366 (
            .O(N__26857),
            .I(N__26851));
    LocalMux I__4365 (
            .O(N__26854),
            .I(N__26848));
    Span4Mux_h I__4364 (
            .O(N__26851),
            .I(N__26842));
    Span4Mux_v I__4363 (
            .O(N__26848),
            .I(N__26842));
    InMux I__4362 (
            .O(N__26847),
            .I(N__26839));
    Odrv4 I__4361 (
            .O(N__26842),
            .I(elapsed_time_ns_1_RNIP1MD11_0_12));
    LocalMux I__4360 (
            .O(N__26839),
            .I(elapsed_time_ns_1_RNIP1MD11_0_12));
    InMux I__4359 (
            .O(N__26834),
            .I(N__26831));
    LocalMux I__4358 (
            .O(N__26831),
            .I(\current_shift_inst.PI_CTRL.integrator_i_10 ));
    InMux I__4357 (
            .O(N__26828),
            .I(N__26825));
    LocalMux I__4356 (
            .O(N__26825),
            .I(N__26822));
    Odrv12 I__4355 (
            .O(N__26822),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    CascadeMux I__4354 (
            .O(N__26819),
            .I(N__26816));
    InMux I__4353 (
            .O(N__26816),
            .I(N__26812));
    InMux I__4352 (
            .O(N__26815),
            .I(N__26808));
    LocalMux I__4351 (
            .O(N__26812),
            .I(N__26805));
    InMux I__4350 (
            .O(N__26811),
            .I(N__26800));
    LocalMux I__4349 (
            .O(N__26808),
            .I(N__26797));
    Span4Mux_h I__4348 (
            .O(N__26805),
            .I(N__26794));
    InMux I__4347 (
            .O(N__26804),
            .I(N__26791));
    InMux I__4346 (
            .O(N__26803),
            .I(N__26788));
    LocalMux I__4345 (
            .O(N__26800),
            .I(N__26785));
    Span4Mux_h I__4344 (
            .O(N__26797),
            .I(N__26778));
    Span4Mux_h I__4343 (
            .O(N__26794),
            .I(N__26778));
    LocalMux I__4342 (
            .O(N__26791),
            .I(N__26778));
    LocalMux I__4341 (
            .O(N__26788),
            .I(N__26775));
    Odrv12 I__4340 (
            .O(N__26785),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__4339 (
            .O(N__26778),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__4338 (
            .O(N__26775),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    InMux I__4337 (
            .O(N__26768),
            .I(N__26765));
    LocalMux I__4336 (
            .O(N__26765),
            .I(N__26762));
    Odrv4 I__4335 (
            .O(N__26762),
            .I(\current_shift_inst.PI_CTRL.integrator_i_20 ));
    InMux I__4334 (
            .O(N__26759),
            .I(N__26755));
    InMux I__4333 (
            .O(N__26758),
            .I(N__26751));
    LocalMux I__4332 (
            .O(N__26755),
            .I(N__26748));
    InMux I__4331 (
            .O(N__26754),
            .I(N__26745));
    LocalMux I__4330 (
            .O(N__26751),
            .I(N__26742));
    Span4Mux_h I__4329 (
            .O(N__26748),
            .I(N__26739));
    LocalMux I__4328 (
            .O(N__26745),
            .I(N__26736));
    Odrv12 I__4327 (
            .O(N__26742),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    Odrv4 I__4326 (
            .O(N__26739),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    Odrv12 I__4325 (
            .O(N__26736),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__4324 (
            .O(N__26729),
            .I(N__26726));
    LocalMux I__4323 (
            .O(N__26726),
            .I(N__26723));
    Odrv4 I__4322 (
            .O(N__26723),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ));
    InMux I__4321 (
            .O(N__26720),
            .I(N__26717));
    LocalMux I__4320 (
            .O(N__26717),
            .I(N__26714));
    Odrv12 I__4319 (
            .O(N__26714),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__4318 (
            .O(N__26711),
            .I(N__26707));
    InMux I__4317 (
            .O(N__26710),
            .I(N__26704));
    LocalMux I__4316 (
            .O(N__26707),
            .I(N__26698));
    LocalMux I__4315 (
            .O(N__26704),
            .I(N__26698));
    InMux I__4314 (
            .O(N__26703),
            .I(N__26695));
    Span4Mux_v I__4313 (
            .O(N__26698),
            .I(N__26692));
    LocalMux I__4312 (
            .O(N__26695),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    Odrv4 I__4311 (
            .O(N__26692),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    CascadeMux I__4310 (
            .O(N__26687),
            .I(N__26684));
    InMux I__4309 (
            .O(N__26684),
            .I(N__26681));
    LocalMux I__4308 (
            .O(N__26681),
            .I(N__26675));
    InMux I__4307 (
            .O(N__26680),
            .I(N__26672));
    InMux I__4306 (
            .O(N__26679),
            .I(N__26669));
    InMux I__4305 (
            .O(N__26678),
            .I(N__26665));
    Span4Mux_h I__4304 (
            .O(N__26675),
            .I(N__26658));
    LocalMux I__4303 (
            .O(N__26672),
            .I(N__26658));
    LocalMux I__4302 (
            .O(N__26669),
            .I(N__26658));
    InMux I__4301 (
            .O(N__26668),
            .I(N__26655));
    LocalMux I__4300 (
            .O(N__26665),
            .I(N__26650));
    Span4Mux_h I__4299 (
            .O(N__26658),
            .I(N__26650));
    LocalMux I__4298 (
            .O(N__26655),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__4297 (
            .O(N__26650),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__4296 (
            .O(N__26645),
            .I(N__26642));
    LocalMux I__4295 (
            .O(N__26642),
            .I(N__26639));
    Span4Mux_v I__4294 (
            .O(N__26639),
            .I(N__26634));
    InMux I__4293 (
            .O(N__26638),
            .I(N__26631));
    InMux I__4292 (
            .O(N__26637),
            .I(N__26628));
    Span4Mux_h I__4291 (
            .O(N__26634),
            .I(N__26625));
    LocalMux I__4290 (
            .O(N__26631),
            .I(N__26622));
    LocalMux I__4289 (
            .O(N__26628),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    Odrv4 I__4288 (
            .O(N__26625),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    Odrv12 I__4287 (
            .O(N__26622),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    InMux I__4286 (
            .O(N__26615),
            .I(N__26612));
    LocalMux I__4285 (
            .O(N__26612),
            .I(N__26609));
    Span4Mux_h I__4284 (
            .O(N__26609),
            .I(N__26606));
    Odrv4 I__4283 (
            .O(N__26606),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ));
    CascadeMux I__4282 (
            .O(N__26603),
            .I(N__26600));
    InMux I__4281 (
            .O(N__26600),
            .I(N__26597));
    LocalMux I__4280 (
            .O(N__26597),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0 ));
    InMux I__4279 (
            .O(N__26594),
            .I(N__26590));
    InMux I__4278 (
            .O(N__26593),
            .I(N__26587));
    LocalMux I__4277 (
            .O(N__26590),
            .I(N__26583));
    LocalMux I__4276 (
            .O(N__26587),
            .I(N__26580));
    InMux I__4275 (
            .O(N__26586),
            .I(N__26577));
    Span4Mux_h I__4274 (
            .O(N__26583),
            .I(N__26574));
    Span4Mux_v I__4273 (
            .O(N__26580),
            .I(N__26571));
    LocalMux I__4272 (
            .O(N__26577),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    Odrv4 I__4271 (
            .O(N__26574),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    Odrv4 I__4270 (
            .O(N__26571),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    CascadeMux I__4269 (
            .O(N__26564),
            .I(N__26560));
    InMux I__4268 (
            .O(N__26563),
            .I(N__26556));
    InMux I__4267 (
            .O(N__26560),
            .I(N__26553));
    CascadeMux I__4266 (
            .O(N__26559),
            .I(N__26550));
    LocalMux I__4265 (
            .O(N__26556),
            .I(N__26546));
    LocalMux I__4264 (
            .O(N__26553),
            .I(N__26543));
    InMux I__4263 (
            .O(N__26550),
            .I(N__26540));
    InMux I__4262 (
            .O(N__26549),
            .I(N__26537));
    Span4Mux_h I__4261 (
            .O(N__26546),
            .I(N__26534));
    Span4Mux_v I__4260 (
            .O(N__26543),
            .I(N__26528));
    LocalMux I__4259 (
            .O(N__26540),
            .I(N__26528));
    LocalMux I__4258 (
            .O(N__26537),
            .I(N__26523));
    Span4Mux_h I__4257 (
            .O(N__26534),
            .I(N__26523));
    InMux I__4256 (
            .O(N__26533),
            .I(N__26520));
    Span4Mux_h I__4255 (
            .O(N__26528),
            .I(N__26517));
    Odrv4 I__4254 (
            .O(N__26523),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__4253 (
            .O(N__26520),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__4252 (
            .O(N__26517),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    CascadeMux I__4251 (
            .O(N__26510),
            .I(N__26507));
    InMux I__4250 (
            .O(N__26507),
            .I(N__26504));
    LocalMux I__4249 (
            .O(N__26504),
            .I(N__26501));
    Span4Mux_h I__4248 (
            .O(N__26501),
            .I(N__26498));
    Odrv4 I__4247 (
            .O(N__26498),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ));
    CascadeMux I__4246 (
            .O(N__26495),
            .I(N__26492));
    InMux I__4245 (
            .O(N__26492),
            .I(N__26489));
    LocalMux I__4244 (
            .O(N__26489),
            .I(N__26486));
    Odrv4 I__4243 (
            .O(N__26486),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0 ));
    InMux I__4242 (
            .O(N__26483),
            .I(N__26480));
    LocalMux I__4241 (
            .O(N__26480),
            .I(N__26477));
    Odrv4 I__4240 (
            .O(N__26477),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    CascadeMux I__4239 (
            .O(N__26474),
            .I(N__26471));
    InMux I__4238 (
            .O(N__26471),
            .I(N__26468));
    LocalMux I__4237 (
            .O(N__26468),
            .I(N__26465));
    Odrv4 I__4236 (
            .O(N__26465),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__4235 (
            .O(N__26462),
            .I(N__26457));
    InMux I__4234 (
            .O(N__26461),
            .I(N__26454));
    InMux I__4233 (
            .O(N__26460),
            .I(N__26451));
    LocalMux I__4232 (
            .O(N__26457),
            .I(N__26448));
    LocalMux I__4231 (
            .O(N__26454),
            .I(N__26445));
    LocalMux I__4230 (
            .O(N__26451),
            .I(N__26442));
    Span4Mux_v I__4229 (
            .O(N__26448),
            .I(N__26439));
    Span4Mux_h I__4228 (
            .O(N__26445),
            .I(N__26436));
    Span4Mux_h I__4227 (
            .O(N__26442),
            .I(N__26433));
    Odrv4 I__4226 (
            .O(N__26439),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv4 I__4225 (
            .O(N__26436),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv4 I__4224 (
            .O(N__26433),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__4223 (
            .O(N__26426),
            .I(N__26423));
    LocalMux I__4222 (
            .O(N__26423),
            .I(N__26420));
    Span4Mux_h I__4221 (
            .O(N__26420),
            .I(N__26417));
    Odrv4 I__4220 (
            .O(N__26417),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ));
    CascadeMux I__4219 (
            .O(N__26414),
            .I(N__26411));
    InMux I__4218 (
            .O(N__26411),
            .I(N__26407));
    InMux I__4217 (
            .O(N__26410),
            .I(N__26404));
    LocalMux I__4216 (
            .O(N__26407),
            .I(N__26401));
    LocalMux I__4215 (
            .O(N__26404),
            .I(N__26397));
    Span4Mux_h I__4214 (
            .O(N__26401),
            .I(N__26394));
    InMux I__4213 (
            .O(N__26400),
            .I(N__26390));
    Span4Mux_h I__4212 (
            .O(N__26397),
            .I(N__26387));
    Span4Mux_h I__4211 (
            .O(N__26394),
            .I(N__26384));
    InMux I__4210 (
            .O(N__26393),
            .I(N__26381));
    LocalMux I__4209 (
            .O(N__26390),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__4208 (
            .O(N__26387),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__4207 (
            .O(N__26384),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__4206 (
            .O(N__26381),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    CascadeMux I__4205 (
            .O(N__26372),
            .I(N__26369));
    InMux I__4204 (
            .O(N__26369),
            .I(N__26366));
    LocalMux I__4203 (
            .O(N__26366),
            .I(\current_shift_inst.PI_CTRL.integrator_i_1 ));
    InMux I__4202 (
            .O(N__26363),
            .I(N__26360));
    LocalMux I__4201 (
            .O(N__26360),
            .I(\current_shift_inst.PI_CTRL.integrator_i_21 ));
    CascadeMux I__4200 (
            .O(N__26357),
            .I(N__26354));
    InMux I__4199 (
            .O(N__26354),
            .I(N__26350));
    InMux I__4198 (
            .O(N__26353),
            .I(N__26347));
    LocalMux I__4197 (
            .O(N__26350),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_12 ));
    LocalMux I__4196 (
            .O(N__26347),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_12 ));
    CascadeMux I__4195 (
            .O(N__26342),
            .I(N__26339));
    InMux I__4194 (
            .O(N__26339),
            .I(N__26335));
    InMux I__4193 (
            .O(N__26338),
            .I(N__26332));
    LocalMux I__4192 (
            .O(N__26335),
            .I(N__26328));
    LocalMux I__4191 (
            .O(N__26332),
            .I(N__26323));
    InMux I__4190 (
            .O(N__26331),
            .I(N__26320));
    Span4Mux_h I__4189 (
            .O(N__26328),
            .I(N__26317));
    InMux I__4188 (
            .O(N__26327),
            .I(N__26312));
    InMux I__4187 (
            .O(N__26326),
            .I(N__26312));
    Span4Mux_h I__4186 (
            .O(N__26323),
            .I(N__26309));
    LocalMux I__4185 (
            .O(N__26320),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__4184 (
            .O(N__26317),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__4183 (
            .O(N__26312),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__4182 (
            .O(N__26309),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__4181 (
            .O(N__26300),
            .I(N__26297));
    LocalMux I__4180 (
            .O(N__26297),
            .I(\current_shift_inst.PI_CTRL.integrator_i_14 ));
    InMux I__4179 (
            .O(N__26294),
            .I(N__26291));
    LocalMux I__4178 (
            .O(N__26291),
            .I(\current_shift_inst.PI_CTRL.integrator_i_22 ));
    InMux I__4177 (
            .O(N__26288),
            .I(N__26284));
    InMux I__4176 (
            .O(N__26287),
            .I(N__26280));
    LocalMux I__4175 (
            .O(N__26284),
            .I(N__26277));
    InMux I__4174 (
            .O(N__26283),
            .I(N__26274));
    LocalMux I__4173 (
            .O(N__26280),
            .I(N__26269));
    Span4Mux_h I__4172 (
            .O(N__26277),
            .I(N__26264));
    LocalMux I__4171 (
            .O(N__26274),
            .I(N__26264));
    InMux I__4170 (
            .O(N__26273),
            .I(N__26261));
    InMux I__4169 (
            .O(N__26272),
            .I(N__26258));
    Span4Mux_h I__4168 (
            .O(N__26269),
            .I(N__26253));
    Span4Mux_h I__4167 (
            .O(N__26264),
            .I(N__26253));
    LocalMux I__4166 (
            .O(N__26261),
            .I(N__26250));
    LocalMux I__4165 (
            .O(N__26258),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__4164 (
            .O(N__26253),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv12 I__4163 (
            .O(N__26250),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__4162 (
            .O(N__26243),
            .I(N__26240));
    LocalMux I__4161 (
            .O(N__26240),
            .I(\current_shift_inst.PI_CTRL.integrator_i_19 ));
    InMux I__4160 (
            .O(N__26237),
            .I(N__26234));
    LocalMux I__4159 (
            .O(N__26234),
            .I(N__26231));
    Odrv4 I__4158 (
            .O(N__26231),
            .I(\current_shift_inst.PI_CTRL.integrator_i_6 ));
    InMux I__4157 (
            .O(N__26228),
            .I(N__26225));
    LocalMux I__4156 (
            .O(N__26225),
            .I(N__26222));
    Span4Mux_v I__4155 (
            .O(N__26222),
            .I(N__26219));
    Odrv4 I__4154 (
            .O(N__26219),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    CascadeMux I__4153 (
            .O(N__26216),
            .I(N__26213));
    InMux I__4152 (
            .O(N__26213),
            .I(N__26209));
    InMux I__4151 (
            .O(N__26212),
            .I(N__26206));
    LocalMux I__4150 (
            .O(N__26209),
            .I(N__26203));
    LocalMux I__4149 (
            .O(N__26206),
            .I(N__26199));
    Span4Mux_h I__4148 (
            .O(N__26203),
            .I(N__26196));
    InMux I__4147 (
            .O(N__26202),
            .I(N__26193));
    Odrv12 I__4146 (
            .O(N__26199),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv4 I__4145 (
            .O(N__26196),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    LocalMux I__4144 (
            .O(N__26193),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__4143 (
            .O(N__26186),
            .I(N__26183));
    LocalMux I__4142 (
            .O(N__26183),
            .I(N__26180));
    Span4Mux_h I__4141 (
            .O(N__26180),
            .I(N__26177));
    Odrv4 I__4140 (
            .O(N__26177),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_9 ));
    CascadeMux I__4139 (
            .O(N__26174),
            .I(N__26171));
    InMux I__4138 (
            .O(N__26171),
            .I(N__26168));
    LocalMux I__4137 (
            .O(N__26168),
            .I(N__26165));
    Odrv4 I__4136 (
            .O(N__26165),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9 ));
    CascadeMux I__4135 (
            .O(N__26162),
            .I(N__26159));
    InMux I__4134 (
            .O(N__26159),
            .I(N__26156));
    LocalMux I__4133 (
            .O(N__26156),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    CascadeMux I__4132 (
            .O(N__26153),
            .I(N__26150));
    InMux I__4131 (
            .O(N__26150),
            .I(N__26146));
    InMux I__4130 (
            .O(N__26149),
            .I(N__26143));
    LocalMux I__4129 (
            .O(N__26146),
            .I(N__26139));
    LocalMux I__4128 (
            .O(N__26143),
            .I(N__26135));
    InMux I__4127 (
            .O(N__26142),
            .I(N__26131));
    Span4Mux_v I__4126 (
            .O(N__26139),
            .I(N__26128));
    InMux I__4125 (
            .O(N__26138),
            .I(N__26125));
    Span4Mux_h I__4124 (
            .O(N__26135),
            .I(N__26122));
    InMux I__4123 (
            .O(N__26134),
            .I(N__26119));
    LocalMux I__4122 (
            .O(N__26131),
            .I(N__26116));
    Span4Mux_h I__4121 (
            .O(N__26128),
            .I(N__26111));
    LocalMux I__4120 (
            .O(N__26125),
            .I(N__26111));
    Span4Mux_h I__4119 (
            .O(N__26122),
            .I(N__26108));
    LocalMux I__4118 (
            .O(N__26119),
            .I(N__26101));
    Span4Mux_v I__4117 (
            .O(N__26116),
            .I(N__26101));
    Span4Mux_h I__4116 (
            .O(N__26111),
            .I(N__26101));
    Odrv4 I__4115 (
            .O(N__26108),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__4114 (
            .O(N__26101),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__4113 (
            .O(N__26096),
            .I(N__26093));
    LocalMux I__4112 (
            .O(N__26093),
            .I(N__26090));
    Odrv4 I__4111 (
            .O(N__26090),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    CascadeMux I__4110 (
            .O(N__26087),
            .I(N__26084));
    InMux I__4109 (
            .O(N__26084),
            .I(N__26081));
    LocalMux I__4108 (
            .O(N__26081),
            .I(N__26078));
    Odrv4 I__4107 (
            .O(N__26078),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__4106 (
            .O(N__26075),
            .I(N__26070));
    InMux I__4105 (
            .O(N__26074),
            .I(N__26067));
    InMux I__4104 (
            .O(N__26073),
            .I(N__26064));
    LocalMux I__4103 (
            .O(N__26070),
            .I(N__26061));
    LocalMux I__4102 (
            .O(N__26067),
            .I(N__26054));
    LocalMux I__4101 (
            .O(N__26064),
            .I(N__26054));
    Span4Mux_h I__4100 (
            .O(N__26061),
            .I(N__26054));
    Odrv4 I__4099 (
            .O(N__26054),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__4098 (
            .O(N__26051),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__4097 (
            .O(N__26048),
            .I(N__26044));
    InMux I__4096 (
            .O(N__26047),
            .I(N__26040));
    LocalMux I__4095 (
            .O(N__26044),
            .I(N__26037));
    InMux I__4094 (
            .O(N__26043),
            .I(N__26034));
    LocalMux I__4093 (
            .O(N__26040),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__4092 (
            .O(N__26037),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__4091 (
            .O(N__26034),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__4090 (
            .O(N__26027),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__4089 (
            .O(N__26024),
            .I(N__26021));
    LocalMux I__4088 (
            .O(N__26021),
            .I(N__26016));
    InMux I__4087 (
            .O(N__26020),
            .I(N__26013));
    InMux I__4086 (
            .O(N__26019),
            .I(N__26010));
    Span4Mux_h I__4085 (
            .O(N__26016),
            .I(N__26007));
    LocalMux I__4084 (
            .O(N__26013),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__4083 (
            .O(N__26010),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__4082 (
            .O(N__26007),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__4081 (
            .O(N__26000),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__4080 (
            .O(N__25997),
            .I(N__25992));
    InMux I__4079 (
            .O(N__25996),
            .I(N__25989));
    InMux I__4078 (
            .O(N__25995),
            .I(N__25986));
    LocalMux I__4077 (
            .O(N__25992),
            .I(N__25983));
    LocalMux I__4076 (
            .O(N__25989),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__4075 (
            .O(N__25986),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__4074 (
            .O(N__25983),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__4073 (
            .O(N__25976),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__4072 (
            .O(N__25973),
            .I(N__25968));
    InMux I__4071 (
            .O(N__25972),
            .I(N__25965));
    InMux I__4070 (
            .O(N__25971),
            .I(N__25962));
    LocalMux I__4069 (
            .O(N__25968),
            .I(N__25959));
    LocalMux I__4068 (
            .O(N__25965),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__4067 (
            .O(N__25962),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv12 I__4066 (
            .O(N__25959),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__4065 (
            .O(N__25952),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__4064 (
            .O(N__25949),
            .I(N__25945));
    InMux I__4063 (
            .O(N__25948),
            .I(N__25941));
    LocalMux I__4062 (
            .O(N__25945),
            .I(N__25938));
    InMux I__4061 (
            .O(N__25944),
            .I(N__25935));
    LocalMux I__4060 (
            .O(N__25941),
            .I(N__25930));
    Span4Mux_h I__4059 (
            .O(N__25938),
            .I(N__25930));
    LocalMux I__4058 (
            .O(N__25935),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    Odrv4 I__4057 (
            .O(N__25930),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__4056 (
            .O(N__25925),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__4055 (
            .O(N__25922),
            .I(N__25917));
    InMux I__4054 (
            .O(N__25921),
            .I(N__25914));
    InMux I__4053 (
            .O(N__25920),
            .I(N__25911));
    LocalMux I__4052 (
            .O(N__25917),
            .I(N__25908));
    LocalMux I__4051 (
            .O(N__25914),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__4050 (
            .O(N__25911),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__4049 (
            .O(N__25908),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__4048 (
            .O(N__25901),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__4047 (
            .O(N__25898),
            .I(N__25894));
    InMux I__4046 (
            .O(N__25897),
            .I(N__25890));
    LocalMux I__4045 (
            .O(N__25894),
            .I(N__25887));
    InMux I__4044 (
            .O(N__25893),
            .I(N__25884));
    LocalMux I__4043 (
            .O(N__25890),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__4042 (
            .O(N__25887),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__4041 (
            .O(N__25884),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__4040 (
            .O(N__25877),
            .I(bfn_11_7_0_));
    InMux I__4039 (
            .O(N__25874),
            .I(N__25856));
    InMux I__4038 (
            .O(N__25873),
            .I(N__25856));
    InMux I__4037 (
            .O(N__25872),
            .I(N__25856));
    InMux I__4036 (
            .O(N__25871),
            .I(N__25856));
    InMux I__4035 (
            .O(N__25870),
            .I(N__25851));
    InMux I__4034 (
            .O(N__25869),
            .I(N__25851));
    InMux I__4033 (
            .O(N__25868),
            .I(N__25842));
    InMux I__4032 (
            .O(N__25867),
            .I(N__25842));
    InMux I__4031 (
            .O(N__25866),
            .I(N__25842));
    InMux I__4030 (
            .O(N__25865),
            .I(N__25842));
    LocalMux I__4029 (
            .O(N__25856),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__4028 (
            .O(N__25851),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__4027 (
            .O(N__25842),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__4026 (
            .O(N__25835),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__4025 (
            .O(N__25832),
            .I(N__25828));
    InMux I__4024 (
            .O(N__25831),
            .I(N__25824));
    LocalMux I__4023 (
            .O(N__25828),
            .I(N__25821));
    InMux I__4022 (
            .O(N__25827),
            .I(N__25818));
    LocalMux I__4021 (
            .O(N__25824),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__4020 (
            .O(N__25821),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__4019 (
            .O(N__25818),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__4018 (
            .O(N__25811),
            .I(N__25807));
    InMux I__4017 (
            .O(N__25810),
            .I(N__25804));
    LocalMux I__4016 (
            .O(N__25807),
            .I(N__25801));
    LocalMux I__4015 (
            .O(N__25804),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__4014 (
            .O(N__25801),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__4013 (
            .O(N__25796),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__4012 (
            .O(N__25793),
            .I(N__25789));
    InMux I__4011 (
            .O(N__25792),
            .I(N__25786));
    LocalMux I__4010 (
            .O(N__25789),
            .I(N__25783));
    LocalMux I__4009 (
            .O(N__25786),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__4008 (
            .O(N__25783),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__4007 (
            .O(N__25778),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__4006 (
            .O(N__25775),
            .I(N__25772));
    LocalMux I__4005 (
            .O(N__25772),
            .I(N__25768));
    InMux I__4004 (
            .O(N__25771),
            .I(N__25765));
    Span4Mux_h I__4003 (
            .O(N__25768),
            .I(N__25762));
    LocalMux I__4002 (
            .O(N__25765),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__4001 (
            .O(N__25762),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__4000 (
            .O(N__25757),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__3999 (
            .O(N__25754),
            .I(N__25750));
    InMux I__3998 (
            .O(N__25753),
            .I(N__25747));
    LocalMux I__3997 (
            .O(N__25750),
            .I(N__25744));
    LocalMux I__3996 (
            .O(N__25747),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv12 I__3995 (
            .O(N__25744),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__3994 (
            .O(N__25739),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__3993 (
            .O(N__25736),
            .I(N__25732));
    InMux I__3992 (
            .O(N__25735),
            .I(N__25729));
    LocalMux I__3991 (
            .O(N__25732),
            .I(N__25726));
    LocalMux I__3990 (
            .O(N__25729),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__3989 (
            .O(N__25726),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__3988 (
            .O(N__25721),
            .I(bfn_10_26_0_));
    InMux I__3987 (
            .O(N__25718),
            .I(N__25714));
    InMux I__3986 (
            .O(N__25717),
            .I(N__25711));
    LocalMux I__3985 (
            .O(N__25714),
            .I(N__25708));
    LocalMux I__3984 (
            .O(N__25711),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__3983 (
            .O(N__25708),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__3982 (
            .O(N__25703),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__3981 (
            .O(N__25700),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__3980 (
            .O(N__25697),
            .I(N__25693));
    InMux I__3979 (
            .O(N__25696),
            .I(N__25690));
    LocalMux I__3978 (
            .O(N__25693),
            .I(N__25687));
    LocalMux I__3977 (
            .O(N__25690),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__3976 (
            .O(N__25687),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__3975 (
            .O(N__25682),
            .I(N__25678));
    InMux I__3974 (
            .O(N__25681),
            .I(N__25674));
    LocalMux I__3973 (
            .O(N__25678),
            .I(N__25671));
    InMux I__3972 (
            .O(N__25677),
            .I(N__25668));
    LocalMux I__3971 (
            .O(N__25674),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__3970 (
            .O(N__25671),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__3969 (
            .O(N__25668),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__3968 (
            .O(N__25661),
            .I(bfn_11_6_0_));
    InMux I__3967 (
            .O(N__25658),
            .I(N__25654));
    InMux I__3966 (
            .O(N__25657),
            .I(N__25651));
    LocalMux I__3965 (
            .O(N__25654),
            .I(N__25648));
    LocalMux I__3964 (
            .O(N__25651),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv4 I__3963 (
            .O(N__25648),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__3962 (
            .O(N__25643),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__3961 (
            .O(N__25640),
            .I(N__25636));
    InMux I__3960 (
            .O(N__25639),
            .I(N__25633));
    LocalMux I__3959 (
            .O(N__25636),
            .I(N__25630));
    LocalMux I__3958 (
            .O(N__25633),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv4 I__3957 (
            .O(N__25630),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__3956 (
            .O(N__25625),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__3955 (
            .O(N__25622),
            .I(N__25618));
    InMux I__3954 (
            .O(N__25621),
            .I(N__25615));
    LocalMux I__3953 (
            .O(N__25618),
            .I(N__25612));
    LocalMux I__3952 (
            .O(N__25615),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv12 I__3951 (
            .O(N__25612),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__3950 (
            .O(N__25607),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__3949 (
            .O(N__25604),
            .I(N__25600));
    InMux I__3948 (
            .O(N__25603),
            .I(N__25597));
    LocalMux I__3947 (
            .O(N__25600),
            .I(N__25594));
    LocalMux I__3946 (
            .O(N__25597),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv12 I__3945 (
            .O(N__25594),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__3944 (
            .O(N__25589),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__3943 (
            .O(N__25586),
            .I(N__25582));
    InMux I__3942 (
            .O(N__25585),
            .I(N__25579));
    LocalMux I__3941 (
            .O(N__25582),
            .I(N__25576));
    LocalMux I__3940 (
            .O(N__25579),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__3939 (
            .O(N__25576),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__3938 (
            .O(N__25571),
            .I(bfn_10_25_0_));
    InMux I__3937 (
            .O(N__25568),
            .I(N__25564));
    InMux I__3936 (
            .O(N__25567),
            .I(N__25561));
    LocalMux I__3935 (
            .O(N__25564),
            .I(N__25558));
    LocalMux I__3934 (
            .O(N__25561),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv4 I__3933 (
            .O(N__25558),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__3932 (
            .O(N__25553),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__3931 (
            .O(N__25550),
            .I(N__25546));
    InMux I__3930 (
            .O(N__25549),
            .I(N__25543));
    LocalMux I__3929 (
            .O(N__25546),
            .I(N__25540));
    LocalMux I__3928 (
            .O(N__25543),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__3927 (
            .O(N__25540),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__3926 (
            .O(N__25535),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__3925 (
            .O(N__25532),
            .I(N__25528));
    InMux I__3924 (
            .O(N__25531),
            .I(N__25525));
    LocalMux I__3923 (
            .O(N__25528),
            .I(N__25522));
    LocalMux I__3922 (
            .O(N__25525),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__3921 (
            .O(N__25522),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__3920 (
            .O(N__25517),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__3919 (
            .O(N__25514),
            .I(N__25511));
    LocalMux I__3918 (
            .O(N__25511),
            .I(\phase_controller_inst2.stoper_hc.un6_running_19 ));
    CascadeMux I__3917 (
            .O(N__25508),
            .I(N__25505));
    InMux I__3916 (
            .O(N__25505),
            .I(N__25502));
    LocalMux I__3915 (
            .O(N__25502),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_19 ));
    InMux I__3914 (
            .O(N__25499),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_19 ));
    CascadeMux I__3913 (
            .O(N__25496),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    InMux I__3912 (
            .O(N__25493),
            .I(N__25490));
    LocalMux I__3911 (
            .O(N__25490),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ));
    InMux I__3910 (
            .O(N__25487),
            .I(N__25483));
    InMux I__3909 (
            .O(N__25486),
            .I(N__25480));
    LocalMux I__3908 (
            .O(N__25483),
            .I(N__25477));
    LocalMux I__3907 (
            .O(N__25480),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__3906 (
            .O(N__25477),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__3905 (
            .O(N__25472),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__3904 (
            .O(N__25469),
            .I(N__25466));
    InMux I__3903 (
            .O(N__25466),
            .I(N__25463));
    LocalMux I__3902 (
            .O(N__25463),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJBZ0Z21 ));
    InMux I__3901 (
            .O(N__25460),
            .I(N__25456));
    InMux I__3900 (
            .O(N__25459),
            .I(N__25453));
    LocalMux I__3899 (
            .O(N__25456),
            .I(N__25450));
    LocalMux I__3898 (
            .O(N__25453),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__3897 (
            .O(N__25450),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__3896 (
            .O(N__25445),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__3895 (
            .O(N__25442),
            .I(N__25438));
    InMux I__3894 (
            .O(N__25441),
            .I(N__25435));
    LocalMux I__3893 (
            .O(N__25438),
            .I(N__25432));
    LocalMux I__3892 (
            .O(N__25435),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv4 I__3891 (
            .O(N__25432),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__3890 (
            .O(N__25427),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__3889 (
            .O(N__25424),
            .I(N__25421));
    LocalMux I__3888 (
            .O(N__25421),
            .I(\phase_controller_inst2.stoper_hc.un6_running_11 ));
    CascadeMux I__3887 (
            .O(N__25418),
            .I(N__25415));
    InMux I__3886 (
            .O(N__25415),
            .I(N__25412));
    LocalMux I__3885 (
            .O(N__25412),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__3884 (
            .O(N__25409),
            .I(N__25406));
    InMux I__3883 (
            .O(N__25406),
            .I(N__25403));
    LocalMux I__3882 (
            .O(N__25403),
            .I(\phase_controller_inst2.stoper_hc.un6_running_12 ));
    InMux I__3881 (
            .O(N__25400),
            .I(N__25397));
    LocalMux I__3880 (
            .O(N__25397),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    InMux I__3879 (
            .O(N__25394),
            .I(N__25391));
    LocalMux I__3878 (
            .O(N__25391),
            .I(\phase_controller_inst2.stoper_hc.un6_running_13 ));
    CascadeMux I__3877 (
            .O(N__25388),
            .I(N__25385));
    InMux I__3876 (
            .O(N__25385),
            .I(N__25382));
    LocalMux I__3875 (
            .O(N__25382),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__3874 (
            .O(N__25379),
            .I(N__25376));
    LocalMux I__3873 (
            .O(N__25376),
            .I(\phase_controller_inst2.stoper_hc.un6_running_14 ));
    CascadeMux I__3872 (
            .O(N__25373),
            .I(N__25370));
    InMux I__3871 (
            .O(N__25370),
            .I(N__25367));
    LocalMux I__3870 (
            .O(N__25367),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    InMux I__3869 (
            .O(N__25364),
            .I(N__25361));
    LocalMux I__3868 (
            .O(N__25361),
            .I(\phase_controller_inst2.stoper_hc.un6_running_15 ));
    CascadeMux I__3867 (
            .O(N__25358),
            .I(N__25355));
    InMux I__3866 (
            .O(N__25355),
            .I(N__25352));
    LocalMux I__3865 (
            .O(N__25352),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__3864 (
            .O(N__25349),
            .I(N__25346));
    LocalMux I__3863 (
            .O(N__25346),
            .I(\phase_controller_inst2.stoper_hc.un6_running_16 ));
    CascadeMux I__3862 (
            .O(N__25343),
            .I(N__25340));
    InMux I__3861 (
            .O(N__25340),
            .I(N__25337));
    LocalMux I__3860 (
            .O(N__25337),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_16 ));
    CascadeMux I__3859 (
            .O(N__25334),
            .I(N__25331));
    InMux I__3858 (
            .O(N__25331),
            .I(N__25328));
    LocalMux I__3857 (
            .O(N__25328),
            .I(\phase_controller_inst2.stoper_hc.un6_running_17 ));
    InMux I__3856 (
            .O(N__25325),
            .I(N__25322));
    LocalMux I__3855 (
            .O(N__25322),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_17 ));
    InMux I__3854 (
            .O(N__25319),
            .I(N__25316));
    LocalMux I__3853 (
            .O(N__25316),
            .I(\phase_controller_inst2.stoper_hc.un6_running_18 ));
    CascadeMux I__3852 (
            .O(N__25313),
            .I(N__25310));
    InMux I__3851 (
            .O(N__25310),
            .I(N__25307));
    LocalMux I__3850 (
            .O(N__25307),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_18 ));
    InMux I__3849 (
            .O(N__25304),
            .I(N__25301));
    LocalMux I__3848 (
            .O(N__25301),
            .I(N__25298));
    Odrv4 I__3847 (
            .O(N__25298),
            .I(\phase_controller_inst2.stoper_hc.un6_running_3 ));
    CascadeMux I__3846 (
            .O(N__25295),
            .I(N__25292));
    InMux I__3845 (
            .O(N__25292),
            .I(N__25289));
    LocalMux I__3844 (
            .O(N__25289),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__3843 (
            .O(N__25286),
            .I(N__25283));
    LocalMux I__3842 (
            .O(N__25283),
            .I(N__25280));
    Odrv4 I__3841 (
            .O(N__25280),
            .I(\phase_controller_inst2.stoper_hc.un6_running_4 ));
    CascadeMux I__3840 (
            .O(N__25277),
            .I(N__25274));
    InMux I__3839 (
            .O(N__25274),
            .I(N__25271));
    LocalMux I__3838 (
            .O(N__25271),
            .I(N__25268));
    Odrv4 I__3837 (
            .O(N__25268),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__3836 (
            .O(N__25265),
            .I(N__25262));
    LocalMux I__3835 (
            .O(N__25262),
            .I(N__25259));
    Odrv4 I__3834 (
            .O(N__25259),
            .I(\phase_controller_inst2.stoper_hc.un6_running_5 ));
    CascadeMux I__3833 (
            .O(N__25256),
            .I(N__25253));
    InMux I__3832 (
            .O(N__25253),
            .I(N__25250));
    LocalMux I__3831 (
            .O(N__25250),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    InMux I__3830 (
            .O(N__25247),
            .I(N__25244));
    LocalMux I__3829 (
            .O(N__25244),
            .I(N__25241));
    Odrv4 I__3828 (
            .O(N__25241),
            .I(\phase_controller_inst2.stoper_hc.un6_running_6 ));
    CascadeMux I__3827 (
            .O(N__25238),
            .I(N__25235));
    InMux I__3826 (
            .O(N__25235),
            .I(N__25232));
    LocalMux I__3825 (
            .O(N__25232),
            .I(N__25229));
    Odrv4 I__3824 (
            .O(N__25229),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    InMux I__3823 (
            .O(N__25226),
            .I(N__25223));
    LocalMux I__3822 (
            .O(N__25223),
            .I(N__25220));
    Odrv4 I__3821 (
            .O(N__25220),
            .I(\phase_controller_inst2.stoper_hc.un6_running_7 ));
    CascadeMux I__3820 (
            .O(N__25217),
            .I(N__25214));
    InMux I__3819 (
            .O(N__25214),
            .I(N__25211));
    LocalMux I__3818 (
            .O(N__25211),
            .I(N__25208));
    Odrv4 I__3817 (
            .O(N__25208),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    CascadeMux I__3816 (
            .O(N__25205),
            .I(N__25202));
    InMux I__3815 (
            .O(N__25202),
            .I(N__25199));
    LocalMux I__3814 (
            .O(N__25199),
            .I(N__25196));
    Odrv4 I__3813 (
            .O(N__25196),
            .I(\phase_controller_inst2.stoper_hc.un6_running_8 ));
    InMux I__3812 (
            .O(N__25193),
            .I(N__25190));
    LocalMux I__3811 (
            .O(N__25190),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    InMux I__3810 (
            .O(N__25187),
            .I(N__25184));
    LocalMux I__3809 (
            .O(N__25184),
            .I(N__25181));
    Span4Mux_v I__3808 (
            .O(N__25181),
            .I(N__25178));
    Span4Mux_h I__3807 (
            .O(N__25178),
            .I(N__25175));
    Odrv4 I__3806 (
            .O(N__25175),
            .I(\phase_controller_inst2.stoper_hc.un6_running_9 ));
    CascadeMux I__3805 (
            .O(N__25172),
            .I(N__25169));
    InMux I__3804 (
            .O(N__25169),
            .I(N__25166));
    LocalMux I__3803 (
            .O(N__25166),
            .I(N__25163));
    Odrv4 I__3802 (
            .O(N__25163),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__3801 (
            .O(N__25160),
            .I(N__25157));
    LocalMux I__3800 (
            .O(N__25157),
            .I(\phase_controller_inst2.stoper_hc.un6_running_10 ));
    CascadeMux I__3799 (
            .O(N__25154),
            .I(N__25151));
    InMux I__3798 (
            .O(N__25151),
            .I(N__25148));
    LocalMux I__3797 (
            .O(N__25148),
            .I(N__25145));
    Odrv4 I__3796 (
            .O(N__25145),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    InMux I__3795 (
            .O(N__25142),
            .I(N__25139));
    LocalMux I__3794 (
            .O(N__25139),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15 ));
    InMux I__3793 (
            .O(N__25136),
            .I(N__25132));
    InMux I__3792 (
            .O(N__25135),
            .I(N__25129));
    LocalMux I__3791 (
            .O(N__25132),
            .I(elapsed_time_ns_1_RNI0AND11_0_28));
    LocalMux I__3790 (
            .O(N__25129),
            .I(elapsed_time_ns_1_RNI0AND11_0_28));
    InMux I__3789 (
            .O(N__25124),
            .I(N__25121));
    LocalMux I__3788 (
            .O(N__25121),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15 ));
    InMux I__3787 (
            .O(N__25118),
            .I(N__25112));
    InMux I__3786 (
            .O(N__25117),
            .I(N__25112));
    LocalMux I__3785 (
            .O(N__25112),
            .I(elapsed_time_ns_1_RNI1BND11_0_29));
    InMux I__3784 (
            .O(N__25109),
            .I(N__25105));
    InMux I__3783 (
            .O(N__25108),
            .I(N__25102));
    LocalMux I__3782 (
            .O(N__25105),
            .I(elapsed_time_ns_1_RNIO1ND11_0_20));
    LocalMux I__3781 (
            .O(N__25102),
            .I(elapsed_time_ns_1_RNIO1ND11_0_20));
    CascadeMux I__3780 (
            .O(N__25097),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15_cascade_ ));
    InMux I__3779 (
            .O(N__25094),
            .I(N__25088));
    InMux I__3778 (
            .O(N__25093),
            .I(N__25088));
    LocalMux I__3777 (
            .O(N__25088),
            .I(elapsed_time_ns_1_RNIV8ND11_0_27));
    CascadeMux I__3776 (
            .O(N__25085),
            .I(N__25082));
    InMux I__3775 (
            .O(N__25082),
            .I(N__25079));
    LocalMux I__3774 (
            .O(N__25079),
            .I(N__25076));
    Odrv4 I__3773 (
            .O(N__25076),
            .I(\phase_controller_inst2.stoper_hc.un6_running_1 ));
    InMux I__3772 (
            .O(N__25073),
            .I(N__25070));
    LocalMux I__3771 (
            .O(N__25070),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    InMux I__3770 (
            .O(N__25067),
            .I(N__25064));
    LocalMux I__3769 (
            .O(N__25064),
            .I(N__25061));
    Odrv4 I__3768 (
            .O(N__25061),
            .I(\phase_controller_inst2.stoper_hc.un6_running_2 ));
    CascadeMux I__3767 (
            .O(N__25058),
            .I(N__25055));
    InMux I__3766 (
            .O(N__25055),
            .I(N__25052));
    LocalMux I__3765 (
            .O(N__25052),
            .I(N__25049));
    Odrv4 I__3764 (
            .O(N__25049),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__3763 (
            .O(N__25046),
            .I(N__25043));
    InMux I__3762 (
            .O(N__25043),
            .I(N__25039));
    InMux I__3761 (
            .O(N__25042),
            .I(N__25035));
    LocalMux I__3760 (
            .O(N__25039),
            .I(N__25032));
    InMux I__3759 (
            .O(N__25038),
            .I(N__25028));
    LocalMux I__3758 (
            .O(N__25035),
            .I(N__25023));
    Span4Mux_v I__3757 (
            .O(N__25032),
            .I(N__25023));
    InMux I__3756 (
            .O(N__25031),
            .I(N__25020));
    LocalMux I__3755 (
            .O(N__25028),
            .I(elapsed_time_ns_1_RNINVLD11_0_10));
    Odrv4 I__3754 (
            .O(N__25023),
            .I(elapsed_time_ns_1_RNINVLD11_0_10));
    LocalMux I__3753 (
            .O(N__25020),
            .I(elapsed_time_ns_1_RNINVLD11_0_10));
    InMux I__3752 (
            .O(N__25013),
            .I(N__25010));
    LocalMux I__3751 (
            .O(N__25010),
            .I(elapsed_time_ns_1_RNIP2ND11_0_21));
    CascadeMux I__3750 (
            .O(N__25007),
            .I(elapsed_time_ns_1_RNIP2ND11_0_21_cascade_));
    CascadeMux I__3749 (
            .O(N__25004),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15_cascade_ ));
    InMux I__3748 (
            .O(N__25001),
            .I(N__24995));
    InMux I__3747 (
            .O(N__25000),
            .I(N__24995));
    LocalMux I__3746 (
            .O(N__24995),
            .I(elapsed_time_ns_1_RNIU7ND11_0_26));
    InMux I__3745 (
            .O(N__24992),
            .I(N__24989));
    LocalMux I__3744 (
            .O(N__24989),
            .I(elapsed_time_ns_1_RNIR4ND11_0_23));
    CascadeMux I__3743 (
            .O(N__24986),
            .I(elapsed_time_ns_1_RNIR4ND11_0_23_cascade_));
    CascadeMux I__3742 (
            .O(N__24983),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_ ));
    CascadeMux I__3741 (
            .O(N__24980),
            .I(elapsed_time_ns_1_RNIP1MD11_0_12_cascade_));
    InMux I__3740 (
            .O(N__24977),
            .I(N__24972));
    InMux I__3739 (
            .O(N__24976),
            .I(N__24969));
    InMux I__3738 (
            .O(N__24975),
            .I(N__24966));
    LocalMux I__3737 (
            .O(N__24972),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2 ));
    LocalMux I__3736 (
            .O(N__24969),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2 ));
    LocalMux I__3735 (
            .O(N__24966),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2 ));
    InMux I__3734 (
            .O(N__24959),
            .I(N__24954));
    InMux I__3733 (
            .O(N__24958),
            .I(N__24949));
    InMux I__3732 (
            .O(N__24957),
            .I(N__24949));
    LocalMux I__3731 (
            .O(N__24954),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ));
    LocalMux I__3730 (
            .O(N__24949),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ));
    CascadeMux I__3729 (
            .O(N__24944),
            .I(N__24940));
    CascadeMux I__3728 (
            .O(N__24943),
            .I(N__24936));
    InMux I__3727 (
            .O(N__24940),
            .I(N__24933));
    InMux I__3726 (
            .O(N__24939),
            .I(N__24928));
    InMux I__3725 (
            .O(N__24936),
            .I(N__24928));
    LocalMux I__3724 (
            .O(N__24933),
            .I(N__24925));
    LocalMux I__3723 (
            .O(N__24928),
            .I(N__24922));
    Span4Mux_h I__3722 (
            .O(N__24925),
            .I(N__24919));
    Odrv4 I__3721 (
            .O(N__24922),
            .I(\phase_controller_inst1.stoper_hc.N_337 ));
    Odrv4 I__3720 (
            .O(N__24919),
            .I(\phase_controller_inst1.stoper_hc.N_337 ));
    InMux I__3719 (
            .O(N__24914),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ));
    CascadeMux I__3718 (
            .O(N__24911),
            .I(N__24908));
    InMux I__3717 (
            .O(N__24908),
            .I(N__24905));
    LocalMux I__3716 (
            .O(N__24905),
            .I(N__24902));
    Odrv4 I__3715 (
            .O(N__24902),
            .I(\current_shift_inst.PI_CTRL.integrator_i_29 ));
    InMux I__3714 (
            .O(N__24899),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ));
    InMux I__3713 (
            .O(N__24896),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ));
    InMux I__3712 (
            .O(N__24893),
            .I(bfn_10_17_0_));
    InMux I__3711 (
            .O(N__24890),
            .I(N__24887));
    LocalMux I__3710 (
            .O(N__24887),
            .I(\current_shift_inst.PI_CTRL.integrator_i_23 ));
    InMux I__3709 (
            .O(N__24884),
            .I(N__24875));
    InMux I__3708 (
            .O(N__24883),
            .I(N__24875));
    InMux I__3707 (
            .O(N__24882),
            .I(N__24872));
    InMux I__3706 (
            .O(N__24881),
            .I(N__24869));
    InMux I__3705 (
            .O(N__24880),
            .I(N__24866));
    LocalMux I__3704 (
            .O(N__24875),
            .I(N__24863));
    LocalMux I__3703 (
            .O(N__24872),
            .I(N__24860));
    LocalMux I__3702 (
            .O(N__24869),
            .I(N__24855));
    LocalMux I__3701 (
            .O(N__24866),
            .I(N__24855));
    Span4Mux_h I__3700 (
            .O(N__24863),
            .I(N__24852));
    Span4Mux_h I__3699 (
            .O(N__24860),
            .I(N__24847));
    Span4Mux_h I__3698 (
            .O(N__24855),
            .I(N__24847));
    Odrv4 I__3697 (
            .O(N__24852),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__3696 (
            .O(N__24847),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    CascadeMux I__3695 (
            .O(N__24842),
            .I(N__24839));
    InMux I__3694 (
            .O(N__24839),
            .I(N__24836));
    LocalMux I__3693 (
            .O(N__24836),
            .I(N__24833));
    Span4Mux_h I__3692 (
            .O(N__24833),
            .I(N__24830));
    Odrv4 I__3691 (
            .O(N__24830),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ));
    InMux I__3690 (
            .O(N__24827),
            .I(N__24823));
    InMux I__3689 (
            .O(N__24826),
            .I(N__24819));
    LocalMux I__3688 (
            .O(N__24823),
            .I(N__24816));
    InMux I__3687 (
            .O(N__24822),
            .I(N__24813));
    LocalMux I__3686 (
            .O(N__24819),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    Odrv12 I__3685 (
            .O(N__24816),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    LocalMux I__3684 (
            .O(N__24813),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    CascadeMux I__3683 (
            .O(N__24806),
            .I(N__24803));
    InMux I__3682 (
            .O(N__24803),
            .I(N__24800));
    LocalMux I__3681 (
            .O(N__24800),
            .I(N__24797));
    Odrv4 I__3680 (
            .O(N__24797),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0 ));
    CascadeMux I__3679 (
            .O(N__24794),
            .I(N__24791));
    InMux I__3678 (
            .O(N__24791),
            .I(N__24788));
    LocalMux I__3677 (
            .O(N__24788),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0 ));
    InMux I__3676 (
            .O(N__24785),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ));
    InMux I__3675 (
            .O(N__24782),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ));
    InMux I__3674 (
            .O(N__24779),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ));
    InMux I__3673 (
            .O(N__24776),
            .I(N__24773));
    LocalMux I__3672 (
            .O(N__24773),
            .I(N__24770));
    Span4Mux_h I__3671 (
            .O(N__24770),
            .I(N__24767));
    Odrv4 I__3670 (
            .O(N__24767),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__3669 (
            .O(N__24764),
            .I(bfn_10_16_0_));
    InMux I__3668 (
            .O(N__24761),
            .I(N__24758));
    LocalMux I__3667 (
            .O(N__24758),
            .I(N__24755));
    Span4Mux_h I__3666 (
            .O(N__24755),
            .I(N__24752));
    Odrv4 I__3665 (
            .O(N__24752),
            .I(\current_shift_inst.PI_CTRL.integrator_i_24 ));
    CascadeMux I__3664 (
            .O(N__24749),
            .I(N__24746));
    InMux I__3663 (
            .O(N__24746),
            .I(N__24743));
    LocalMux I__3662 (
            .O(N__24743),
            .I(N__24740));
    Odrv4 I__3661 (
            .O(N__24740),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0 ));
    CascadeMux I__3660 (
            .O(N__24737),
            .I(N__24734));
    InMux I__3659 (
            .O(N__24734),
            .I(N__24731));
    LocalMux I__3658 (
            .O(N__24731),
            .I(N__24728));
    Span4Mux_v I__3657 (
            .O(N__24728),
            .I(N__24725));
    Odrv4 I__3656 (
            .O(N__24725),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__3655 (
            .O(N__24722),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ));
    InMux I__3654 (
            .O(N__24719),
            .I(N__24716));
    LocalMux I__3653 (
            .O(N__24716),
            .I(N__24713));
    Span4Mux_v I__3652 (
            .O(N__24713),
            .I(N__24710));
    Odrv4 I__3651 (
            .O(N__24710),
            .I(\current_shift_inst.PI_CTRL.integrator_i_25 ));
    CascadeMux I__3650 (
            .O(N__24707),
            .I(N__24704));
    InMux I__3649 (
            .O(N__24704),
            .I(N__24701));
    LocalMux I__3648 (
            .O(N__24701),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0 ));
    InMux I__3647 (
            .O(N__24698),
            .I(N__24695));
    LocalMux I__3646 (
            .O(N__24695),
            .I(N__24692));
    Span4Mux_v I__3645 (
            .O(N__24692),
            .I(N__24689));
    Odrv4 I__3644 (
            .O(N__24689),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__3643 (
            .O(N__24686),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ));
    InMux I__3642 (
            .O(N__24683),
            .I(N__24680));
    LocalMux I__3641 (
            .O(N__24680),
            .I(N__24677));
    Span12Mux_h I__3640 (
            .O(N__24677),
            .I(N__24674));
    Odrv12 I__3639 (
            .O(N__24674),
            .I(\current_shift_inst.PI_CTRL.integrator_i_26 ));
    CascadeMux I__3638 (
            .O(N__24671),
            .I(N__24668));
    InMux I__3637 (
            .O(N__24668),
            .I(N__24665));
    LocalMux I__3636 (
            .O(N__24665),
            .I(N__24662));
    Odrv4 I__3635 (
            .O(N__24662),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0 ));
    CascadeMux I__3634 (
            .O(N__24659),
            .I(N__24656));
    InMux I__3633 (
            .O(N__24656),
            .I(N__24653));
    LocalMux I__3632 (
            .O(N__24653),
            .I(N__24650));
    Span4Mux_v I__3631 (
            .O(N__24650),
            .I(N__24647));
    Odrv4 I__3630 (
            .O(N__24647),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__3629 (
            .O(N__24644),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ));
    CascadeMux I__3628 (
            .O(N__24641),
            .I(N__24638));
    InMux I__3627 (
            .O(N__24638),
            .I(N__24635));
    LocalMux I__3626 (
            .O(N__24635),
            .I(N__24632));
    Span4Mux_h I__3625 (
            .O(N__24632),
            .I(N__24629));
    Odrv4 I__3624 (
            .O(N__24629),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0 ));
    CascadeMux I__3623 (
            .O(N__24626),
            .I(N__24623));
    InMux I__3622 (
            .O(N__24623),
            .I(N__24620));
    LocalMux I__3621 (
            .O(N__24620),
            .I(N__24617));
    Odrv12 I__3620 (
            .O(N__24617),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__3619 (
            .O(N__24614),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ));
    InMux I__3618 (
            .O(N__24611),
            .I(N__24608));
    LocalMux I__3617 (
            .O(N__24608),
            .I(N__24605));
    Odrv4 I__3616 (
            .O(N__24605),
            .I(\current_shift_inst.PI_CTRL.integrator_i_12 ));
    CascadeMux I__3615 (
            .O(N__24602),
            .I(N__24599));
    InMux I__3614 (
            .O(N__24599),
            .I(N__24596));
    LocalMux I__3613 (
            .O(N__24596),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0 ));
    InMux I__3612 (
            .O(N__24593),
            .I(N__24590));
    LocalMux I__3611 (
            .O(N__24590),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__3610 (
            .O(N__24587),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ));
    InMux I__3609 (
            .O(N__24584),
            .I(N__24581));
    LocalMux I__3608 (
            .O(N__24581),
            .I(N__24578));
    Odrv4 I__3607 (
            .O(N__24578),
            .I(\current_shift_inst.PI_CTRL.integrator_i_13 ));
    CascadeMux I__3606 (
            .O(N__24575),
            .I(N__24572));
    InMux I__3605 (
            .O(N__24572),
            .I(N__24569));
    LocalMux I__3604 (
            .O(N__24569),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0 ));
    InMux I__3603 (
            .O(N__24566),
            .I(N__24563));
    LocalMux I__3602 (
            .O(N__24563),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__3601 (
            .O(N__24560),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ));
    CascadeMux I__3600 (
            .O(N__24557),
            .I(N__24554));
    InMux I__3599 (
            .O(N__24554),
            .I(N__24551));
    LocalMux I__3598 (
            .O(N__24551),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0 ));
    InMux I__3597 (
            .O(N__24548),
            .I(N__24545));
    LocalMux I__3596 (
            .O(N__24545),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__3595 (
            .O(N__24542),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ));
    InMux I__3594 (
            .O(N__24539),
            .I(N__24536));
    LocalMux I__3593 (
            .O(N__24536),
            .I(N__24533));
    Span4Mux_h I__3592 (
            .O(N__24533),
            .I(N__24530));
    Odrv4 I__3591 (
            .O(N__24530),
            .I(\current_shift_inst.PI_CTRL.integrator_i_15 ));
    CascadeMux I__3590 (
            .O(N__24527),
            .I(N__24524));
    InMux I__3589 (
            .O(N__24524),
            .I(N__24521));
    LocalMux I__3588 (
            .O(N__24521),
            .I(N__24518));
    Odrv4 I__3587 (
            .O(N__24518),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0 ));
    CascadeMux I__3586 (
            .O(N__24515),
            .I(N__24512));
    InMux I__3585 (
            .O(N__24512),
            .I(N__24509));
    LocalMux I__3584 (
            .O(N__24509),
            .I(N__24506));
    Span4Mux_v I__3583 (
            .O(N__24506),
            .I(N__24503));
    Odrv4 I__3582 (
            .O(N__24503),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__3581 (
            .O(N__24500),
            .I(bfn_10_15_0_));
    InMux I__3580 (
            .O(N__24497),
            .I(N__24494));
    LocalMux I__3579 (
            .O(N__24494),
            .I(N__24491));
    Span4Mux_h I__3578 (
            .O(N__24491),
            .I(N__24488));
    Odrv4 I__3577 (
            .O(N__24488),
            .I(\current_shift_inst.PI_CTRL.integrator_i_16 ));
    CascadeMux I__3576 (
            .O(N__24485),
            .I(N__24482));
    InMux I__3575 (
            .O(N__24482),
            .I(N__24479));
    LocalMux I__3574 (
            .O(N__24479),
            .I(N__24476));
    Span4Mux_h I__3573 (
            .O(N__24476),
            .I(N__24473));
    Odrv4 I__3572 (
            .O(N__24473),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0 ));
    InMux I__3571 (
            .O(N__24470),
            .I(N__24467));
    LocalMux I__3570 (
            .O(N__24467),
            .I(N__24464));
    Span4Mux_v I__3569 (
            .O(N__24464),
            .I(N__24461));
    Odrv4 I__3568 (
            .O(N__24461),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__3567 (
            .O(N__24458),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ));
    InMux I__3566 (
            .O(N__24455),
            .I(N__24452));
    LocalMux I__3565 (
            .O(N__24452),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0 ));
    CascadeMux I__3564 (
            .O(N__24449),
            .I(N__24446));
    InMux I__3563 (
            .O(N__24446),
            .I(N__24443));
    LocalMux I__3562 (
            .O(N__24443),
            .I(\current_shift_inst.PI_CTRL.integrator_i_17 ));
    CascadeMux I__3561 (
            .O(N__24440),
            .I(N__24437));
    InMux I__3560 (
            .O(N__24437),
            .I(N__24434));
    LocalMux I__3559 (
            .O(N__24434),
            .I(N__24431));
    Span4Mux_h I__3558 (
            .O(N__24431),
            .I(N__24428));
    Span4Mux_h I__3557 (
            .O(N__24428),
            .I(N__24425));
    Odrv4 I__3556 (
            .O(N__24425),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__3555 (
            .O(N__24422),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ));
    InMux I__3554 (
            .O(N__24419),
            .I(N__24416));
    LocalMux I__3553 (
            .O(N__24416),
            .I(N__24413));
    Span4Mux_v I__3552 (
            .O(N__24413),
            .I(N__24410));
    Odrv4 I__3551 (
            .O(N__24410),
            .I(\current_shift_inst.PI_CTRL.integrator_i_18 ));
    CascadeMux I__3550 (
            .O(N__24407),
            .I(N__24404));
    InMux I__3549 (
            .O(N__24404),
            .I(N__24401));
    LocalMux I__3548 (
            .O(N__24401),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0 ));
    InMux I__3547 (
            .O(N__24398),
            .I(N__24395));
    LocalMux I__3546 (
            .O(N__24395),
            .I(N__24392));
    Span4Mux_h I__3545 (
            .O(N__24392),
            .I(N__24389));
    Odrv4 I__3544 (
            .O(N__24389),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__3543 (
            .O(N__24386),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ));
    CascadeMux I__3542 (
            .O(N__24383),
            .I(N__24380));
    InMux I__3541 (
            .O(N__24380),
            .I(N__24377));
    LocalMux I__3540 (
            .O(N__24377),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0 ));
    InMux I__3539 (
            .O(N__24374),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ));
    InMux I__3538 (
            .O(N__24371),
            .I(N__24368));
    LocalMux I__3537 (
            .O(N__24368),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__3536 (
            .O(N__24365),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ));
    InMux I__3535 (
            .O(N__24362),
            .I(N__24359));
    LocalMux I__3534 (
            .O(N__24359),
            .I(N__24356));
    Span4Mux_v I__3533 (
            .O(N__24356),
            .I(N__24353));
    Odrv4 I__3532 (
            .O(N__24353),
            .I(\current_shift_inst.PI_CTRL.integrator_i_5 ));
    InMux I__3531 (
            .O(N__24350),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ));
    InMux I__3530 (
            .O(N__24347),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ));
    InMux I__3529 (
            .O(N__24344),
            .I(N__24341));
    LocalMux I__3528 (
            .O(N__24341),
            .I(N__24338));
    Odrv4 I__3527 (
            .O(N__24338),
            .I(\current_shift_inst.PI_CTRL.integrator_i_7 ));
    CascadeMux I__3526 (
            .O(N__24335),
            .I(N__24332));
    InMux I__3525 (
            .O(N__24332),
            .I(N__24329));
    LocalMux I__3524 (
            .O(N__24329),
            .I(N__24326));
    Span4Mux_h I__3523 (
            .O(N__24326),
            .I(N__24323));
    Odrv4 I__3522 (
            .O(N__24323),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11 ));
    InMux I__3521 (
            .O(N__24320),
            .I(N__24317));
    LocalMux I__3520 (
            .O(N__24317),
            .I(N__24314));
    Odrv4 I__3519 (
            .O(N__24314),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__3518 (
            .O(N__24311),
            .I(bfn_10_14_0_));
    InMux I__3517 (
            .O(N__24308),
            .I(N__24305));
    LocalMux I__3516 (
            .O(N__24305),
            .I(N__24302));
    Odrv4 I__3515 (
            .O(N__24302),
            .I(\current_shift_inst.PI_CTRL.integrator_i_8 ));
    CascadeMux I__3514 (
            .O(N__24299),
            .I(N__24296));
    InMux I__3513 (
            .O(N__24296),
            .I(N__24293));
    LocalMux I__3512 (
            .O(N__24293),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0 ));
    InMux I__3511 (
            .O(N__24290),
            .I(N__24287));
    LocalMux I__3510 (
            .O(N__24287),
            .I(N__24284));
    Odrv4 I__3509 (
            .O(N__24284),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__3508 (
            .O(N__24281),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ));
    InMux I__3507 (
            .O(N__24278),
            .I(N__24275));
    LocalMux I__3506 (
            .O(N__24275),
            .I(N__24272));
    Span4Mux_v I__3505 (
            .O(N__24272),
            .I(N__24269));
    Odrv4 I__3504 (
            .O(N__24269),
            .I(\current_shift_inst.PI_CTRL.integrator_i_9 ));
    CascadeMux I__3503 (
            .O(N__24266),
            .I(N__24263));
    InMux I__3502 (
            .O(N__24263),
            .I(N__24260));
    LocalMux I__3501 (
            .O(N__24260),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0 ));
    CascadeMux I__3500 (
            .O(N__24257),
            .I(N__24254));
    InMux I__3499 (
            .O(N__24254),
            .I(N__24251));
    LocalMux I__3498 (
            .O(N__24251),
            .I(N__24248));
    Odrv4 I__3497 (
            .O(N__24248),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__3496 (
            .O(N__24245),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ));
    CascadeMux I__3495 (
            .O(N__24242),
            .I(N__24239));
    InMux I__3494 (
            .O(N__24239),
            .I(N__24236));
    LocalMux I__3493 (
            .O(N__24236),
            .I(N__24233));
    Odrv4 I__3492 (
            .O(N__24233),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0 ));
    InMux I__3491 (
            .O(N__24230),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ));
    InMux I__3490 (
            .O(N__24227),
            .I(N__24224));
    LocalMux I__3489 (
            .O(N__24224),
            .I(N__24221));
    Odrv12 I__3488 (
            .O(N__24221),
            .I(\current_shift_inst.PI_CTRL.integrator_i_11 ));
    CascadeMux I__3487 (
            .O(N__24218),
            .I(N__24215));
    InMux I__3486 (
            .O(N__24215),
            .I(N__24212));
    LocalMux I__3485 (
            .O(N__24212),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0 ));
    CascadeMux I__3484 (
            .O(N__24209),
            .I(N__24206));
    InMux I__3483 (
            .O(N__24206),
            .I(N__24203));
    LocalMux I__3482 (
            .O(N__24203),
            .I(N__24200));
    Odrv4 I__3481 (
            .O(N__24200),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__3480 (
            .O(N__24197),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ));
    CascadeMux I__3479 (
            .O(N__24194),
            .I(N__24191));
    InMux I__3478 (
            .O(N__24191),
            .I(N__24187));
    InMux I__3477 (
            .O(N__24190),
            .I(N__24184));
    LocalMux I__3476 (
            .O(N__24187),
            .I(N__24181));
    LocalMux I__3475 (
            .O(N__24184),
            .I(N__24176));
    Span4Mux_h I__3474 (
            .O(N__24181),
            .I(N__24173));
    InMux I__3473 (
            .O(N__24180),
            .I(N__24168));
    InMux I__3472 (
            .O(N__24179),
            .I(N__24168));
    Span4Mux_h I__3471 (
            .O(N__24176),
            .I(N__24162));
    Span4Mux_h I__3470 (
            .O(N__24173),
            .I(N__24162));
    LocalMux I__3469 (
            .O(N__24168),
            .I(N__24159));
    InMux I__3468 (
            .O(N__24167),
            .I(N__24156));
    Odrv4 I__3467 (
            .O(N__24162),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__3466 (
            .O(N__24159),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__3465 (
            .O(N__24156),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__3464 (
            .O(N__24149),
            .I(N__24145));
    InMux I__3463 (
            .O(N__24148),
            .I(N__24142));
    LocalMux I__3462 (
            .O(N__24145),
            .I(N__24139));
    LocalMux I__3461 (
            .O(N__24142),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0 ));
    Odrv4 I__3460 (
            .O(N__24139),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0 ));
    CascadeMux I__3459 (
            .O(N__24134),
            .I(N__24131));
    InMux I__3458 (
            .O(N__24131),
            .I(N__24128));
    LocalMux I__3457 (
            .O(N__24128),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4 ));
    CascadeMux I__3456 (
            .O(N__24125),
            .I(N__24121));
    CascadeMux I__3455 (
            .O(N__24124),
            .I(N__24118));
    InMux I__3454 (
            .O(N__24121),
            .I(N__24115));
    InMux I__3453 (
            .O(N__24118),
            .I(N__24112));
    LocalMux I__3452 (
            .O(N__24115),
            .I(N__24108));
    LocalMux I__3451 (
            .O(N__24112),
            .I(N__24105));
    InMux I__3450 (
            .O(N__24111),
            .I(N__24102));
    Span12Mux_s10_h I__3449 (
            .O(N__24108),
            .I(N__24099));
    Span4Mux_v I__3448 (
            .O(N__24105),
            .I(N__24094));
    LocalMux I__3447 (
            .O(N__24102),
            .I(N__24094));
    Odrv12 I__3446 (
            .O(N__24099),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    Odrv4 I__3445 (
            .O(N__24094),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    InMux I__3444 (
            .O(N__24089),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ));
    InMux I__3443 (
            .O(N__24086),
            .I(N__24083));
    LocalMux I__3442 (
            .O(N__24083),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5 ));
    InMux I__3441 (
            .O(N__24080),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ));
    InMux I__3440 (
            .O(N__24077),
            .I(N__24074));
    LocalMux I__3439 (
            .O(N__24074),
            .I(N__24071));
    Span4Mux_h I__3438 (
            .O(N__24071),
            .I(N__24068));
    Span4Mux_h I__3437 (
            .O(N__24068),
            .I(N__24065));
    Odrv4 I__3436 (
            .O(N__24065),
            .I(\current_shift_inst.PI_CTRL.integrator_i_2 ));
    CascadeMux I__3435 (
            .O(N__24062),
            .I(N__24059));
    InMux I__3434 (
            .O(N__24059),
            .I(N__24056));
    LocalMux I__3433 (
            .O(N__24056),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6 ));
    CascadeMux I__3432 (
            .O(N__24053),
            .I(N__24050));
    InMux I__3431 (
            .O(N__24050),
            .I(N__24045));
    InMux I__3430 (
            .O(N__24049),
            .I(N__24042));
    InMux I__3429 (
            .O(N__24048),
            .I(N__24039));
    LocalMux I__3428 (
            .O(N__24045),
            .I(N__24035));
    LocalMux I__3427 (
            .O(N__24042),
            .I(N__24032));
    LocalMux I__3426 (
            .O(N__24039),
            .I(N__24029));
    InMux I__3425 (
            .O(N__24038),
            .I(N__24026));
    Span4Mux_h I__3424 (
            .O(N__24035),
            .I(N__24023));
    Span4Mux_h I__3423 (
            .O(N__24032),
            .I(N__24020));
    Span4Mux_v I__3422 (
            .O(N__24029),
            .I(N__24017));
    LocalMux I__3421 (
            .O(N__24026),
            .I(N__24010));
    Span4Mux_h I__3420 (
            .O(N__24023),
            .I(N__24010));
    Span4Mux_h I__3419 (
            .O(N__24020),
            .I(N__24010));
    Odrv4 I__3418 (
            .O(N__24017),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__3417 (
            .O(N__24010),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__3416 (
            .O(N__24005),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ));
    InMux I__3415 (
            .O(N__24002),
            .I(N__23999));
    LocalMux I__3414 (
            .O(N__23999),
            .I(N__23996));
    Odrv12 I__3413 (
            .O(N__23996),
            .I(\current_shift_inst.PI_CTRL.integrator_i_3 ));
    CascadeMux I__3412 (
            .O(N__23993),
            .I(N__23990));
    InMux I__3411 (
            .O(N__23990),
            .I(N__23987));
    LocalMux I__3410 (
            .O(N__23987),
            .I(N__23984));
    Odrv4 I__3409 (
            .O(N__23984),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7 ));
    CascadeMux I__3408 (
            .O(N__23981),
            .I(N__23977));
    CascadeMux I__3407 (
            .O(N__23980),
            .I(N__23974));
    InMux I__3406 (
            .O(N__23977),
            .I(N__23970));
    InMux I__3405 (
            .O(N__23974),
            .I(N__23966));
    InMux I__3404 (
            .O(N__23973),
            .I(N__23963));
    LocalMux I__3403 (
            .O(N__23970),
            .I(N__23960));
    InMux I__3402 (
            .O(N__23969),
            .I(N__23956));
    LocalMux I__3401 (
            .O(N__23966),
            .I(N__23951));
    LocalMux I__3400 (
            .O(N__23963),
            .I(N__23951));
    Span4Mux_v I__3399 (
            .O(N__23960),
            .I(N__23948));
    InMux I__3398 (
            .O(N__23959),
            .I(N__23945));
    LocalMux I__3397 (
            .O(N__23956),
            .I(N__23938));
    Span4Mux_h I__3396 (
            .O(N__23951),
            .I(N__23938));
    Span4Mux_h I__3395 (
            .O(N__23948),
            .I(N__23938));
    LocalMux I__3394 (
            .O(N__23945),
            .I(N__23935));
    Odrv4 I__3393 (
            .O(N__23938),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__3392 (
            .O(N__23935),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__3391 (
            .O(N__23930),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ));
    InMux I__3390 (
            .O(N__23927),
            .I(N__23924));
    LocalMux I__3389 (
            .O(N__23924),
            .I(\current_shift_inst.PI_CTRL.integrator_i_4 ));
    CascadeMux I__3388 (
            .O(N__23921),
            .I(N__23918));
    InMux I__3387 (
            .O(N__23918),
            .I(N__23915));
    LocalMux I__3386 (
            .O(N__23915),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8 ));
    CascadeMux I__3385 (
            .O(N__23912),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    InMux I__3384 (
            .O(N__23909),
            .I(N__23906));
    LocalMux I__3383 (
            .O(N__23906),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    CascadeMux I__3382 (
            .O(N__23903),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__3381 (
            .O(N__23900),
            .I(N__23897));
    LocalMux I__3380 (
            .O(N__23897),
            .I(N__23894));
    Span4Mux_h I__3379 (
            .O(N__23894),
            .I(N__23891));
    Odrv4 I__3378 (
            .O(N__23891),
            .I(il_max_comp2_D1));
    InMux I__3377 (
            .O(N__23888),
            .I(N__23885));
    LocalMux I__3376 (
            .O(N__23885),
            .I(il_min_comp1_D1));
    InMux I__3375 (
            .O(N__23882),
            .I(N__23879));
    LocalMux I__3374 (
            .O(N__23879),
            .I(N__23875));
    InMux I__3373 (
            .O(N__23878),
            .I(N__23872));
    Span4Mux_h I__3372 (
            .O(N__23875),
            .I(N__23869));
    LocalMux I__3371 (
            .O(N__23872),
            .I(N__23861));
    Span4Mux_h I__3370 (
            .O(N__23869),
            .I(N__23861));
    InMux I__3369 (
            .O(N__23868),
            .I(N__23856));
    InMux I__3368 (
            .O(N__23867),
            .I(N__23856));
    InMux I__3367 (
            .O(N__23866),
            .I(N__23853));
    Odrv4 I__3366 (
            .O(N__23861),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__3365 (
            .O(N__23856),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__3364 (
            .O(N__23853),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__3363 (
            .O(N__23846),
            .I(N__23842));
    InMux I__3362 (
            .O(N__23845),
            .I(N__23839));
    LocalMux I__3361 (
            .O(N__23842),
            .I(\phase_controller_inst1.stoper_hc.N_287 ));
    LocalMux I__3360 (
            .O(N__23839),
            .I(\phase_controller_inst1.stoper_hc.N_287 ));
    CascadeMux I__3359 (
            .O(N__23834),
            .I(N__23830));
    CascadeMux I__3358 (
            .O(N__23833),
            .I(N__23824));
    InMux I__3357 (
            .O(N__23830),
            .I(N__23821));
    InMux I__3356 (
            .O(N__23829),
            .I(N__23818));
    InMux I__3355 (
            .O(N__23828),
            .I(N__23815));
    InMux I__3354 (
            .O(N__23827),
            .I(N__23810));
    InMux I__3353 (
            .O(N__23824),
            .I(N__23807));
    LocalMux I__3352 (
            .O(N__23821),
            .I(N__23804));
    LocalMux I__3351 (
            .O(N__23818),
            .I(N__23801));
    LocalMux I__3350 (
            .O(N__23815),
            .I(N__23798));
    InMux I__3349 (
            .O(N__23814),
            .I(N__23795));
    InMux I__3348 (
            .O(N__23813),
            .I(N__23792));
    LocalMux I__3347 (
            .O(N__23810),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14));
    LocalMux I__3346 (
            .O(N__23807),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14));
    Odrv4 I__3345 (
            .O(N__23804),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14));
    Odrv4 I__3344 (
            .O(N__23801),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14));
    Odrv4 I__3343 (
            .O(N__23798),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14));
    LocalMux I__3342 (
            .O(N__23795),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14));
    LocalMux I__3341 (
            .O(N__23792),
            .I(elapsed_time_ns_1_RNI1TBED1_0_14));
    InMux I__3340 (
            .O(N__23777),
            .I(N__23773));
    InMux I__3339 (
            .O(N__23776),
            .I(N__23770));
    LocalMux I__3338 (
            .O(N__23773),
            .I(N__23764));
    LocalMux I__3337 (
            .O(N__23770),
            .I(N__23764));
    InMux I__3336 (
            .O(N__23769),
            .I(N__23759));
    Span4Mux_v I__3335 (
            .O(N__23764),
            .I(N__23756));
    InMux I__3334 (
            .O(N__23763),
            .I(N__23751));
    InMux I__3333 (
            .O(N__23762),
            .I(N__23751));
    LocalMux I__3332 (
            .O(N__23759),
            .I(elapsed_time_ns_1_RNI51CED1_0_18));
    Odrv4 I__3331 (
            .O(N__23756),
            .I(elapsed_time_ns_1_RNI51CED1_0_18));
    LocalMux I__3330 (
            .O(N__23751),
            .I(elapsed_time_ns_1_RNI51CED1_0_18));
    InMux I__3329 (
            .O(N__23744),
            .I(N__23739));
    InMux I__3328 (
            .O(N__23743),
            .I(N__23736));
    InMux I__3327 (
            .O(N__23742),
            .I(N__23733));
    LocalMux I__3326 (
            .O(N__23739),
            .I(N__23727));
    LocalMux I__3325 (
            .O(N__23736),
            .I(N__23727));
    LocalMux I__3324 (
            .O(N__23733),
            .I(N__23724));
    InMux I__3323 (
            .O(N__23732),
            .I(N__23721));
    Odrv4 I__3322 (
            .O(N__23727),
            .I(elapsed_time_ns_1_RNI40CED1_0_17));
    Odrv4 I__3321 (
            .O(N__23724),
            .I(elapsed_time_ns_1_RNI40CED1_0_17));
    LocalMux I__3320 (
            .O(N__23721),
            .I(elapsed_time_ns_1_RNI40CED1_0_17));
    CascadeMux I__3319 (
            .O(N__23714),
            .I(N__23709));
    InMux I__3318 (
            .O(N__23713),
            .I(N__23704));
    InMux I__3317 (
            .O(N__23712),
            .I(N__23701));
    InMux I__3316 (
            .O(N__23709),
            .I(N__23696));
    InMux I__3315 (
            .O(N__23708),
            .I(N__23696));
    InMux I__3314 (
            .O(N__23707),
            .I(N__23693));
    LocalMux I__3313 (
            .O(N__23704),
            .I(N__23690));
    LocalMux I__3312 (
            .O(N__23701),
            .I(N__23685));
    LocalMux I__3311 (
            .O(N__23696),
            .I(N__23685));
    LocalMux I__3310 (
            .O(N__23693),
            .I(elapsed_time_ns_1_RNI62CED1_0_19));
    Odrv4 I__3309 (
            .O(N__23690),
            .I(elapsed_time_ns_1_RNI62CED1_0_19));
    Odrv4 I__3308 (
            .O(N__23685),
            .I(elapsed_time_ns_1_RNI62CED1_0_19));
    InMux I__3307 (
            .O(N__23678),
            .I(N__23674));
    InMux I__3306 (
            .O(N__23677),
            .I(N__23671));
    LocalMux I__3305 (
            .O(N__23674),
            .I(N__23666));
    LocalMux I__3304 (
            .O(N__23671),
            .I(N__23666));
    Span4Mux_v I__3303 (
            .O(N__23666),
            .I(N__23661));
    InMux I__3302 (
            .O(N__23665),
            .I(N__23658));
    InMux I__3301 (
            .O(N__23664),
            .I(N__23655));
    Span4Mux_h I__3300 (
            .O(N__23661),
            .I(N__23652));
    LocalMux I__3299 (
            .O(N__23658),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    LocalMux I__3298 (
            .O(N__23655),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__3297 (
            .O(N__23652),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__3296 (
            .O(N__23645),
            .I(N__23641));
    InMux I__3295 (
            .O(N__23644),
            .I(N__23637));
    LocalMux I__3294 (
            .O(N__23641),
            .I(N__23634));
    InMux I__3293 (
            .O(N__23640),
            .I(N__23631));
    LocalMux I__3292 (
            .O(N__23637),
            .I(N__23624));
    Span4Mux_h I__3291 (
            .O(N__23634),
            .I(N__23624));
    LocalMux I__3290 (
            .O(N__23631),
            .I(N__23624));
    Span4Mux_h I__3289 (
            .O(N__23624),
            .I(N__23621));
    Span4Mux_v I__3288 (
            .O(N__23621),
            .I(N__23618));
    Odrv4 I__3287 (
            .O(N__23618),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    IoInMux I__3286 (
            .O(N__23615),
            .I(N__23612));
    LocalMux I__3285 (
            .O(N__23612),
            .I(N__23609));
    Odrv4 I__3284 (
            .O(N__23609),
            .I(s3_phy_c));
    CascadeMux I__3283 (
            .O(N__23606),
            .I(N__23602));
    InMux I__3282 (
            .O(N__23605),
            .I(N__23596));
    InMux I__3281 (
            .O(N__23602),
            .I(N__23593));
    InMux I__3280 (
            .O(N__23601),
            .I(N__23590));
    InMux I__3279 (
            .O(N__23600),
            .I(N__23585));
    InMux I__3278 (
            .O(N__23599),
            .I(N__23585));
    LocalMux I__3277 (
            .O(N__23596),
            .I(elapsed_time_ns_1_RNIL13KD1_0_9));
    LocalMux I__3276 (
            .O(N__23593),
            .I(elapsed_time_ns_1_RNIL13KD1_0_9));
    LocalMux I__3275 (
            .O(N__23590),
            .I(elapsed_time_ns_1_RNIL13KD1_0_9));
    LocalMux I__3274 (
            .O(N__23585),
            .I(elapsed_time_ns_1_RNIL13KD1_0_9));
    InMux I__3273 (
            .O(N__23576),
            .I(N__23573));
    LocalMux I__3272 (
            .O(N__23573),
            .I(N__23569));
    InMux I__3271 (
            .O(N__23572),
            .I(N__23566));
    Span4Mux_v I__3270 (
            .O(N__23569),
            .I(N__23563));
    LocalMux I__3269 (
            .O(N__23566),
            .I(N__23560));
    Odrv4 I__3268 (
            .O(N__23563),
            .I(\phase_controller_inst1.stoper_hc.N_266_iZ0Z_1 ));
    Odrv4 I__3267 (
            .O(N__23560),
            .I(\phase_controller_inst1.stoper_hc.N_266_iZ0Z_1 ));
    InMux I__3266 (
            .O(N__23555),
            .I(N__23551));
    InMux I__3265 (
            .O(N__23554),
            .I(N__23546));
    LocalMux I__3264 (
            .O(N__23551),
            .I(N__23543));
    InMux I__3263 (
            .O(N__23550),
            .I(N__23538));
    InMux I__3262 (
            .O(N__23549),
            .I(N__23538));
    LocalMux I__3261 (
            .O(N__23546),
            .I(elapsed_time_ns_1_RNI3VBED1_0_16));
    Odrv4 I__3260 (
            .O(N__23543),
            .I(elapsed_time_ns_1_RNI3VBED1_0_16));
    LocalMux I__3259 (
            .O(N__23538),
            .I(elapsed_time_ns_1_RNI3VBED1_0_16));
    CascadeMux I__3258 (
            .O(N__23531),
            .I(\phase_controller_inst1.stoper_hc.N_325_cascade_ ));
    CascadeMux I__3257 (
            .O(N__23528),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1_cascade_ ));
    CascadeMux I__3256 (
            .O(N__23525),
            .I(elapsed_time_ns_1_RNIB4DJ11_0_5_cascade_));
    CascadeMux I__3255 (
            .O(N__23522),
            .I(N__23518));
    InMux I__3254 (
            .O(N__23521),
            .I(N__23515));
    InMux I__3253 (
            .O(N__23518),
            .I(N__23512));
    LocalMux I__3252 (
            .O(N__23515),
            .I(N__23508));
    LocalMux I__3251 (
            .O(N__23512),
            .I(N__23505));
    InMux I__3250 (
            .O(N__23511),
            .I(N__23502));
    Span4Mux_h I__3249 (
            .O(N__23508),
            .I(N__23495));
    Span4Mux_h I__3248 (
            .O(N__23505),
            .I(N__23495));
    LocalMux I__3247 (
            .O(N__23502),
            .I(N__23492));
    InMux I__3246 (
            .O(N__23501),
            .I(N__23487));
    InMux I__3245 (
            .O(N__23500),
            .I(N__23487));
    Odrv4 I__3244 (
            .O(N__23495),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__3243 (
            .O(N__23492),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__3242 (
            .O(N__23487),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__3241 (
            .O(N__23480),
            .I(N__23476));
    InMux I__3240 (
            .O(N__23479),
            .I(N__23472));
    LocalMux I__3239 (
            .O(N__23476),
            .I(N__23469));
    InMux I__3238 (
            .O(N__23475),
            .I(N__23466));
    LocalMux I__3237 (
            .O(N__23472),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    Odrv4 I__3236 (
            .O(N__23469),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    LocalMux I__3235 (
            .O(N__23466),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    InMux I__3234 (
            .O(N__23459),
            .I(N__23456));
    LocalMux I__3233 (
            .O(N__23456),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ));
    InMux I__3232 (
            .O(N__23453),
            .I(N__23449));
    InMux I__3231 (
            .O(N__23452),
            .I(N__23446));
    LocalMux I__3230 (
            .O(N__23449),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    LocalMux I__3229 (
            .O(N__23446),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    InMux I__3228 (
            .O(N__23441),
            .I(N__23438));
    LocalMux I__3227 (
            .O(N__23438),
            .I(N__23435));
    Odrv4 I__3226 (
            .O(N__23435),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ));
    CascadeMux I__3225 (
            .O(N__23432),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29_cascade_ ));
    InMux I__3224 (
            .O(N__23429),
            .I(N__23424));
    InMux I__3223 (
            .O(N__23428),
            .I(N__23421));
    InMux I__3222 (
            .O(N__23427),
            .I(N__23418));
    LocalMux I__3221 (
            .O(N__23424),
            .I(N__23413));
    LocalMux I__3220 (
            .O(N__23421),
            .I(N__23410));
    LocalMux I__3219 (
            .O(N__23418),
            .I(N__23407));
    InMux I__3218 (
            .O(N__23417),
            .I(N__23402));
    InMux I__3217 (
            .O(N__23416),
            .I(N__23402));
    Span4Mux_h I__3216 (
            .O(N__23413),
            .I(N__23397));
    Span4Mux_h I__3215 (
            .O(N__23410),
            .I(N__23397));
    Span4Mux_h I__3214 (
            .O(N__23407),
            .I(N__23392));
    LocalMux I__3213 (
            .O(N__23402),
            .I(N__23392));
    Odrv4 I__3212 (
            .O(N__23397),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__3211 (
            .O(N__23392),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__3210 (
            .O(N__23387),
            .I(N__23383));
    InMux I__3209 (
            .O(N__23386),
            .I(N__23380));
    LocalMux I__3208 (
            .O(N__23383),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    LocalMux I__3207 (
            .O(N__23380),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    InMux I__3206 (
            .O(N__23375),
            .I(N__23371));
    CascadeMux I__3205 (
            .O(N__23374),
            .I(N__23368));
    LocalMux I__3204 (
            .O(N__23371),
            .I(N__23365));
    InMux I__3203 (
            .O(N__23368),
            .I(N__23362));
    Span4Mux_v I__3202 (
            .O(N__23365),
            .I(N__23357));
    LocalMux I__3201 (
            .O(N__23362),
            .I(N__23354));
    InMux I__3200 (
            .O(N__23361),
            .I(N__23351));
    InMux I__3199 (
            .O(N__23360),
            .I(N__23348));
    Span4Mux_h I__3198 (
            .O(N__23357),
            .I(N__23342));
    Span4Mux_v I__3197 (
            .O(N__23354),
            .I(N__23342));
    LocalMux I__3196 (
            .O(N__23351),
            .I(N__23339));
    LocalMux I__3195 (
            .O(N__23348),
            .I(N__23336));
    InMux I__3194 (
            .O(N__23347),
            .I(N__23333));
    Odrv4 I__3193 (
            .O(N__23342),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__3192 (
            .O(N__23339),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__3191 (
            .O(N__23336),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__3190 (
            .O(N__23333),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    CascadeMux I__3189 (
            .O(N__23324),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_ ));
    InMux I__3188 (
            .O(N__23321),
            .I(N__23318));
    LocalMux I__3187 (
            .O(N__23318),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ));
    InMux I__3186 (
            .O(N__23315),
            .I(N__23311));
    InMux I__3185 (
            .O(N__23314),
            .I(N__23307));
    LocalMux I__3184 (
            .O(N__23311),
            .I(N__23304));
    InMux I__3183 (
            .O(N__23310),
            .I(N__23301));
    LocalMux I__3182 (
            .O(N__23307),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    Odrv12 I__3181 (
            .O(N__23304),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    LocalMux I__3180 (
            .O(N__23301),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    CascadeMux I__3179 (
            .O(N__23294),
            .I(N__23291));
    InMux I__3178 (
            .O(N__23291),
            .I(N__23286));
    InMux I__3177 (
            .O(N__23290),
            .I(N__23283));
    CascadeMux I__3176 (
            .O(N__23289),
            .I(N__23280));
    LocalMux I__3175 (
            .O(N__23286),
            .I(N__23276));
    LocalMux I__3174 (
            .O(N__23283),
            .I(N__23273));
    InMux I__3173 (
            .O(N__23280),
            .I(N__23270));
    InMux I__3172 (
            .O(N__23279),
            .I(N__23267));
    Span4Mux_h I__3171 (
            .O(N__23276),
            .I(N__23263));
    Span4Mux_v I__3170 (
            .O(N__23273),
            .I(N__23256));
    LocalMux I__3169 (
            .O(N__23270),
            .I(N__23256));
    LocalMux I__3168 (
            .O(N__23267),
            .I(N__23256));
    InMux I__3167 (
            .O(N__23266),
            .I(N__23253));
    Odrv4 I__3166 (
            .O(N__23263),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__3165 (
            .O(N__23256),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__3164 (
            .O(N__23253),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    CascadeMux I__3163 (
            .O(N__23246),
            .I(N__23243));
    InMux I__3162 (
            .O(N__23243),
            .I(N__23240));
    LocalMux I__3161 (
            .O(N__23240),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ));
    CascadeMux I__3160 (
            .O(N__23237),
            .I(\phase_controller_inst1.stoper_hc.N_275_cascade_ ));
    InMux I__3159 (
            .O(N__23234),
            .I(N__23230));
    InMux I__3158 (
            .O(N__23233),
            .I(N__23227));
    LocalMux I__3157 (
            .O(N__23230),
            .I(N__23224));
    LocalMux I__3156 (
            .O(N__23227),
            .I(N__23218));
    Span4Mux_h I__3155 (
            .O(N__23224),
            .I(N__23215));
    InMux I__3154 (
            .O(N__23223),
            .I(N__23212));
    InMux I__3153 (
            .O(N__23222),
            .I(N__23209));
    InMux I__3152 (
            .O(N__23221),
            .I(N__23206));
    Odrv4 I__3151 (
            .O(N__23218),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__3150 (
            .O(N__23215),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__3149 (
            .O(N__23212),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__3148 (
            .O(N__23209),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__3147 (
            .O(N__23206),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__3146 (
            .O(N__23195),
            .I(N__23191));
    InMux I__3145 (
            .O(N__23194),
            .I(N__23188));
    LocalMux I__3144 (
            .O(N__23191),
            .I(N__23182));
    LocalMux I__3143 (
            .O(N__23188),
            .I(N__23182));
    InMux I__3142 (
            .O(N__23187),
            .I(N__23179));
    Sp12to4 I__3141 (
            .O(N__23182),
            .I(N__23176));
    LocalMux I__3140 (
            .O(N__23179),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    Odrv12 I__3139 (
            .O(N__23176),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    InMux I__3138 (
            .O(N__23171),
            .I(N__23168));
    LocalMux I__3137 (
            .O(N__23168),
            .I(N__23165));
    Odrv4 I__3136 (
            .O(N__23165),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ));
    InMux I__3135 (
            .O(N__23162),
            .I(N__23159));
    LocalMux I__3134 (
            .O(N__23159),
            .I(N__23156));
    Span4Mux_v I__3133 (
            .O(N__23156),
            .I(N__23153));
    Odrv4 I__3132 (
            .O(N__23153),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__3131 (
            .O(N__23150),
            .I(N__23147));
    LocalMux I__3130 (
            .O(N__23147),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ));
    InMux I__3129 (
            .O(N__23144),
            .I(N__23140));
    InMux I__3128 (
            .O(N__23143),
            .I(N__23135));
    LocalMux I__3127 (
            .O(N__23140),
            .I(N__23132));
    CascadeMux I__3126 (
            .O(N__23139),
            .I(N__23129));
    InMux I__3125 (
            .O(N__23138),
            .I(N__23125));
    LocalMux I__3124 (
            .O(N__23135),
            .I(N__23122));
    Span4Mux_h I__3123 (
            .O(N__23132),
            .I(N__23119));
    InMux I__3122 (
            .O(N__23129),
            .I(N__23116));
    InMux I__3121 (
            .O(N__23128),
            .I(N__23113));
    LocalMux I__3120 (
            .O(N__23125),
            .I(N__23110));
    Odrv4 I__3119 (
            .O(N__23122),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__3118 (
            .O(N__23119),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__3117 (
            .O(N__23116),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__3116 (
            .O(N__23113),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__3115 (
            .O(N__23110),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    CascadeMux I__3114 (
            .O(N__23099),
            .I(N__23096));
    InMux I__3113 (
            .O(N__23096),
            .I(N__23093));
    LocalMux I__3112 (
            .O(N__23093),
            .I(N__23089));
    InMux I__3111 (
            .O(N__23092),
            .I(N__23085));
    Span4Mux_h I__3110 (
            .O(N__23089),
            .I(N__23082));
    InMux I__3109 (
            .O(N__23088),
            .I(N__23079));
    LocalMux I__3108 (
            .O(N__23085),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    Odrv4 I__3107 (
            .O(N__23082),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    LocalMux I__3106 (
            .O(N__23079),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    InMux I__3105 (
            .O(N__23072),
            .I(N__23069));
    LocalMux I__3104 (
            .O(N__23069),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ));
    CascadeMux I__3103 (
            .O(N__23066),
            .I(N__23062));
    InMux I__3102 (
            .O(N__23065),
            .I(N__23058));
    InMux I__3101 (
            .O(N__23062),
            .I(N__23055));
    InMux I__3100 (
            .O(N__23061),
            .I(N__23052));
    LocalMux I__3099 (
            .O(N__23058),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    LocalMux I__3098 (
            .O(N__23055),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    LocalMux I__3097 (
            .O(N__23052),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    InMux I__3096 (
            .O(N__23045),
            .I(N__23042));
    LocalMux I__3095 (
            .O(N__23042),
            .I(N__23039));
    Odrv4 I__3094 (
            .O(N__23039),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ));
    InMux I__3093 (
            .O(N__23036),
            .I(N__23033));
    LocalMux I__3092 (
            .O(N__23033),
            .I(N__23028));
    InMux I__3091 (
            .O(N__23032),
            .I(N__23025));
    InMux I__3090 (
            .O(N__23031),
            .I(N__23022));
    Span4Mux_h I__3089 (
            .O(N__23028),
            .I(N__23017));
    LocalMux I__3088 (
            .O(N__23025),
            .I(N__23017));
    LocalMux I__3087 (
            .O(N__23022),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    Odrv4 I__3086 (
            .O(N__23017),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    InMux I__3085 (
            .O(N__23012),
            .I(N__23007));
    InMux I__3084 (
            .O(N__23011),
            .I(N__23004));
    InMux I__3083 (
            .O(N__23010),
            .I(N__23001));
    LocalMux I__3082 (
            .O(N__23007),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    LocalMux I__3081 (
            .O(N__23004),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    LocalMux I__3080 (
            .O(N__23001),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    CascadeMux I__3079 (
            .O(N__22994),
            .I(N__22991));
    InMux I__3078 (
            .O(N__22991),
            .I(N__22986));
    InMux I__3077 (
            .O(N__22990),
            .I(N__22982));
    InMux I__3076 (
            .O(N__22989),
            .I(N__22979));
    LocalMux I__3075 (
            .O(N__22986),
            .I(N__22976));
    CascadeMux I__3074 (
            .O(N__22985),
            .I(N__22972));
    LocalMux I__3073 (
            .O(N__22982),
            .I(N__22969));
    LocalMux I__3072 (
            .O(N__22979),
            .I(N__22966));
    Span4Mux_h I__3071 (
            .O(N__22976),
            .I(N__22963));
    InMux I__3070 (
            .O(N__22975),
            .I(N__22960));
    InMux I__3069 (
            .O(N__22972),
            .I(N__22957));
    Span4Mux_v I__3068 (
            .O(N__22969),
            .I(N__22954));
    Odrv4 I__3067 (
            .O(N__22966),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__3066 (
            .O(N__22963),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__3065 (
            .O(N__22960),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__3064 (
            .O(N__22957),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__3063 (
            .O(N__22954),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__3062 (
            .O(N__22943),
            .I(N__22940));
    LocalMux I__3061 (
            .O(N__22940),
            .I(N__22936));
    InMux I__3060 (
            .O(N__22939),
            .I(N__22932));
    Span4Mux_v I__3059 (
            .O(N__22936),
            .I(N__22929));
    InMux I__3058 (
            .O(N__22935),
            .I(N__22926));
    LocalMux I__3057 (
            .O(N__22932),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    Odrv4 I__3056 (
            .O(N__22929),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    LocalMux I__3055 (
            .O(N__22926),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    CascadeMux I__3054 (
            .O(N__22919),
            .I(N__22916));
    InMux I__3053 (
            .O(N__22916),
            .I(N__22913));
    LocalMux I__3052 (
            .O(N__22913),
            .I(N__22910));
    Odrv4 I__3051 (
            .O(N__22910),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ));
    CascadeMux I__3050 (
            .O(N__22907),
            .I(N__22903));
    InMux I__3049 (
            .O(N__22906),
            .I(N__22900));
    InMux I__3048 (
            .O(N__22903),
            .I(N__22897));
    LocalMux I__3047 (
            .O(N__22900),
            .I(N__22892));
    LocalMux I__3046 (
            .O(N__22897),
            .I(N__22889));
    InMux I__3045 (
            .O(N__22896),
            .I(N__22885));
    InMux I__3044 (
            .O(N__22895),
            .I(N__22882));
    Span4Mux_v I__3043 (
            .O(N__22892),
            .I(N__22879));
    Span4Mux_v I__3042 (
            .O(N__22889),
            .I(N__22876));
    InMux I__3041 (
            .O(N__22888),
            .I(N__22873));
    LocalMux I__3040 (
            .O(N__22885),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__3039 (
            .O(N__22882),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__3038 (
            .O(N__22879),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__3037 (
            .O(N__22876),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__3036 (
            .O(N__22873),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    CascadeMux I__3035 (
            .O(N__22862),
            .I(N__22858));
    InMux I__3034 (
            .O(N__22861),
            .I(N__22855));
    InMux I__3033 (
            .O(N__22858),
            .I(N__22852));
    LocalMux I__3032 (
            .O(N__22855),
            .I(N__22849));
    LocalMux I__3031 (
            .O(N__22852),
            .I(N__22846));
    Span4Mux_v I__3030 (
            .O(N__22849),
            .I(N__22842));
    Span4Mux_h I__3029 (
            .O(N__22846),
            .I(N__22839));
    InMux I__3028 (
            .O(N__22845),
            .I(N__22836));
    Odrv4 I__3027 (
            .O(N__22842),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    Odrv4 I__3026 (
            .O(N__22839),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    LocalMux I__3025 (
            .O(N__22836),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__3024 (
            .O(N__22829),
            .I(N__22826));
    LocalMux I__3023 (
            .O(N__22826),
            .I(N__22823));
    Odrv4 I__3022 (
            .O(N__22823),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_8 ));
    CascadeMux I__3021 (
            .O(N__22820),
            .I(N__22817));
    InMux I__3020 (
            .O(N__22817),
            .I(N__22813));
    InMux I__3019 (
            .O(N__22816),
            .I(N__22809));
    LocalMux I__3018 (
            .O(N__22813),
            .I(N__22806));
    InMux I__3017 (
            .O(N__22812),
            .I(N__22803));
    LocalMux I__3016 (
            .O(N__22809),
            .I(N__22800));
    Span4Mux_v I__3015 (
            .O(N__22806),
            .I(N__22797));
    LocalMux I__3014 (
            .O(N__22803),
            .I(N__22794));
    Odrv12 I__3013 (
            .O(N__22800),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    Odrv4 I__3012 (
            .O(N__22797),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    Odrv4 I__3011 (
            .O(N__22794),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__3010 (
            .O(N__22787),
            .I(N__22784));
    LocalMux I__3009 (
            .O(N__22784),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ));
    InMux I__3008 (
            .O(N__22781),
            .I(N__22778));
    LocalMux I__3007 (
            .O(N__22778),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO ));
    CascadeMux I__3006 (
            .O(N__22775),
            .I(N__22772));
    InMux I__3005 (
            .O(N__22772),
            .I(N__22767));
    InMux I__3004 (
            .O(N__22771),
            .I(N__22764));
    InMux I__3003 (
            .O(N__22770),
            .I(N__22761));
    LocalMux I__3002 (
            .O(N__22767),
            .I(N__22758));
    LocalMux I__3001 (
            .O(N__22764),
            .I(N__22755));
    LocalMux I__3000 (
            .O(N__22761),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    Odrv4 I__2999 (
            .O(N__22758),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    Odrv12 I__2998 (
            .O(N__22755),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    InMux I__2997 (
            .O(N__22748),
            .I(N__22745));
    LocalMux I__2996 (
            .O(N__22745),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ));
    InMux I__2995 (
            .O(N__22742),
            .I(N__22738));
    InMux I__2994 (
            .O(N__22741),
            .I(N__22735));
    LocalMux I__2993 (
            .O(N__22738),
            .I(N__22732));
    LocalMux I__2992 (
            .O(N__22735),
            .I(N__22726));
    Span4Mux_v I__2991 (
            .O(N__22732),
            .I(N__22723));
    InMux I__2990 (
            .O(N__22731),
            .I(N__22720));
    InMux I__2989 (
            .O(N__22730),
            .I(N__22715));
    InMux I__2988 (
            .O(N__22729),
            .I(N__22715));
    Odrv4 I__2987 (
            .O(N__22726),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__2986 (
            .O(N__22723),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__2985 (
            .O(N__22720),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__2984 (
            .O(N__22715),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    InMux I__2983 (
            .O(N__22706),
            .I(N__22702));
    InMux I__2982 (
            .O(N__22705),
            .I(N__22699));
    LocalMux I__2981 (
            .O(N__22702),
            .I(N__22696));
    LocalMux I__2980 (
            .O(N__22699),
            .I(N__22690));
    Span4Mux_v I__2979 (
            .O(N__22696),
            .I(N__22690));
    InMux I__2978 (
            .O(N__22695),
            .I(N__22687));
    Odrv4 I__2977 (
            .O(N__22690),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    LocalMux I__2976 (
            .O(N__22687),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    InMux I__2975 (
            .O(N__22682),
            .I(N__22679));
    LocalMux I__2974 (
            .O(N__22679),
            .I(N__22676));
    Odrv4 I__2973 (
            .O(N__22676),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ));
    InMux I__2972 (
            .O(N__22673),
            .I(N__22669));
    InMux I__2971 (
            .O(N__22672),
            .I(N__22666));
    LocalMux I__2970 (
            .O(N__22669),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    LocalMux I__2969 (
            .O(N__22666),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    CascadeMux I__2968 (
            .O(N__22661),
            .I(N__22657));
    InMux I__2967 (
            .O(N__22660),
            .I(N__22654));
    InMux I__2966 (
            .O(N__22657),
            .I(N__22651));
    LocalMux I__2965 (
            .O(N__22654),
            .I(N__22645));
    LocalMux I__2964 (
            .O(N__22651),
            .I(N__22642));
    InMux I__2963 (
            .O(N__22650),
            .I(N__22639));
    InMux I__2962 (
            .O(N__22649),
            .I(N__22633));
    InMux I__2961 (
            .O(N__22648),
            .I(N__22633));
    Span4Mux_h I__2960 (
            .O(N__22645),
            .I(N__22626));
    Span4Mux_h I__2959 (
            .O(N__22642),
            .I(N__22626));
    LocalMux I__2958 (
            .O(N__22639),
            .I(N__22626));
    InMux I__2957 (
            .O(N__22638),
            .I(N__22623));
    LocalMux I__2956 (
            .O(N__22633),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__2955 (
            .O(N__22626),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__2954 (
            .O(N__22623),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    CascadeMux I__2953 (
            .O(N__22616),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_ ));
    InMux I__2952 (
            .O(N__22613),
            .I(N__22610));
    LocalMux I__2951 (
            .O(N__22610),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ));
    CascadeMux I__2950 (
            .O(N__22607),
            .I(N__22604));
    InMux I__2949 (
            .O(N__22604),
            .I(N__22601));
    LocalMux I__2948 (
            .O(N__22601),
            .I(N__22598));
    Odrv12 I__2947 (
            .O(N__22598),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_7 ));
    InMux I__2946 (
            .O(N__22595),
            .I(N__22592));
    LocalMux I__2945 (
            .O(N__22592),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO ));
    InMux I__2944 (
            .O(N__22589),
            .I(N__22586));
    LocalMux I__2943 (
            .O(N__22586),
            .I(N__22583));
    Span4Mux_h I__2942 (
            .O(N__22583),
            .I(N__22580));
    Odrv4 I__2941 (
            .O(N__22580),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ));
    InMux I__2940 (
            .O(N__22577),
            .I(N__22574));
    LocalMux I__2939 (
            .O(N__22574),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_4 ));
    InMux I__2938 (
            .O(N__22571),
            .I(N__22568));
    LocalMux I__2937 (
            .O(N__22568),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_5 ));
    InMux I__2936 (
            .O(N__22565),
            .I(N__22562));
    LocalMux I__2935 (
            .O(N__22562),
            .I(N__22559));
    Span4Mux_v I__2934 (
            .O(N__22559),
            .I(N__22555));
    InMux I__2933 (
            .O(N__22558),
            .I(N__22551));
    Span4Mux_h I__2932 (
            .O(N__22555),
            .I(N__22548));
    InMux I__2931 (
            .O(N__22554),
            .I(N__22545));
    LocalMux I__2930 (
            .O(N__22551),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    Odrv4 I__2929 (
            .O(N__22548),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    LocalMux I__2928 (
            .O(N__22545),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    InMux I__2927 (
            .O(N__22538),
            .I(N__22535));
    LocalMux I__2926 (
            .O(N__22535),
            .I(N__22532));
    Odrv4 I__2925 (
            .O(N__22532),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ));
    InMux I__2924 (
            .O(N__22529),
            .I(N__22526));
    LocalMux I__2923 (
            .O(N__22526),
            .I(N__22522));
    InMux I__2922 (
            .O(N__22525),
            .I(N__22518));
    Span4Mux_h I__2921 (
            .O(N__22522),
            .I(N__22515));
    InMux I__2920 (
            .O(N__22521),
            .I(N__22512));
    LocalMux I__2919 (
            .O(N__22518),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    Odrv4 I__2918 (
            .O(N__22515),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    LocalMux I__2917 (
            .O(N__22512),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    CascadeMux I__2916 (
            .O(N__22505),
            .I(N__22502));
    InMux I__2915 (
            .O(N__22502),
            .I(N__22499));
    LocalMux I__2914 (
            .O(N__22499),
            .I(N__22493));
    CascadeMux I__2913 (
            .O(N__22498),
            .I(N__22490));
    CascadeMux I__2912 (
            .O(N__22497),
            .I(N__22487));
    InMux I__2911 (
            .O(N__22496),
            .I(N__22483));
    Span4Mux_v I__2910 (
            .O(N__22493),
            .I(N__22480));
    InMux I__2909 (
            .O(N__22490),
            .I(N__22475));
    InMux I__2908 (
            .O(N__22487),
            .I(N__22475));
    InMux I__2907 (
            .O(N__22486),
            .I(N__22472));
    LocalMux I__2906 (
            .O(N__22483),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__2905 (
            .O(N__22480),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__2904 (
            .O(N__22475),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__2903 (
            .O(N__22472),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    InMux I__2902 (
            .O(N__22463),
            .I(N__22460));
    LocalMux I__2901 (
            .O(N__22460),
            .I(N__22457));
    Odrv4 I__2900 (
            .O(N__22457),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ));
    InMux I__2899 (
            .O(N__22454),
            .I(N__22451));
    LocalMux I__2898 (
            .O(N__22451),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_6 ));
    CascadeMux I__2897 (
            .O(N__22448),
            .I(N__22445));
    InMux I__2896 (
            .O(N__22445),
            .I(N__22441));
    InMux I__2895 (
            .O(N__22444),
            .I(N__22437));
    LocalMux I__2894 (
            .O(N__22441),
            .I(N__22434));
    InMux I__2893 (
            .O(N__22440),
            .I(N__22431));
    LocalMux I__2892 (
            .O(N__22437),
            .I(N__22428));
    Span4Mux_h I__2891 (
            .O(N__22434),
            .I(N__22425));
    LocalMux I__2890 (
            .O(N__22431),
            .I(N__22422));
    Odrv12 I__2889 (
            .O(N__22428),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv4 I__2888 (
            .O(N__22425),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv4 I__2887 (
            .O(N__22422),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__2886 (
            .O(N__22415),
            .I(N__22412));
    LocalMux I__2885 (
            .O(N__22412),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0 ));
    InMux I__2884 (
            .O(N__22409),
            .I(N__22406));
    LocalMux I__2883 (
            .O(N__22406),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ));
    InMux I__2882 (
            .O(N__22403),
            .I(N__22400));
    LocalMux I__2881 (
            .O(N__22400),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ));
    InMux I__2880 (
            .O(N__22397),
            .I(N__22394));
    LocalMux I__2879 (
            .O(N__22394),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    InMux I__2878 (
            .O(N__22391),
            .I(N__22388));
    LocalMux I__2877 (
            .O(N__22388),
            .I(N__22385));
    Odrv12 I__2876 (
            .O(N__22385),
            .I(\pwm_generator_inst.thresholdZ0Z_8 ));
    CascadeMux I__2875 (
            .O(N__22382),
            .I(N__22379));
    InMux I__2874 (
            .O(N__22379),
            .I(N__22376));
    LocalMux I__2873 (
            .O(N__22376),
            .I(\pwm_generator_inst.counter_i_8 ));
    InMux I__2872 (
            .O(N__22373),
            .I(N__22370));
    LocalMux I__2871 (
            .O(N__22370),
            .I(N__22367));
    Span4Mux_h I__2870 (
            .O(N__22367),
            .I(N__22364));
    Odrv4 I__2869 (
            .O(N__22364),
            .I(\pwm_generator_inst.thresholdZ0Z_9 ));
    CascadeMux I__2868 (
            .O(N__22361),
            .I(N__22358));
    InMux I__2867 (
            .O(N__22358),
            .I(N__22355));
    LocalMux I__2866 (
            .O(N__22355),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__2865 (
            .O(N__22352),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__2864 (
            .O(N__22349),
            .I(N__22346));
    LocalMux I__2863 (
            .O(N__22346),
            .I(N__22343));
    Span4Mux_s0_v I__2862 (
            .O(N__22343),
            .I(N__22340));
    Span4Mux_v I__2861 (
            .O(N__22340),
            .I(N__22337));
    Sp12to4 I__2860 (
            .O(N__22337),
            .I(N__22334));
    Span12Mux_h I__2859 (
            .O(N__22334),
            .I(N__22331));
    Odrv12 I__2858 (
            .O(N__22331),
            .I(pwm_output_c));
    InMux I__2857 (
            .O(N__22328),
            .I(N__22325));
    LocalMux I__2856 (
            .O(N__22325),
            .I(N__22322));
    Odrv12 I__2855 (
            .O(N__22322),
            .I(il_min_comp1_c));
    CascadeMux I__2854 (
            .O(N__22319),
            .I(N__22315));
    InMux I__2853 (
            .O(N__22318),
            .I(N__22312));
    InMux I__2852 (
            .O(N__22315),
            .I(N__22309));
    LocalMux I__2851 (
            .O(N__22312),
            .I(N__22305));
    LocalMux I__2850 (
            .O(N__22309),
            .I(N__22302));
    InMux I__2849 (
            .O(N__22308),
            .I(N__22299));
    Span4Mux_v I__2848 (
            .O(N__22305),
            .I(N__22294));
    Span4Mux_h I__2847 (
            .O(N__22302),
            .I(N__22289));
    LocalMux I__2846 (
            .O(N__22299),
            .I(N__22289));
    InMux I__2845 (
            .O(N__22298),
            .I(N__22284));
    InMux I__2844 (
            .O(N__22297),
            .I(N__22284));
    Odrv4 I__2843 (
            .O(N__22294),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__2842 (
            .O(N__22289),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__2841 (
            .O(N__22284),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__2840 (
            .O(N__22277),
            .I(N__22274));
    LocalMux I__2839 (
            .O(N__22274),
            .I(N__22271));
    Odrv12 I__2838 (
            .O(N__22271),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ));
    InMux I__2837 (
            .O(N__22268),
            .I(N__22265));
    LocalMux I__2836 (
            .O(N__22265),
            .I(N__22262));
    Odrv12 I__2835 (
            .O(N__22262),
            .I(\pwm_generator_inst.thresholdZ0Z_1 ));
    CascadeMux I__2834 (
            .O(N__22259),
            .I(N__22256));
    InMux I__2833 (
            .O(N__22256),
            .I(N__22253));
    LocalMux I__2832 (
            .O(N__22253),
            .I(\pwm_generator_inst.counter_i_1 ));
    InMux I__2831 (
            .O(N__22250),
            .I(N__22247));
    LocalMux I__2830 (
            .O(N__22247),
            .I(N__22244));
    Odrv12 I__2829 (
            .O(N__22244),
            .I(\pwm_generator_inst.thresholdZ0Z_2 ));
    CascadeMux I__2828 (
            .O(N__22241),
            .I(N__22238));
    InMux I__2827 (
            .O(N__22238),
            .I(N__22235));
    LocalMux I__2826 (
            .O(N__22235),
            .I(\pwm_generator_inst.counter_i_2 ));
    InMux I__2825 (
            .O(N__22232),
            .I(N__22229));
    LocalMux I__2824 (
            .O(N__22229),
            .I(N__22226));
    Span4Mux_h I__2823 (
            .O(N__22226),
            .I(N__22223));
    Span4Mux_h I__2822 (
            .O(N__22223),
            .I(N__22220));
    Odrv4 I__2821 (
            .O(N__22220),
            .I(\pwm_generator_inst.thresholdZ0Z_3 ));
    CascadeMux I__2820 (
            .O(N__22217),
            .I(N__22214));
    InMux I__2819 (
            .O(N__22214),
            .I(N__22211));
    LocalMux I__2818 (
            .O(N__22211),
            .I(\pwm_generator_inst.counter_i_3 ));
    InMux I__2817 (
            .O(N__22208),
            .I(N__22205));
    LocalMux I__2816 (
            .O(N__22205),
            .I(N__22202));
    Span4Mux_h I__2815 (
            .O(N__22202),
            .I(N__22199));
    Odrv4 I__2814 (
            .O(N__22199),
            .I(\pwm_generator_inst.thresholdZ0Z_4 ));
    CascadeMux I__2813 (
            .O(N__22196),
            .I(N__22193));
    InMux I__2812 (
            .O(N__22193),
            .I(N__22190));
    LocalMux I__2811 (
            .O(N__22190),
            .I(\pwm_generator_inst.counter_i_4 ));
    InMux I__2810 (
            .O(N__22187),
            .I(N__22184));
    LocalMux I__2809 (
            .O(N__22184),
            .I(N__22181));
    Odrv12 I__2808 (
            .O(N__22181),
            .I(\pwm_generator_inst.thresholdZ0Z_5 ));
    CascadeMux I__2807 (
            .O(N__22178),
            .I(N__22175));
    InMux I__2806 (
            .O(N__22175),
            .I(N__22172));
    LocalMux I__2805 (
            .O(N__22172),
            .I(\pwm_generator_inst.counter_i_5 ));
    CascadeMux I__2804 (
            .O(N__22169),
            .I(N__22166));
    InMux I__2803 (
            .O(N__22166),
            .I(N__22163));
    LocalMux I__2802 (
            .O(N__22163),
            .I(N__22160));
    Odrv4 I__2801 (
            .O(N__22160),
            .I(\pwm_generator_inst.thresholdZ0Z_6 ));
    InMux I__2800 (
            .O(N__22157),
            .I(N__22154));
    LocalMux I__2799 (
            .O(N__22154),
            .I(\pwm_generator_inst.counter_i_6 ));
    CascadeMux I__2798 (
            .O(N__22151),
            .I(N__22148));
    InMux I__2797 (
            .O(N__22148),
            .I(N__22145));
    LocalMux I__2796 (
            .O(N__22145),
            .I(N__22142));
    Odrv12 I__2795 (
            .O(N__22142),
            .I(\pwm_generator_inst.thresholdZ0Z_7 ));
    InMux I__2794 (
            .O(N__22139),
            .I(N__22136));
    LocalMux I__2793 (
            .O(N__22136),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__2792 (
            .O(N__22133),
            .I(elapsed_time_ns_1_RNI40CED1_0_17_cascade_));
    InMux I__2791 (
            .O(N__22130),
            .I(N__22127));
    LocalMux I__2790 (
            .O(N__22127),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17 ));
    CascadeMux I__2789 (
            .O(N__22124),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3_cascade_ ));
    CascadeMux I__2788 (
            .O(N__22121),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21_cascade_ ));
    InMux I__2787 (
            .O(N__22118),
            .I(N__22115));
    LocalMux I__2786 (
            .O(N__22115),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24 ));
    InMux I__2785 (
            .O(N__22112),
            .I(N__22109));
    LocalMux I__2784 (
            .O(N__22109),
            .I(N__22106));
    Odrv4 I__2783 (
            .O(N__22106),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19 ));
    CascadeMux I__2782 (
            .O(N__22103),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_cascade_ ));
    InMux I__2781 (
            .O(N__22100),
            .I(N__22097));
    LocalMux I__2780 (
            .O(N__22097),
            .I(N__22094));
    Odrv12 I__2779 (
            .O(N__22094),
            .I(\pwm_generator_inst.thresholdZ0Z_0 ));
    CascadeMux I__2778 (
            .O(N__22091),
            .I(N__22088));
    InMux I__2777 (
            .O(N__22088),
            .I(N__22085));
    LocalMux I__2776 (
            .O(N__22085),
            .I(N__22082));
    Odrv4 I__2775 (
            .O(N__22082),
            .I(\pwm_generator_inst.counter_i_0 ));
    InMux I__2774 (
            .O(N__22079),
            .I(N__22076));
    LocalMux I__2773 (
            .O(N__22076),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9 ));
    InMux I__2772 (
            .O(N__22073),
            .I(N__22070));
    LocalMux I__2771 (
            .O(N__22070),
            .I(N__22067));
    Span4Mux_h I__2770 (
            .O(N__22067),
            .I(N__22064));
    Odrv4 I__2769 (
            .O(N__22064),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__2768 (
            .O(N__22061),
            .I(N__22058));
    LocalMux I__2767 (
            .O(N__22058),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14 ));
    CascadeMux I__2766 (
            .O(N__22055),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_ ));
    CascadeMux I__2765 (
            .O(N__22052),
            .I(elapsed_time_ns_1_RNI3VBED1_0_16_cascade_));
    CascadeMux I__2764 (
            .O(N__22049),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_ ));
    InMux I__2763 (
            .O(N__22046),
            .I(N__22043));
    LocalMux I__2762 (
            .O(N__22043),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2 ));
    InMux I__2761 (
            .O(N__22040),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ));
    InMux I__2760 (
            .O(N__22037),
            .I(bfn_8_18_0_));
    InMux I__2759 (
            .O(N__22034),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ));
    InMux I__2758 (
            .O(N__22031),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ));
    InMux I__2757 (
            .O(N__22028),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ));
    InMux I__2756 (
            .O(N__22025),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ));
    InMux I__2755 (
            .O(N__22022),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ));
    InMux I__2754 (
            .O(N__22019),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ));
    InMux I__2753 (
            .O(N__22016),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_31 ));
    InMux I__2752 (
            .O(N__22013),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ));
    InMux I__2751 (
            .O(N__22010),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ));
    InMux I__2750 (
            .O(N__22007),
            .I(bfn_8_17_0_));
    InMux I__2749 (
            .O(N__22004),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ));
    InMux I__2748 (
            .O(N__22001),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ));
    InMux I__2747 (
            .O(N__21998),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ));
    InMux I__2746 (
            .O(N__21995),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ));
    InMux I__2745 (
            .O(N__21992),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ));
    InMux I__2744 (
            .O(N__21989),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ));
    InMux I__2743 (
            .O(N__21986),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ));
    InMux I__2742 (
            .O(N__21983),
            .I(N__21980));
    LocalMux I__2741 (
            .O(N__21980),
            .I(N__21977));
    Odrv4 I__2740 (
            .O(N__21977),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ));
    InMux I__2739 (
            .O(N__21974),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ));
    InMux I__2738 (
            .O(N__21971),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ));
    InMux I__2737 (
            .O(N__21968),
            .I(N__21965));
    LocalMux I__2736 (
            .O(N__21965),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ));
    InMux I__2735 (
            .O(N__21962),
            .I(bfn_8_16_0_));
    InMux I__2734 (
            .O(N__21959),
            .I(N__21956));
    LocalMux I__2733 (
            .O(N__21956),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ));
    InMux I__2732 (
            .O(N__21953),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ));
    InMux I__2731 (
            .O(N__21950),
            .I(N__21947));
    LocalMux I__2730 (
            .O(N__21947),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ));
    InMux I__2729 (
            .O(N__21944),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ));
    InMux I__2728 (
            .O(N__21941),
            .I(N__21938));
    LocalMux I__2727 (
            .O(N__21938),
            .I(N__21935));
    Odrv12 I__2726 (
            .O(N__21935),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ));
    InMux I__2725 (
            .O(N__21932),
            .I(N__21929));
    LocalMux I__2724 (
            .O(N__21929),
            .I(N__21926));
    Odrv4 I__2723 (
            .O(N__21926),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_11 ));
    InMux I__2722 (
            .O(N__21923),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ));
    InMux I__2721 (
            .O(N__21920),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ));
    InMux I__2720 (
            .O(N__21917),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ));
    InMux I__2719 (
            .O(N__21914),
            .I(N__21910));
    InMux I__2718 (
            .O(N__21913),
            .I(N__21907));
    LocalMux I__2717 (
            .O(N__21910),
            .I(N__21904));
    LocalMux I__2716 (
            .O(N__21907),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    Odrv4 I__2715 (
            .O(N__21904),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__2714 (
            .O(N__21899),
            .I(N__21896));
    LocalMux I__2713 (
            .O(N__21896),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ));
    InMux I__2712 (
            .O(N__21893),
            .I(N__21890));
    LocalMux I__2711 (
            .O(N__21890),
            .I(N__21886));
    InMux I__2710 (
            .O(N__21889),
            .I(N__21883));
    Odrv4 I__2709 (
            .O(N__21886),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    LocalMux I__2708 (
            .O(N__21883),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__2707 (
            .O(N__21878),
            .I(N__21875));
    LocalMux I__2706 (
            .O(N__21875),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ));
    InMux I__2705 (
            .O(N__21872),
            .I(N__21869));
    LocalMux I__2704 (
            .O(N__21869),
            .I(N__21865));
    InMux I__2703 (
            .O(N__21868),
            .I(N__21862));
    Odrv12 I__2702 (
            .O(N__21865),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    LocalMux I__2701 (
            .O(N__21862),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__2700 (
            .O(N__21857),
            .I(N__21854));
    LocalMux I__2699 (
            .O(N__21854),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ));
    InMux I__2698 (
            .O(N__21851),
            .I(N__21848));
    LocalMux I__2697 (
            .O(N__21848),
            .I(N__21845));
    Span4Mux_v I__2696 (
            .O(N__21845),
            .I(N__21841));
    InMux I__2695 (
            .O(N__21844),
            .I(N__21838));
    Odrv4 I__2694 (
            .O(N__21841),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    LocalMux I__2693 (
            .O(N__21838),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__2692 (
            .O(N__21833),
            .I(N__21830));
    LocalMux I__2691 (
            .O(N__21830),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ));
    InMux I__2690 (
            .O(N__21827),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ));
    InMux I__2689 (
            .O(N__21824),
            .I(N__21821));
    LocalMux I__2688 (
            .O(N__21821),
            .I(N__21818));
    Odrv4 I__2687 (
            .O(N__21818),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__2686 (
            .O(N__21815),
            .I(N__21810));
    InMux I__2685 (
            .O(N__21814),
            .I(N__21807));
    InMux I__2684 (
            .O(N__21813),
            .I(N__21804));
    LocalMux I__2683 (
            .O(N__21810),
            .I(N__21799));
    LocalMux I__2682 (
            .O(N__21807),
            .I(N__21799));
    LocalMux I__2681 (
            .O(N__21804),
            .I(N__21794));
    Span4Mux_v I__2680 (
            .O(N__21799),
            .I(N__21794));
    Odrv4 I__2679 (
            .O(N__21794),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__2678 (
            .O(N__21791),
            .I(N__21788));
    LocalMux I__2677 (
            .O(N__21788),
            .I(N__21785));
    Odrv4 I__2676 (
            .O(N__21785),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    CascadeMux I__2675 (
            .O(N__21782),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16_cascade_ ));
    InMux I__2674 (
            .O(N__21779),
            .I(N__21776));
    LocalMux I__2673 (
            .O(N__21776),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18 ));
    CascadeMux I__2672 (
            .O(N__21773),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_ ));
    InMux I__2671 (
            .O(N__21770),
            .I(N__21767));
    LocalMux I__2670 (
            .O(N__21767),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    InMux I__2669 (
            .O(N__21764),
            .I(N__21761));
    LocalMux I__2668 (
            .O(N__21761),
            .I(\current_shift_inst.PI_CTRL.N_62 ));
    InMux I__2667 (
            .O(N__21758),
            .I(N__21755));
    LocalMux I__2666 (
            .O(N__21755),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ));
    InMux I__2665 (
            .O(N__21752),
            .I(N__21749));
    LocalMux I__2664 (
            .O(N__21749),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    CascadeMux I__2663 (
            .O(N__21746),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18_cascade_ ));
    IoInMux I__2662 (
            .O(N__21743),
            .I(N__21740));
    LocalMux I__2661 (
            .O(N__21740),
            .I(N__21737));
    IoSpan4Mux I__2660 (
            .O(N__21737),
            .I(N__21734));
    Span4Mux_s2_v I__2659 (
            .O(N__21734),
            .I(N__21731));
    Odrv4 I__2658 (
            .O(N__21731),
            .I(\delay_measurement_inst.delay_hc_timer.N_432_i ));
    InMux I__2657 (
            .O(N__21728),
            .I(N__21725));
    LocalMux I__2656 (
            .O(N__21725),
            .I(N__21722));
    Odrv12 I__2655 (
            .O(N__21722),
            .I(il_max_comp1_c));
    InMux I__2654 (
            .O(N__21719),
            .I(N__21716));
    LocalMux I__2653 (
            .O(N__21716),
            .I(N__21713));
    Span4Mux_h I__2652 (
            .O(N__21713),
            .I(N__21710));
    Span4Mux_v I__2651 (
            .O(N__21710),
            .I(N__21707));
    Odrv4 I__2650 (
            .O(N__21707),
            .I(il_max_comp2_c));
    InMux I__2649 (
            .O(N__21704),
            .I(N__21701));
    LocalMux I__2648 (
            .O(N__21701),
            .I(N__21698));
    Span12Mux_h I__2647 (
            .O(N__21698),
            .I(N__21695));
    Odrv12 I__2646 (
            .O(N__21695),
            .I(il_min_comp2_c));
    InMux I__2645 (
            .O(N__21692),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__2644 (
            .O(N__21689),
            .I(bfn_7_16_0_));
    InMux I__2643 (
            .O(N__21686),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__2642 (
            .O(N__21683),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__2641 (
            .O(N__21680),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__2640 (
            .O(N__21677),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__2639 (
            .O(N__21674),
            .I(N__21671));
    LocalMux I__2638 (
            .O(N__21671),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__2637 (
            .O(N__21668),
            .I(N__21665));
    LocalMux I__2636 (
            .O(N__21665),
            .I(N__21662));
    Odrv12 I__2635 (
            .O(N__21662),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__2634 (
            .O(N__21659),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__2633 (
            .O(N__21656),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__2632 (
            .O(N__21653),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__2631 (
            .O(N__21650),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__2630 (
            .O(N__21647),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__2629 (
            .O(N__21644),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__2628 (
            .O(N__21641),
            .I(N__21638));
    LocalMux I__2627 (
            .O(N__21638),
            .I(\current_shift_inst.PI_CTRL.N_74_16 ));
    InMux I__2626 (
            .O(N__21635),
            .I(N__21629));
    InMux I__2625 (
            .O(N__21634),
            .I(N__21629));
    LocalMux I__2624 (
            .O(N__21629),
            .I(\current_shift_inst.PI_CTRL.N_74_21 ));
    InMux I__2623 (
            .O(N__21626),
            .I(N__21620));
    InMux I__2622 (
            .O(N__21625),
            .I(N__21620));
    LocalMux I__2621 (
            .O(N__21620),
            .I(\current_shift_inst.PI_CTRL.N_72 ));
    CascadeMux I__2620 (
            .O(N__21617),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_1_cascade_ ));
    InMux I__2619 (
            .O(N__21614),
            .I(N__21611));
    LocalMux I__2618 (
            .O(N__21611),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    CascadeMux I__2617 (
            .O(N__21608),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31_cascade_ ));
    InMux I__2616 (
            .O(N__21605),
            .I(N__21602));
    LocalMux I__2615 (
            .O(N__21602),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ));
    CascadeMux I__2614 (
            .O(N__21599),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7_cascade_ ));
    CascadeMux I__2613 (
            .O(N__21596),
            .I(\current_shift_inst.PI_CTRL.N_74_16_cascade_ ));
    InMux I__2612 (
            .O(N__21593),
            .I(N__21590));
    LocalMux I__2611 (
            .O(N__21590),
            .I(N__21587));
    Odrv4 I__2610 (
            .O(N__21587),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    InMux I__2609 (
            .O(N__21584),
            .I(N__21581));
    LocalMux I__2608 (
            .O(N__21581),
            .I(N__21578));
    Odrv4 I__2607 (
            .O(N__21578),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    InMux I__2606 (
            .O(N__21575),
            .I(N__21572));
    LocalMux I__2605 (
            .O(N__21572),
            .I(N__21569));
    Odrv4 I__2604 (
            .O(N__21569),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    InMux I__2603 (
            .O(N__21566),
            .I(N__21563));
    LocalMux I__2602 (
            .O(N__21563),
            .I(N__21560));
    Odrv4 I__2601 (
            .O(N__21560),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    InMux I__2600 (
            .O(N__21557),
            .I(N__21554));
    LocalMux I__2599 (
            .O(N__21554),
            .I(N__21551));
    Odrv4 I__2598 (
            .O(N__21551),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    InMux I__2597 (
            .O(N__21548),
            .I(N__21545));
    LocalMux I__2596 (
            .O(N__21545),
            .I(N__21542));
    Odrv4 I__2595 (
            .O(N__21542),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__2594 (
            .O(N__21539),
            .I(N__21536));
    LocalMux I__2593 (
            .O(N__21536),
            .I(N__21533));
    Span4Mux_h I__2592 (
            .O(N__21533),
            .I(N__21530));
    Odrv4 I__2591 (
            .O(N__21530),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    CascadeMux I__2590 (
            .O(N__21527),
            .I(N__21516));
    CascadeMux I__2589 (
            .O(N__21526),
            .I(N__21512));
    CascadeMux I__2588 (
            .O(N__21525),
            .I(N__21508));
    CascadeMux I__2587 (
            .O(N__21524),
            .I(N__21504));
    CascadeMux I__2586 (
            .O(N__21523),
            .I(N__21500));
    CascadeMux I__2585 (
            .O(N__21522),
            .I(N__21496));
    CascadeMux I__2584 (
            .O(N__21521),
            .I(N__21492));
    InMux I__2583 (
            .O(N__21520),
            .I(N__21472));
    InMux I__2582 (
            .O(N__21519),
            .I(N__21472));
    InMux I__2581 (
            .O(N__21516),
            .I(N__21472));
    InMux I__2580 (
            .O(N__21515),
            .I(N__21472));
    InMux I__2579 (
            .O(N__21512),
            .I(N__21472));
    InMux I__2578 (
            .O(N__21511),
            .I(N__21472));
    InMux I__2577 (
            .O(N__21508),
            .I(N__21472));
    InMux I__2576 (
            .O(N__21507),
            .I(N__21472));
    InMux I__2575 (
            .O(N__21504),
            .I(N__21455));
    InMux I__2574 (
            .O(N__21503),
            .I(N__21455));
    InMux I__2573 (
            .O(N__21500),
            .I(N__21455));
    InMux I__2572 (
            .O(N__21499),
            .I(N__21455));
    InMux I__2571 (
            .O(N__21496),
            .I(N__21455));
    InMux I__2570 (
            .O(N__21495),
            .I(N__21455));
    InMux I__2569 (
            .O(N__21492),
            .I(N__21455));
    InMux I__2568 (
            .O(N__21491),
            .I(N__21455));
    CascadeMux I__2567 (
            .O(N__21490),
            .I(N__21452));
    CascadeMux I__2566 (
            .O(N__21489),
            .I(N__21448));
    LocalMux I__2565 (
            .O(N__21472),
            .I(N__21442));
    LocalMux I__2564 (
            .O(N__21455),
            .I(N__21442));
    InMux I__2563 (
            .O(N__21452),
            .I(N__21433));
    InMux I__2562 (
            .O(N__21451),
            .I(N__21433));
    InMux I__2561 (
            .O(N__21448),
            .I(N__21433));
    InMux I__2560 (
            .O(N__21447),
            .I(N__21433));
    Span4Mux_v I__2559 (
            .O(N__21442),
            .I(N__21428));
    LocalMux I__2558 (
            .O(N__21433),
            .I(N__21428));
    Odrv4 I__2557 (
            .O(N__21428),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__2556 (
            .O(N__21425),
            .I(N__21422));
    LocalMux I__2555 (
            .O(N__21422),
            .I(N__21419));
    Odrv12 I__2554 (
            .O(N__21419),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    InMux I__2553 (
            .O(N__21416),
            .I(N__21413));
    LocalMux I__2552 (
            .O(N__21413),
            .I(N__21410));
    Odrv12 I__2551 (
            .O(N__21410),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__2550 (
            .O(N__21407),
            .I(N__21404));
    LocalMux I__2549 (
            .O(N__21404),
            .I(N__21401));
    Odrv12 I__2548 (
            .O(N__21401),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    CascadeMux I__2547 (
            .O(N__21398),
            .I(N__21395));
    InMux I__2546 (
            .O(N__21395),
            .I(N__21392));
    LocalMux I__2545 (
            .O(N__21392),
            .I(N__21389));
    Odrv12 I__2544 (
            .O(N__21389),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    ClkMux I__2543 (
            .O(N__21386),
            .I(N__21380));
    ClkMux I__2542 (
            .O(N__21385),
            .I(N__21380));
    GlobalMux I__2541 (
            .O(N__21380),
            .I(N__21377));
    gio2CtrlBuf I__2540 (
            .O(N__21377),
            .I(delay_hc_input_c_g));
    InMux I__2539 (
            .O(N__21374),
            .I(N__21371));
    LocalMux I__2538 (
            .O(N__21371),
            .I(N__21368));
    Glb2LocalMux I__2537 (
            .O(N__21368),
            .I(N__21365));
    GlobalMux I__2536 (
            .O(N__21365),
            .I(clk_12mhz));
    IoInMux I__2535 (
            .O(N__21362),
            .I(N__21359));
    LocalMux I__2534 (
            .O(N__21359),
            .I(N__21356));
    IoSpan4Mux I__2533 (
            .O(N__21356),
            .I(N__21353));
    Span4Mux_s0_v I__2532 (
            .O(N__21353),
            .I(N__21350));
    Odrv4 I__2531 (
            .O(N__21350),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__2530 (
            .O(N__21347),
            .I(N__21344));
    LocalMux I__2529 (
            .O(N__21344),
            .I(N__21341));
    Span4Mux_h I__2528 (
            .O(N__21341),
            .I(N__21338));
    Odrv4 I__2527 (
            .O(N__21338),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_6 ));
    InMux I__2526 (
            .O(N__21335),
            .I(N__21332));
    LocalMux I__2525 (
            .O(N__21332),
            .I(N__21329));
    Span4Mux_h I__2524 (
            .O(N__21329),
            .I(N__21326));
    Odrv4 I__2523 (
            .O(N__21326),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_4 ));
    InMux I__2522 (
            .O(N__21323),
            .I(N__21320));
    LocalMux I__2521 (
            .O(N__21320),
            .I(N__21317));
    Odrv12 I__2520 (
            .O(N__21317),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_9 ));
    CascadeMux I__2519 (
            .O(N__21314),
            .I(N__21310));
    InMux I__2518 (
            .O(N__21313),
            .I(N__21307));
    InMux I__2517 (
            .O(N__21310),
            .I(N__21304));
    LocalMux I__2516 (
            .O(N__21307),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    LocalMux I__2515 (
            .O(N__21304),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2514 (
            .O(N__21299),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__2513 (
            .O(N__21296),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__2512 (
            .O(N__21293),
            .I(N__21287));
    InMux I__2511 (
            .O(N__21292),
            .I(N__21287));
    LocalMux I__2510 (
            .O(N__21287),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2509 (
            .O(N__21284),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2508 (
            .O(N__21281),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2507 (
            .O(N__21278),
            .I(N__21274));
    InMux I__2506 (
            .O(N__21277),
            .I(N__21266));
    LocalMux I__2505 (
            .O(N__21274),
            .I(N__21261));
    InMux I__2504 (
            .O(N__21273),
            .I(N__21254));
    InMux I__2503 (
            .O(N__21272),
            .I(N__21254));
    InMux I__2502 (
            .O(N__21271),
            .I(N__21254));
    InMux I__2501 (
            .O(N__21270),
            .I(N__21248));
    InMux I__2500 (
            .O(N__21269),
            .I(N__21248));
    LocalMux I__2499 (
            .O(N__21266),
            .I(N__21245));
    InMux I__2498 (
            .O(N__21265),
            .I(N__21240));
    InMux I__2497 (
            .O(N__21264),
            .I(N__21240));
    Span4Mux_h I__2496 (
            .O(N__21261),
            .I(N__21237));
    LocalMux I__2495 (
            .O(N__21254),
            .I(N__21234));
    InMux I__2494 (
            .O(N__21253),
            .I(N__21231));
    LocalMux I__2493 (
            .O(N__21248),
            .I(N__21226));
    Span4Mux_h I__2492 (
            .O(N__21245),
            .I(N__21226));
    LocalMux I__2491 (
            .O(N__21240),
            .I(N__21223));
    Span4Mux_v I__2490 (
            .O(N__21237),
            .I(N__21216));
    Span4Mux_h I__2489 (
            .O(N__21234),
            .I(N__21216));
    LocalMux I__2488 (
            .O(N__21231),
            .I(N__21216));
    Span4Mux_v I__2487 (
            .O(N__21226),
            .I(N__21213));
    Odrv12 I__2486 (
            .O(N__21223),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2485 (
            .O(N__21216),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2484 (
            .O(N__21213),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__2483 (
            .O(N__21206),
            .I(N__21203));
    LocalMux I__2482 (
            .O(N__21203),
            .I(N__21199));
    InMux I__2481 (
            .O(N__21202),
            .I(N__21196));
    Odrv4 I__2480 (
            .O(N__21199),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    LocalMux I__2479 (
            .O(N__21196),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2478 (
            .O(N__21191),
            .I(N__21188));
    LocalMux I__2477 (
            .O(N__21188),
            .I(N__21184));
    InMux I__2476 (
            .O(N__21187),
            .I(N__21181));
    Odrv4 I__2475 (
            .O(N__21184),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    LocalMux I__2474 (
            .O(N__21181),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    CascadeMux I__2473 (
            .O(N__21176),
            .I(N__21173));
    InMux I__2472 (
            .O(N__21173),
            .I(N__21170));
    LocalMux I__2471 (
            .O(N__21170),
            .I(N__21166));
    InMux I__2470 (
            .O(N__21169),
            .I(N__21163));
    Odrv4 I__2469 (
            .O(N__21166),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    LocalMux I__2468 (
            .O(N__21163),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    CascadeMux I__2467 (
            .O(N__21158),
            .I(N__21154));
    InMux I__2466 (
            .O(N__21157),
            .I(N__21151));
    InMux I__2465 (
            .O(N__21154),
            .I(N__21148));
    LocalMux I__2464 (
            .O(N__21151),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    LocalMux I__2463 (
            .O(N__21148),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2462 (
            .O(N__21143),
            .I(N__21140));
    LocalMux I__2461 (
            .O(N__21140),
            .I(N__21136));
    InMux I__2460 (
            .O(N__21139),
            .I(N__21133));
    Odrv4 I__2459 (
            .O(N__21136),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    LocalMux I__2458 (
            .O(N__21133),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    CascadeMux I__2457 (
            .O(N__21128),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ));
    InMux I__2456 (
            .O(N__21125),
            .I(N__21122));
    LocalMux I__2455 (
            .O(N__21122),
            .I(N__21118));
    InMux I__2454 (
            .O(N__21121),
            .I(N__21115));
    Odrv4 I__2453 (
            .O(N__21118),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    LocalMux I__2452 (
            .O(N__21115),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2451 (
            .O(N__21110),
            .I(N__21107));
    LocalMux I__2450 (
            .O(N__21107),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    CascadeMux I__2449 (
            .O(N__21104),
            .I(N__21101));
    InMux I__2448 (
            .O(N__21101),
            .I(N__21097));
    InMux I__2447 (
            .O(N__21100),
            .I(N__21094));
    LocalMux I__2446 (
            .O(N__21097),
            .I(N__21089));
    LocalMux I__2445 (
            .O(N__21094),
            .I(N__21089));
    Odrv4 I__2444 (
            .O(N__21089),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2443 (
            .O(N__21086),
            .I(N__21083));
    LocalMux I__2442 (
            .O(N__21083),
            .I(N__21079));
    InMux I__2441 (
            .O(N__21082),
            .I(N__21076));
    Odrv4 I__2440 (
            .O(N__21079),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    LocalMux I__2439 (
            .O(N__21076),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2438 (
            .O(N__21071),
            .I(N__21068));
    LocalMux I__2437 (
            .O(N__21068),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    InMux I__2436 (
            .O(N__21065),
            .I(N__21059));
    InMux I__2435 (
            .O(N__21064),
            .I(N__21059));
    LocalMux I__2434 (
            .O(N__21059),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2433 (
            .O(N__21056),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    InMux I__2432 (
            .O(N__21053),
            .I(N__21050));
    LocalMux I__2431 (
            .O(N__21050),
            .I(N__21047));
    Span4Mux_h I__2430 (
            .O(N__21047),
            .I(N__21043));
    InMux I__2429 (
            .O(N__21046),
            .I(N__21040));
    Odrv4 I__2428 (
            .O(N__21043),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    LocalMux I__2427 (
            .O(N__21040),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2426 (
            .O(N__21035),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__2425 (
            .O(N__21032),
            .I(N__21029));
    LocalMux I__2424 (
            .O(N__21029),
            .I(N__21026));
    Span4Mux_h I__2423 (
            .O(N__21026),
            .I(N__21022));
    InMux I__2422 (
            .O(N__21025),
            .I(N__21019));
    Odrv4 I__2421 (
            .O(N__21022),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    LocalMux I__2420 (
            .O(N__21019),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2419 (
            .O(N__21014),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__2418 (
            .O(N__21011),
            .I(N__21005));
    InMux I__2417 (
            .O(N__21010),
            .I(N__21005));
    LocalMux I__2416 (
            .O(N__21005),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2415 (
            .O(N__21002),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__2414 (
            .O(N__20999),
            .I(N__20993));
    InMux I__2413 (
            .O(N__20998),
            .I(N__20993));
    LocalMux I__2412 (
            .O(N__20993),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2411 (
            .O(N__20990),
            .I(bfn_5_13_0_));
    InMux I__2410 (
            .O(N__20987),
            .I(N__20981));
    InMux I__2409 (
            .O(N__20986),
            .I(N__20981));
    LocalMux I__2408 (
            .O(N__20981),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2407 (
            .O(N__20978),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ));
    InMux I__2406 (
            .O(N__20975),
            .I(N__20969));
    InMux I__2405 (
            .O(N__20974),
            .I(N__20969));
    LocalMux I__2404 (
            .O(N__20969),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2403 (
            .O(N__20966),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__2402 (
            .O(N__20963),
            .I(N__20957));
    InMux I__2401 (
            .O(N__20962),
            .I(N__20957));
    LocalMux I__2400 (
            .O(N__20957),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2399 (
            .O(N__20954),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__2398 (
            .O(N__20951),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__2397 (
            .O(N__20948),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    CascadeMux I__2396 (
            .O(N__20945),
            .I(N__20942));
    InMux I__2395 (
            .O(N__20942),
            .I(N__20939));
    LocalMux I__2394 (
            .O(N__20939),
            .I(N__20935));
    InMux I__2393 (
            .O(N__20938),
            .I(N__20932));
    Span4Mux_h I__2392 (
            .O(N__20935),
            .I(N__20929));
    LocalMux I__2391 (
            .O(N__20932),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    Odrv4 I__2390 (
            .O(N__20929),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2389 (
            .O(N__20924),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    CascadeMux I__2388 (
            .O(N__20921),
            .I(N__20917));
    InMux I__2387 (
            .O(N__20920),
            .I(N__20914));
    InMux I__2386 (
            .O(N__20917),
            .I(N__20911));
    LocalMux I__2385 (
            .O(N__20914),
            .I(N__20908));
    LocalMux I__2384 (
            .O(N__20911),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    Odrv4 I__2383 (
            .O(N__20908),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2382 (
            .O(N__20903),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__2381 (
            .O(N__20900),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__2380 (
            .O(N__20897),
            .I(bfn_5_12_0_));
    InMux I__2379 (
            .O(N__20894),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ));
    InMux I__2378 (
            .O(N__20891),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    CascadeMux I__2377 (
            .O(N__20888),
            .I(N__20884));
    InMux I__2376 (
            .O(N__20887),
            .I(N__20881));
    InMux I__2375 (
            .O(N__20884),
            .I(N__20878));
    LocalMux I__2374 (
            .O(N__20881),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    LocalMux I__2373 (
            .O(N__20878),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2372 (
            .O(N__20873),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__2371 (
            .O(N__20870),
            .I(N__20864));
    InMux I__2370 (
            .O(N__20869),
            .I(N__20864));
    LocalMux I__2369 (
            .O(N__20864),
            .I(N__20860));
    InMux I__2368 (
            .O(N__20863),
            .I(N__20857));
    Odrv4 I__2367 (
            .O(N__20860),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    LocalMux I__2366 (
            .O(N__20857),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2365 (
            .O(N__20852),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__2364 (
            .O(N__20849),
            .I(N__20845));
    InMux I__2363 (
            .O(N__20848),
            .I(N__20842));
    LocalMux I__2362 (
            .O(N__20845),
            .I(N__20839));
    LocalMux I__2361 (
            .O(N__20842),
            .I(N__20836));
    Span4Mux_h I__2360 (
            .O(N__20839),
            .I(N__20831));
    Span4Mux_h I__2359 (
            .O(N__20836),
            .I(N__20828));
    InMux I__2358 (
            .O(N__20835),
            .I(N__20823));
    InMux I__2357 (
            .O(N__20834),
            .I(N__20823));
    Odrv4 I__2356 (
            .O(N__20831),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__2355 (
            .O(N__20828),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    LocalMux I__2354 (
            .O(N__20823),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2353 (
            .O(N__20816),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    CascadeMux I__2352 (
            .O(N__20813),
            .I(N__20810));
    InMux I__2351 (
            .O(N__20810),
            .I(N__20807));
    LocalMux I__2350 (
            .O(N__20807),
            .I(N__20804));
    Span4Mux_h I__2349 (
            .O(N__20804),
            .I(N__20799));
    InMux I__2348 (
            .O(N__20803),
            .I(N__20796));
    InMux I__2347 (
            .O(N__20802),
            .I(N__20793));
    Odrv4 I__2346 (
            .O(N__20799),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    LocalMux I__2345 (
            .O(N__20796),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    LocalMux I__2344 (
            .O(N__20793),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2343 (
            .O(N__20786),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    CascadeMux I__2342 (
            .O(N__20783),
            .I(N__20780));
    InMux I__2341 (
            .O(N__20780),
            .I(N__20775));
    InMux I__2340 (
            .O(N__20779),
            .I(N__20772));
    InMux I__2339 (
            .O(N__20778),
            .I(N__20769));
    LocalMux I__2338 (
            .O(N__20775),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    LocalMux I__2337 (
            .O(N__20772),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    LocalMux I__2336 (
            .O(N__20769),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2335 (
            .O(N__20762),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__2334 (
            .O(N__20759),
            .I(N__20756));
    LocalMux I__2333 (
            .O(N__20756),
            .I(N__20753));
    Span4Mux_h I__2332 (
            .O(N__20753),
            .I(N__20748));
    InMux I__2331 (
            .O(N__20752),
            .I(N__20745));
    InMux I__2330 (
            .O(N__20751),
            .I(N__20742));
    Odrv4 I__2329 (
            .O(N__20748),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    LocalMux I__2328 (
            .O(N__20745),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    LocalMux I__2327 (
            .O(N__20742),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2326 (
            .O(N__20735),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    CascadeMux I__2325 (
            .O(N__20732),
            .I(N__20728));
    InMux I__2324 (
            .O(N__20731),
            .I(N__20724));
    InMux I__2323 (
            .O(N__20728),
            .I(N__20721));
    InMux I__2322 (
            .O(N__20727),
            .I(N__20718));
    LocalMux I__2321 (
            .O(N__20724),
            .I(N__20715));
    LocalMux I__2320 (
            .O(N__20721),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    LocalMux I__2319 (
            .O(N__20718),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__2318 (
            .O(N__20715),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2317 (
            .O(N__20708),
            .I(bfn_5_11_0_));
    InMux I__2316 (
            .O(N__20705),
            .I(N__20701));
    InMux I__2315 (
            .O(N__20704),
            .I(N__20698));
    LocalMux I__2314 (
            .O(N__20701),
            .I(N__20692));
    LocalMux I__2313 (
            .O(N__20698),
            .I(N__20692));
    InMux I__2312 (
            .O(N__20697),
            .I(N__20689));
    Odrv4 I__2311 (
            .O(N__20692),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    LocalMux I__2310 (
            .O(N__20689),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2309 (
            .O(N__20684),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ));
    InMux I__2308 (
            .O(N__20681),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__2307 (
            .O(N__20678),
            .I(N__20675));
    LocalMux I__2306 (
            .O(N__20675),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    CascadeMux I__2305 (
            .O(N__20672),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ));
    InMux I__2304 (
            .O(N__20669),
            .I(N__20658));
    InMux I__2303 (
            .O(N__20668),
            .I(N__20653));
    InMux I__2302 (
            .O(N__20667),
            .I(N__20653));
    InMux I__2301 (
            .O(N__20666),
            .I(N__20646));
    InMux I__2300 (
            .O(N__20665),
            .I(N__20646));
    InMux I__2299 (
            .O(N__20664),
            .I(N__20646));
    InMux I__2298 (
            .O(N__20663),
            .I(N__20643));
    InMux I__2297 (
            .O(N__20662),
            .I(N__20638));
    InMux I__2296 (
            .O(N__20661),
            .I(N__20638));
    LocalMux I__2295 (
            .O(N__20658),
            .I(N__20635));
    LocalMux I__2294 (
            .O(N__20653),
            .I(N__20632));
    LocalMux I__2293 (
            .O(N__20646),
            .I(N__20625));
    LocalMux I__2292 (
            .O(N__20643),
            .I(N__20625));
    LocalMux I__2291 (
            .O(N__20638),
            .I(N__20625));
    Span4Mux_h I__2290 (
            .O(N__20635),
            .I(N__20622));
    Odrv4 I__2289 (
            .O(N__20632),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2288 (
            .O(N__20625),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2287 (
            .O(N__20622),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    InMux I__2286 (
            .O(N__20615),
            .I(N__20612));
    LocalMux I__2285 (
            .O(N__20612),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    InMux I__2284 (
            .O(N__20609),
            .I(N__20606));
    LocalMux I__2283 (
            .O(N__20606),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    InMux I__2282 (
            .O(N__20603),
            .I(N__20600));
    LocalMux I__2281 (
            .O(N__20600),
            .I(N__20597));
    Span4Mux_h I__2280 (
            .O(N__20597),
            .I(N__20594));
    Odrv4 I__2279 (
            .O(N__20594),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_1 ));
    InMux I__2278 (
            .O(N__20591),
            .I(N__20588));
    LocalMux I__2277 (
            .O(N__20588),
            .I(N__20585));
    Span4Mux_h I__2276 (
            .O(N__20585),
            .I(N__20582));
    Odrv4 I__2275 (
            .O(N__20582),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_0 ));
    InMux I__2274 (
            .O(N__20579),
            .I(N__20576));
    LocalMux I__2273 (
            .O(N__20576),
            .I(N__20573));
    Odrv4 I__2272 (
            .O(N__20573),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__2271 (
            .O(N__20570),
            .I(N__20567));
    LocalMux I__2270 (
            .O(N__20567),
            .I(N__20564));
    Odrv4 I__2269 (
            .O(N__20564),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__2268 (
            .O(N__20561),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ));
    InMux I__2267 (
            .O(N__20558),
            .I(N__20555));
    LocalMux I__2266 (
            .O(N__20555),
            .I(N__20552));
    Odrv4 I__2265 (
            .O(N__20552),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2264 (
            .O(N__20549),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__2263 (
            .O(N__20546),
            .I(N__20543));
    LocalMux I__2262 (
            .O(N__20543),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ));
    CascadeMux I__2261 (
            .O(N__20540),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ));
    InMux I__2260 (
            .O(N__20537),
            .I(N__20534));
    LocalMux I__2259 (
            .O(N__20534),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    CascadeMux I__2258 (
            .O(N__20531),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ));
    InMux I__2257 (
            .O(N__20528),
            .I(N__20525));
    LocalMux I__2256 (
            .O(N__20525),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    CascadeMux I__2255 (
            .O(N__20522),
            .I(N__20517));
    CascadeMux I__2254 (
            .O(N__20521),
            .I(N__20512));
    InMux I__2253 (
            .O(N__20520),
            .I(N__20507));
    InMux I__2252 (
            .O(N__20517),
            .I(N__20507));
    InMux I__2251 (
            .O(N__20516),
            .I(N__20499));
    InMux I__2250 (
            .O(N__20515),
            .I(N__20499));
    InMux I__2249 (
            .O(N__20512),
            .I(N__20499));
    LocalMux I__2248 (
            .O(N__20507),
            .I(N__20496));
    InMux I__2247 (
            .O(N__20506),
            .I(N__20492));
    LocalMux I__2246 (
            .O(N__20499),
            .I(N__20487));
    Span4Mux_h I__2245 (
            .O(N__20496),
            .I(N__20487));
    InMux I__2244 (
            .O(N__20495),
            .I(N__20484));
    LocalMux I__2243 (
            .O(N__20492),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv4 I__2242 (
            .O(N__20487),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    LocalMux I__2241 (
            .O(N__20484),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    InMux I__2240 (
            .O(N__20477),
            .I(N__20474));
    LocalMux I__2239 (
            .O(N__20474),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    CascadeMux I__2238 (
            .O(N__20471),
            .I(N__20468));
    InMux I__2237 (
            .O(N__20468),
            .I(N__20465));
    LocalMux I__2236 (
            .O(N__20465),
            .I(N__20462));
    Span4Mux_h I__2235 (
            .O(N__20462),
            .I(N__20459));
    Odrv4 I__2234 (
            .O(N__20459),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9 ));
    InMux I__2233 (
            .O(N__20456),
            .I(N__20453));
    LocalMux I__2232 (
            .O(N__20453),
            .I(N__20448));
    InMux I__2231 (
            .O(N__20452),
            .I(N__20445));
    InMux I__2230 (
            .O(N__20451),
            .I(N__20442));
    Span4Mux_h I__2229 (
            .O(N__20448),
            .I(N__20439));
    LocalMux I__2228 (
            .O(N__20445),
            .I(pwm_duty_input_9));
    LocalMux I__2227 (
            .O(N__20442),
            .I(pwm_duty_input_9));
    Odrv4 I__2226 (
            .O(N__20439),
            .I(pwm_duty_input_9));
    InMux I__2225 (
            .O(N__20432),
            .I(N__20429));
    LocalMux I__2224 (
            .O(N__20429),
            .I(N__20425));
    InMux I__2223 (
            .O(N__20428),
            .I(N__20422));
    Span4Mux_v I__2222 (
            .O(N__20425),
            .I(N__20417));
    LocalMux I__2221 (
            .O(N__20422),
            .I(N__20417));
    Span4Mux_h I__2220 (
            .O(N__20417),
            .I(N__20413));
    InMux I__2219 (
            .O(N__20416),
            .I(N__20410));
    Odrv4 I__2218 (
            .O(N__20413),
            .I(pwm_duty_input_7));
    LocalMux I__2217 (
            .O(N__20410),
            .I(pwm_duty_input_7));
    InMux I__2216 (
            .O(N__20405),
            .I(N__20401));
    CascadeMux I__2215 (
            .O(N__20404),
            .I(N__20398));
    LocalMux I__2214 (
            .O(N__20401),
            .I(N__20394));
    InMux I__2213 (
            .O(N__20398),
            .I(N__20391));
    InMux I__2212 (
            .O(N__20397),
            .I(N__20388));
    Span4Mux_h I__2211 (
            .O(N__20394),
            .I(N__20385));
    LocalMux I__2210 (
            .O(N__20391),
            .I(pwm_duty_input_6));
    LocalMux I__2209 (
            .O(N__20388),
            .I(pwm_duty_input_6));
    Odrv4 I__2208 (
            .O(N__20385),
            .I(pwm_duty_input_6));
    InMux I__2207 (
            .O(N__20378),
            .I(N__20375));
    LocalMux I__2206 (
            .O(N__20375),
            .I(N__20370));
    InMux I__2205 (
            .O(N__20374),
            .I(N__20367));
    InMux I__2204 (
            .O(N__20373),
            .I(N__20364));
    Span4Mux_v I__2203 (
            .O(N__20370),
            .I(N__20361));
    LocalMux I__2202 (
            .O(N__20367),
            .I(pwm_duty_input_8));
    LocalMux I__2201 (
            .O(N__20364),
            .I(pwm_duty_input_8));
    Odrv4 I__2200 (
            .O(N__20361),
            .I(pwm_duty_input_8));
    InMux I__2199 (
            .O(N__20354),
            .I(N__20351));
    LocalMux I__2198 (
            .O(N__20351),
            .I(N__20346));
    InMux I__2197 (
            .O(N__20350),
            .I(N__20343));
    InMux I__2196 (
            .O(N__20349),
            .I(N__20340));
    Span4Mux_h I__2195 (
            .O(N__20346),
            .I(N__20337));
    LocalMux I__2194 (
            .O(N__20343),
            .I(pwm_duty_input_3));
    LocalMux I__2193 (
            .O(N__20340),
            .I(pwm_duty_input_3));
    Odrv4 I__2192 (
            .O(N__20337),
            .I(pwm_duty_input_3));
    InMux I__2191 (
            .O(N__20330),
            .I(N__20325));
    InMux I__2190 (
            .O(N__20329),
            .I(N__20322));
    InMux I__2189 (
            .O(N__20328),
            .I(N__20319));
    LocalMux I__2188 (
            .O(N__20325),
            .I(N__20316));
    LocalMux I__2187 (
            .O(N__20322),
            .I(N__20313));
    LocalMux I__2186 (
            .O(N__20319),
            .I(N__20310));
    Odrv4 I__2185 (
            .O(N__20316),
            .I(pwm_duty_input_4));
    Odrv4 I__2184 (
            .O(N__20313),
            .I(pwm_duty_input_4));
    Odrv12 I__2183 (
            .O(N__20310),
            .I(pwm_duty_input_4));
    CascadeMux I__2182 (
            .O(N__20303),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ));
    InMux I__2181 (
            .O(N__20300),
            .I(N__20297));
    LocalMux I__2180 (
            .O(N__20297),
            .I(N__20293));
    InMux I__2179 (
            .O(N__20296),
            .I(N__20290));
    Span4Mux_v I__2178 (
            .O(N__20293),
            .I(N__20285));
    LocalMux I__2177 (
            .O(N__20290),
            .I(N__20285));
    Span4Mux_h I__2176 (
            .O(N__20285),
            .I(N__20281));
    InMux I__2175 (
            .O(N__20284),
            .I(N__20278));
    Odrv4 I__2174 (
            .O(N__20281),
            .I(pwm_duty_input_5));
    LocalMux I__2173 (
            .O(N__20278),
            .I(pwm_duty_input_5));
    InMux I__2172 (
            .O(N__20273),
            .I(N__20251));
    InMux I__2171 (
            .O(N__20272),
            .I(N__20251));
    InMux I__2170 (
            .O(N__20271),
            .I(N__20251));
    InMux I__2169 (
            .O(N__20270),
            .I(N__20251));
    InMux I__2168 (
            .O(N__20269),
            .I(N__20251));
    InMux I__2167 (
            .O(N__20268),
            .I(N__20251));
    InMux I__2166 (
            .O(N__20267),
            .I(N__20242));
    InMux I__2165 (
            .O(N__20266),
            .I(N__20242));
    InMux I__2164 (
            .O(N__20265),
            .I(N__20242));
    InMux I__2163 (
            .O(N__20264),
            .I(N__20242));
    LocalMux I__2162 (
            .O(N__20251),
            .I(N__20237));
    LocalMux I__2161 (
            .O(N__20242),
            .I(N__20237));
    Odrv4 I__2160 (
            .O(N__20237),
            .I(\pwm_generator_inst.N_17 ));
    CascadeMux I__2159 (
            .O(N__20234),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ));
    CascadeMux I__2158 (
            .O(N__20231),
            .I(N__20228));
    InMux I__2157 (
            .O(N__20228),
            .I(N__20224));
    InMux I__2156 (
            .O(N__20227),
            .I(N__20221));
    LocalMux I__2155 (
            .O(N__20224),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__2154 (
            .O(N__20221),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    CascadeMux I__2153 (
            .O(N__20216),
            .I(N__20213));
    InMux I__2152 (
            .O(N__20213),
            .I(N__20210));
    LocalMux I__2151 (
            .O(N__20210),
            .I(\current_shift_inst.PI_CTRL.N_155 ));
    CascadeMux I__2150 (
            .O(N__20207),
            .I(N__20203));
    InMux I__2149 (
            .O(N__20206),
            .I(N__20200));
    InMux I__2148 (
            .O(N__20203),
            .I(N__20197));
    LocalMux I__2147 (
            .O(N__20200),
            .I(N__20191));
    LocalMux I__2146 (
            .O(N__20197),
            .I(N__20191));
    InMux I__2145 (
            .O(N__20196),
            .I(N__20188));
    Odrv4 I__2144 (
            .O(N__20191),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__2143 (
            .O(N__20188),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    InMux I__2142 (
            .O(N__20183),
            .I(N__20180));
    LocalMux I__2141 (
            .O(N__20180),
            .I(\current_shift_inst.PI_CTRL.N_149 ));
    InMux I__2140 (
            .O(N__20177),
            .I(N__20174));
    LocalMux I__2139 (
            .O(N__20174),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_2 ));
    InMux I__2138 (
            .O(N__20171),
            .I(N__20168));
    LocalMux I__2137 (
            .O(N__20168),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_3 ));
    CascadeMux I__2136 (
            .O(N__20165),
            .I(N__20162));
    InMux I__2135 (
            .O(N__20162),
            .I(N__20159));
    LocalMux I__2134 (
            .O(N__20159),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ));
    CascadeMux I__2133 (
            .O(N__20156),
            .I(N__20153));
    InMux I__2132 (
            .O(N__20153),
            .I(N__20150));
    LocalMux I__2131 (
            .O(N__20150),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ));
    InMux I__2130 (
            .O(N__20147),
            .I(N__20144));
    LocalMux I__2129 (
            .O(N__20144),
            .I(N__20141));
    Odrv4 I__2128 (
            .O(N__20141),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_7 ));
    InMux I__2127 (
            .O(N__20138),
            .I(N__20135));
    LocalMux I__2126 (
            .O(N__20135),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ));
    InMux I__2125 (
            .O(N__20132),
            .I(N__20129));
    LocalMux I__2124 (
            .O(N__20129),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_8 ));
    InMux I__2123 (
            .O(N__20126),
            .I(N__20104));
    InMux I__2122 (
            .O(N__20125),
            .I(N__20104));
    InMux I__2121 (
            .O(N__20124),
            .I(N__20104));
    InMux I__2120 (
            .O(N__20123),
            .I(N__20104));
    InMux I__2119 (
            .O(N__20122),
            .I(N__20104));
    InMux I__2118 (
            .O(N__20121),
            .I(N__20104));
    InMux I__2117 (
            .O(N__20120),
            .I(N__20095));
    InMux I__2116 (
            .O(N__20119),
            .I(N__20095));
    InMux I__2115 (
            .O(N__20118),
            .I(N__20095));
    InMux I__2114 (
            .O(N__20117),
            .I(N__20095));
    LocalMux I__2113 (
            .O(N__20104),
            .I(N__20092));
    LocalMux I__2112 (
            .O(N__20095),
            .I(\pwm_generator_inst.N_16 ));
    Odrv4 I__2111 (
            .O(N__20092),
            .I(\pwm_generator_inst.N_16 ));
    CascadeMux I__2110 (
            .O(N__20087),
            .I(N__20084));
    InMux I__2109 (
            .O(N__20084),
            .I(N__20081));
    LocalMux I__2108 (
            .O(N__20081),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ));
    CascadeMux I__2107 (
            .O(N__20078),
            .I(N__20070));
    CascadeMux I__2106 (
            .O(N__20077),
            .I(N__20059));
    CascadeMux I__2105 (
            .O(N__20076),
            .I(N__20056));
    InMux I__2104 (
            .O(N__20075),
            .I(N__20047));
    InMux I__2103 (
            .O(N__20074),
            .I(N__20047));
    InMux I__2102 (
            .O(N__20073),
            .I(N__20047));
    InMux I__2101 (
            .O(N__20070),
            .I(N__20047));
    CascadeMux I__2100 (
            .O(N__20069),
            .I(N__20042));
    InMux I__2099 (
            .O(N__20068),
            .I(N__20035));
    InMux I__2098 (
            .O(N__20067),
            .I(N__20035));
    InMux I__2097 (
            .O(N__20066),
            .I(N__20035));
    InMux I__2096 (
            .O(N__20065),
            .I(N__20022));
    InMux I__2095 (
            .O(N__20064),
            .I(N__20022));
    InMux I__2094 (
            .O(N__20063),
            .I(N__20022));
    InMux I__2093 (
            .O(N__20062),
            .I(N__20022));
    InMux I__2092 (
            .O(N__20059),
            .I(N__20022));
    InMux I__2091 (
            .O(N__20056),
            .I(N__20022));
    LocalMux I__2090 (
            .O(N__20047),
            .I(N__20019));
    InMux I__2089 (
            .O(N__20046),
            .I(N__20014));
    InMux I__2088 (
            .O(N__20045),
            .I(N__20014));
    InMux I__2087 (
            .O(N__20042),
            .I(N__20011));
    LocalMux I__2086 (
            .O(N__20035),
            .I(N__20008));
    LocalMux I__2085 (
            .O(N__20022),
            .I(N__20005));
    Span4Mux_h I__2084 (
            .O(N__20019),
            .I(N__19984));
    LocalMux I__2083 (
            .O(N__20014),
            .I(N__19984));
    LocalMux I__2082 (
            .O(N__20011),
            .I(N__19979));
    Span4Mux_s1_h I__2081 (
            .O(N__20008),
            .I(N__19979));
    Span4Mux_h I__2080 (
            .O(N__20005),
            .I(N__19976));
    InMux I__2079 (
            .O(N__20004),
            .I(N__19973));
    InMux I__2078 (
            .O(N__20003),
            .I(N__19956));
    InMux I__2077 (
            .O(N__20002),
            .I(N__19956));
    InMux I__2076 (
            .O(N__20001),
            .I(N__19956));
    InMux I__2075 (
            .O(N__20000),
            .I(N__19956));
    InMux I__2074 (
            .O(N__19999),
            .I(N__19956));
    InMux I__2073 (
            .O(N__19998),
            .I(N__19956));
    InMux I__2072 (
            .O(N__19997),
            .I(N__19956));
    InMux I__2071 (
            .O(N__19996),
            .I(N__19956));
    InMux I__2070 (
            .O(N__19995),
            .I(N__19941));
    InMux I__2069 (
            .O(N__19994),
            .I(N__19941));
    InMux I__2068 (
            .O(N__19993),
            .I(N__19941));
    InMux I__2067 (
            .O(N__19992),
            .I(N__19941));
    InMux I__2066 (
            .O(N__19991),
            .I(N__19941));
    InMux I__2065 (
            .O(N__19990),
            .I(N__19941));
    InMux I__2064 (
            .O(N__19989),
            .I(N__19941));
    Span4Mux_v I__2063 (
            .O(N__19984),
            .I(N__19936));
    Span4Mux_v I__2062 (
            .O(N__19979),
            .I(N__19936));
    Odrv4 I__2061 (
            .O(N__19976),
            .I(N_19_1));
    LocalMux I__2060 (
            .O(N__19973),
            .I(N_19_1));
    LocalMux I__2059 (
            .O(N__19956),
            .I(N_19_1));
    LocalMux I__2058 (
            .O(N__19941),
            .I(N_19_1));
    Odrv4 I__2057 (
            .O(N__19936),
            .I(N_19_1));
    CascadeMux I__2056 (
            .O(N__19925),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    InMux I__2055 (
            .O(N__19922),
            .I(N__19916));
    InMux I__2054 (
            .O(N__19921),
            .I(N__19916));
    LocalMux I__2053 (
            .O(N__19916),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    InMux I__2052 (
            .O(N__19913),
            .I(N__19910));
    LocalMux I__2051 (
            .O(N__19910),
            .I(N__19906));
    InMux I__2050 (
            .O(N__19909),
            .I(N__19903));
    Span4Mux_s3_h I__2049 (
            .O(N__19906),
            .I(N__19900));
    LocalMux I__2048 (
            .O(N__19903),
            .I(pwm_duty_input_2));
    Odrv4 I__2047 (
            .O(N__19900),
            .I(pwm_duty_input_2));
    InMux I__2046 (
            .O(N__19895),
            .I(N__19889));
    InMux I__2045 (
            .O(N__19894),
            .I(N__19889));
    LocalMux I__2044 (
            .O(N__19889),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__2043 (
            .O(N__19886),
            .I(N__19883));
    LocalMux I__2042 (
            .O(N__19883),
            .I(N__19879));
    InMux I__2041 (
            .O(N__19882),
            .I(N__19876));
    Span4Mux_s3_h I__2040 (
            .O(N__19879),
            .I(N__19873));
    LocalMux I__2039 (
            .O(N__19876),
            .I(pwm_duty_input_1));
    Odrv4 I__2038 (
            .O(N__19873),
            .I(pwm_duty_input_1));
    CascadeMux I__2037 (
            .O(N__19868),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ));
    InMux I__2036 (
            .O(N__19865),
            .I(N__19862));
    LocalMux I__2035 (
            .O(N__19862),
            .I(N__19859));
    Odrv4 I__2034 (
            .O(N__19859),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ));
    CascadeMux I__2033 (
            .O(N__19856),
            .I(N__19850));
    CascadeMux I__2032 (
            .O(N__19855),
            .I(N__19846));
    CascadeMux I__2031 (
            .O(N__19854),
            .I(N__19843));
    CascadeMux I__2030 (
            .O(N__19853),
            .I(N__19840));
    InMux I__2029 (
            .O(N__19850),
            .I(N__19835));
    InMux I__2028 (
            .O(N__19849),
            .I(N__19835));
    InMux I__2027 (
            .O(N__19846),
            .I(N__19828));
    InMux I__2026 (
            .O(N__19843),
            .I(N__19828));
    InMux I__2025 (
            .O(N__19840),
            .I(N__19828));
    LocalMux I__2024 (
            .O(N__19835),
            .I(\current_shift_inst.PI_CTRL.N_153 ));
    LocalMux I__2023 (
            .O(N__19828),
            .I(\current_shift_inst.PI_CTRL.N_153 ));
    InMux I__2022 (
            .O(N__19823),
            .I(N__19814));
    InMux I__2021 (
            .O(N__19822),
            .I(N__19814));
    InMux I__2020 (
            .O(N__19821),
            .I(N__19814));
    LocalMux I__2019 (
            .O(N__19814),
            .I(\current_shift_inst.PI_CTRL.N_154 ));
    InMux I__2018 (
            .O(N__19811),
            .I(N__19808));
    LocalMux I__2017 (
            .O(N__19808),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_6 ));
    InMux I__2016 (
            .O(N__19805),
            .I(N__19802));
    LocalMux I__2015 (
            .O(N__19802),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ));
    InMux I__2014 (
            .O(N__19799),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_5 ));
    InMux I__2013 (
            .O(N__19796),
            .I(N__19793));
    LocalMux I__2012 (
            .O(N__19793),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_7 ));
    InMux I__2011 (
            .O(N__19790),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_6 ));
    InMux I__2010 (
            .O(N__19787),
            .I(N__19784));
    LocalMux I__2009 (
            .O(N__19784),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_8 ));
    InMux I__2008 (
            .O(N__19781),
            .I(bfn_3_9_0_));
    InMux I__2007 (
            .O(N__19778),
            .I(N__19775));
    LocalMux I__2006 (
            .O(N__19775),
            .I(N__19772));
    Odrv4 I__2005 (
            .O(N__19772),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ));
    InMux I__2004 (
            .O(N__19769),
            .I(N__19766));
    LocalMux I__2003 (
            .O(N__19766),
            .I(N__19763));
    Odrv4 I__2002 (
            .O(N__19763),
            .I(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ));
    CascadeMux I__2001 (
            .O(N__19760),
            .I(N__19755));
    CascadeMux I__2000 (
            .O(N__19759),
            .I(N__19750));
    CascadeMux I__1999 (
            .O(N__19758),
            .I(N__19745));
    InMux I__1998 (
            .O(N__19755),
            .I(N__19741));
    InMux I__1997 (
            .O(N__19754),
            .I(N__19738));
    InMux I__1996 (
            .O(N__19753),
            .I(N__19735));
    InMux I__1995 (
            .O(N__19750),
            .I(N__19732));
    InMux I__1994 (
            .O(N__19749),
            .I(N__19727));
    InMux I__1993 (
            .O(N__19748),
            .I(N__19727));
    InMux I__1992 (
            .O(N__19745),
            .I(N__19723));
    CascadeMux I__1991 (
            .O(N__19744),
            .I(N__19720));
    LocalMux I__1990 (
            .O(N__19741),
            .I(N__19714));
    LocalMux I__1989 (
            .O(N__19738),
            .I(N__19711));
    LocalMux I__1988 (
            .O(N__19735),
            .I(N__19704));
    LocalMux I__1987 (
            .O(N__19732),
            .I(N__19704));
    LocalMux I__1986 (
            .O(N__19727),
            .I(N__19704));
    InMux I__1985 (
            .O(N__19726),
            .I(N__19701));
    LocalMux I__1984 (
            .O(N__19723),
            .I(N__19698));
    InMux I__1983 (
            .O(N__19720),
            .I(N__19689));
    InMux I__1982 (
            .O(N__19719),
            .I(N__19689));
    InMux I__1981 (
            .O(N__19718),
            .I(N__19689));
    InMux I__1980 (
            .O(N__19717),
            .I(N__19689));
    Span4Mux_h I__1979 (
            .O(N__19714),
            .I(N__19680));
    Span4Mux_v I__1978 (
            .O(N__19711),
            .I(N__19680));
    Span4Mux_h I__1977 (
            .O(N__19704),
            .I(N__19680));
    LocalMux I__1976 (
            .O(N__19701),
            .I(N__19680));
    Span4Mux_h I__1975 (
            .O(N__19698),
            .I(N__19677));
    LocalMux I__1974 (
            .O(N__19689),
            .I(N__19672));
    Span4Mux_s2_h I__1973 (
            .O(N__19680),
            .I(N__19672));
    Odrv4 I__1972 (
            .O(N__19677),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__1971 (
            .O(N__19672),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    InMux I__1970 (
            .O(N__19667),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_8 ));
    CascadeMux I__1969 (
            .O(N__19664),
            .I(\pwm_generator_inst.un1_duty_inputlt3_cascade_ ));
    CascadeMux I__1968 (
            .O(N__19661),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3_cascade_ ));
    InMux I__1967 (
            .O(N__19658),
            .I(N__19655));
    LocalMux I__1966 (
            .O(N__19655),
            .I(N__19651));
    InMux I__1965 (
            .O(N__19654),
            .I(N__19648));
    Span4Mux_v I__1964 (
            .O(N__19651),
            .I(N__19645));
    LocalMux I__1963 (
            .O(N__19648),
            .I(pwm_duty_input_0));
    Odrv4 I__1962 (
            .O(N__19645),
            .I(pwm_duty_input_0));
    InMux I__1961 (
            .O(N__19640),
            .I(N__19637));
    LocalMux I__1960 (
            .O(N__19637),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_5 ));
    InMux I__1959 (
            .O(N__19634),
            .I(N__19631));
    LocalMux I__1958 (
            .O(N__19631),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_0 ));
    CascadeMux I__1957 (
            .O(N__19628),
            .I(N__19625));
    InMux I__1956 (
            .O(N__19625),
            .I(N__19622));
    LocalMux I__1955 (
            .O(N__19622),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ));
    InMux I__1954 (
            .O(N__19619),
            .I(N__19616));
    LocalMux I__1953 (
            .O(N__19616),
            .I(N__19613));
    Odrv4 I__1952 (
            .O(N__19613),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_1 ));
    CascadeMux I__1951 (
            .O(N__19610),
            .I(N__19607));
    InMux I__1950 (
            .O(N__19607),
            .I(N__19604));
    LocalMux I__1949 (
            .O(N__19604),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ));
    InMux I__1948 (
            .O(N__19601),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_0 ));
    InMux I__1947 (
            .O(N__19598),
            .I(N__19595));
    LocalMux I__1946 (
            .O(N__19595),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_2 ));
    CascadeMux I__1945 (
            .O(N__19592),
            .I(N__19589));
    InMux I__1944 (
            .O(N__19589),
            .I(N__19586));
    LocalMux I__1943 (
            .O(N__19586),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ));
    InMux I__1942 (
            .O(N__19583),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_1 ));
    InMux I__1941 (
            .O(N__19580),
            .I(N__19577));
    LocalMux I__1940 (
            .O(N__19577),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_3 ));
    CascadeMux I__1939 (
            .O(N__19574),
            .I(N__19571));
    InMux I__1938 (
            .O(N__19571),
            .I(N__19568));
    LocalMux I__1937 (
            .O(N__19568),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ));
    InMux I__1936 (
            .O(N__19565),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_2 ));
    InMux I__1935 (
            .O(N__19562),
            .I(N__19559));
    LocalMux I__1934 (
            .O(N__19559),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_4 ));
    InMux I__1933 (
            .O(N__19556),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_3 ));
    InMux I__1932 (
            .O(N__19553),
            .I(N__19550));
    LocalMux I__1931 (
            .O(N__19550),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_5 ));
    InMux I__1930 (
            .O(N__19547),
            .I(N__19544));
    LocalMux I__1929 (
            .O(N__19544),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ));
    InMux I__1928 (
            .O(N__19541),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_4 ));
    InMux I__1927 (
            .O(N__19538),
            .I(N__19535));
    LocalMux I__1926 (
            .O(N__19535),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ));
    InMux I__1925 (
            .O(N__19532),
            .I(N__19529));
    LocalMux I__1924 (
            .O(N__19529),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ));
    InMux I__1923 (
            .O(N__19526),
            .I(N__19523));
    LocalMux I__1922 (
            .O(N__19523),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ));
    InMux I__1921 (
            .O(N__19520),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19 ));
    InMux I__1920 (
            .O(N__19517),
            .I(N__19514));
    LocalMux I__1919 (
            .O(N__19514),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ));
    InMux I__1918 (
            .O(N__19511),
            .I(N__19508));
    LocalMux I__1917 (
            .O(N__19508),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ));
    InMux I__1916 (
            .O(N__19505),
            .I(N__19502));
    LocalMux I__1915 (
            .O(N__19502),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ));
    InMux I__1914 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__1913 (
            .O(N__19496),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ));
    InMux I__1912 (
            .O(N__19493),
            .I(N__19490));
    LocalMux I__1911 (
            .O(N__19490),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ));
    InMux I__1910 (
            .O(N__19487),
            .I(N__19484));
    LocalMux I__1909 (
            .O(N__19484),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ));
    InMux I__1908 (
            .O(N__19481),
            .I(N__19478));
    LocalMux I__1907 (
            .O(N__19478),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ));
    InMux I__1906 (
            .O(N__19475),
            .I(N__19472));
    LocalMux I__1905 (
            .O(N__19472),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ));
    InMux I__1904 (
            .O(N__19469),
            .I(N__19466));
    LocalMux I__1903 (
            .O(N__19466),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ));
    InMux I__1902 (
            .O(N__19463),
            .I(N__19460));
    LocalMux I__1901 (
            .O(N__19460),
            .I(N__19457));
    Span4Mux_h I__1900 (
            .O(N__19457),
            .I(N__19454));
    Odrv4 I__1899 (
            .O(N__19454),
            .I(\pwm_generator_inst.O_12 ));
    CascadeMux I__1898 (
            .O(N__19451),
            .I(N__19448));
    InMux I__1897 (
            .O(N__19448),
            .I(N__19442));
    InMux I__1896 (
            .O(N__19447),
            .I(N__19442));
    LocalMux I__1895 (
            .O(N__19442),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    InMux I__1894 (
            .O(N__19439),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0 ));
    InMux I__1893 (
            .O(N__19436),
            .I(N__19433));
    LocalMux I__1892 (
            .O(N__19433),
            .I(N__19430));
    Span4Mux_v I__1891 (
            .O(N__19430),
            .I(N__19427));
    Odrv4 I__1890 (
            .O(N__19427),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1889 (
            .O(N__19424),
            .I(N__19418));
    InMux I__1888 (
            .O(N__19423),
            .I(N__19418));
    LocalMux I__1887 (
            .O(N__19418),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    InMux I__1886 (
            .O(N__19415),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1 ));
    InMux I__1885 (
            .O(N__19412),
            .I(N__19409));
    LocalMux I__1884 (
            .O(N__19409),
            .I(N__19406));
    Span4Mux_h I__1883 (
            .O(N__19406),
            .I(N__19403));
    Odrv4 I__1882 (
            .O(N__19403),
            .I(\pwm_generator_inst.O_14 ));
    CascadeMux I__1881 (
            .O(N__19400),
            .I(N__19397));
    InMux I__1880 (
            .O(N__19397),
            .I(N__19393));
    InMux I__1879 (
            .O(N__19396),
            .I(N__19390));
    LocalMux I__1878 (
            .O(N__19393),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    LocalMux I__1877 (
            .O(N__19390),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    InMux I__1876 (
            .O(N__19385),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2 ));
    InMux I__1875 (
            .O(N__19382),
            .I(N__19379));
    LocalMux I__1874 (
            .O(N__19379),
            .I(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ));
    CascadeMux I__1873 (
            .O(N__19376),
            .I(N__19373));
    InMux I__1872 (
            .O(N__19373),
            .I(N__19370));
    LocalMux I__1871 (
            .O(N__19370),
            .I(N__19366));
    InMux I__1870 (
            .O(N__19369),
            .I(N__19363));
    Odrv4 I__1869 (
            .O(N__19366),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    LocalMux I__1868 (
            .O(N__19363),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    InMux I__1867 (
            .O(N__19358),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3 ));
    CascadeMux I__1866 (
            .O(N__19355),
            .I(N__19352));
    InMux I__1865 (
            .O(N__19352),
            .I(N__19349));
    LocalMux I__1864 (
            .O(N__19349),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ));
    InMux I__1863 (
            .O(N__19346),
            .I(N__19340));
    InMux I__1862 (
            .O(N__19345),
            .I(N__19340));
    LocalMux I__1861 (
            .O(N__19340),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    InMux I__1860 (
            .O(N__19337),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4 ));
    InMux I__1859 (
            .O(N__19334),
            .I(N__19331));
    LocalMux I__1858 (
            .O(N__19331),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ));
    InMux I__1857 (
            .O(N__19328),
            .I(N__19324));
    InMux I__1856 (
            .O(N__19327),
            .I(N__19321));
    LocalMux I__1855 (
            .O(N__19324),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    LocalMux I__1854 (
            .O(N__19321),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    InMux I__1853 (
            .O(N__19316),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5 ));
    CascadeMux I__1852 (
            .O(N__19313),
            .I(N__19310));
    InMux I__1851 (
            .O(N__19310),
            .I(N__19307));
    LocalMux I__1850 (
            .O(N__19307),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ));
    InMux I__1849 (
            .O(N__19304),
            .I(N__19301));
    LocalMux I__1848 (
            .O(N__19301),
            .I(N__19297));
    InMux I__1847 (
            .O(N__19300),
            .I(N__19294));
    Odrv4 I__1846 (
            .O(N__19297),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    LocalMux I__1845 (
            .O(N__19294),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    InMux I__1844 (
            .O(N__19289),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6 ));
    InMux I__1843 (
            .O(N__19286),
            .I(N__19283));
    LocalMux I__1842 (
            .O(N__19283),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ));
    InMux I__1841 (
            .O(N__19280),
            .I(bfn_2_11_0_));
    InMux I__1840 (
            .O(N__19277),
            .I(N__19274));
    LocalMux I__1839 (
            .O(N__19274),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ));
    InMux I__1838 (
            .O(N__19271),
            .I(N__19266));
    InMux I__1837 (
            .O(N__19270),
            .I(N__19263));
    InMux I__1836 (
            .O(N__19269),
            .I(N__19260));
    LocalMux I__1835 (
            .O(N__19266),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    LocalMux I__1834 (
            .O(N__19263),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    LocalMux I__1833 (
            .O(N__19260),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    InMux I__1832 (
            .O(N__19253),
            .I(N__19249));
    InMux I__1831 (
            .O(N__19252),
            .I(N__19246));
    LocalMux I__1830 (
            .O(N__19249),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    LocalMux I__1829 (
            .O(N__19246),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    InMux I__1828 (
            .O(N__19241),
            .I(N__19238));
    LocalMux I__1827 (
            .O(N__19238),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ));
    CascadeMux I__1826 (
            .O(N__19235),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13_cascade_ ));
    InMux I__1825 (
            .O(N__19232),
            .I(N__19228));
    InMux I__1824 (
            .O(N__19231),
            .I(N__19225));
    LocalMux I__1823 (
            .O(N__19228),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    LocalMux I__1822 (
            .O(N__19225),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    InMux I__1821 (
            .O(N__19220),
            .I(N__19217));
    LocalMux I__1820 (
            .O(N__19217),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ));
    CascadeMux I__1819 (
            .O(N__19214),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ));
    InMux I__1818 (
            .O(N__19211),
            .I(N__19208));
    LocalMux I__1817 (
            .O(N__19208),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ));
    InMux I__1816 (
            .O(N__19205),
            .I(N__19198));
    InMux I__1815 (
            .O(N__19204),
            .I(N__19198));
    InMux I__1814 (
            .O(N__19203),
            .I(N__19195));
    LocalMux I__1813 (
            .O(N__19198),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    LocalMux I__1812 (
            .O(N__19195),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    InMux I__1811 (
            .O(N__19190),
            .I(N__19187));
    LocalMux I__1810 (
            .O(N__19187),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ));
    InMux I__1809 (
            .O(N__19184),
            .I(N__19179));
    InMux I__1808 (
            .O(N__19183),
            .I(N__19174));
    InMux I__1807 (
            .O(N__19182),
            .I(N__19174));
    LocalMux I__1806 (
            .O(N__19179),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    LocalMux I__1805 (
            .O(N__19174),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    InMux I__1804 (
            .O(N__19169),
            .I(N__19165));
    InMux I__1803 (
            .O(N__19168),
            .I(N__19162));
    LocalMux I__1802 (
            .O(N__19165),
            .I(N__19159));
    LocalMux I__1801 (
            .O(N__19162),
            .I(N__19156));
    Span4Mux_v I__1800 (
            .O(N__19159),
            .I(N__19153));
    Span4Mux_h I__1799 (
            .O(N__19156),
            .I(N__19150));
    Odrv4 I__1798 (
            .O(N__19153),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    Odrv4 I__1797 (
            .O(N__19150),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    InMux I__1796 (
            .O(N__19145),
            .I(N__19142));
    LocalMux I__1795 (
            .O(N__19142),
            .I(N__19139));
    Span4Mux_v I__1794 (
            .O(N__19139),
            .I(N__19135));
    InMux I__1793 (
            .O(N__19138),
            .I(N__19132));
    Odrv4 I__1792 (
            .O(N__19135),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    LocalMux I__1791 (
            .O(N__19132),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    InMux I__1790 (
            .O(N__19127),
            .I(N__19121));
    CascadeMux I__1789 (
            .O(N__19126),
            .I(N__19117));
    CascadeMux I__1788 (
            .O(N__19125),
            .I(N__19113));
    CascadeMux I__1787 (
            .O(N__19124),
            .I(N__19109));
    LocalMux I__1786 (
            .O(N__19121),
            .I(N__19106));
    InMux I__1785 (
            .O(N__19120),
            .I(N__19092));
    InMux I__1784 (
            .O(N__19117),
            .I(N__19092));
    InMux I__1783 (
            .O(N__19116),
            .I(N__19092));
    InMux I__1782 (
            .O(N__19113),
            .I(N__19092));
    InMux I__1781 (
            .O(N__19112),
            .I(N__19092));
    InMux I__1780 (
            .O(N__19109),
            .I(N__19092));
    Span4Mux_v I__1779 (
            .O(N__19106),
            .I(N__19089));
    InMux I__1778 (
            .O(N__19105),
            .I(N__19086));
    LocalMux I__1777 (
            .O(N__19092),
            .I(N__19083));
    Odrv4 I__1776 (
            .O(N__19089),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    LocalMux I__1775 (
            .O(N__19086),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    Odrv4 I__1774 (
            .O(N__19083),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    InMux I__1773 (
            .O(N__19076),
            .I(N__19073));
    LocalMux I__1772 (
            .O(N__19073),
            .I(N__19070));
    Span4Mux_v I__1771 (
            .O(N__19070),
            .I(N__19067));
    Odrv4 I__1770 (
            .O(N__19067),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_16 ));
    InMux I__1769 (
            .O(N__19064),
            .I(N__19061));
    LocalMux I__1768 (
            .O(N__19061),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ));
    InMux I__1767 (
            .O(N__19058),
            .I(N__19055));
    LocalMux I__1766 (
            .O(N__19055),
            .I(rgb_drv_RNOZ0));
    InMux I__1765 (
            .O(N__19052),
            .I(N__19049));
    LocalMux I__1764 (
            .O(N__19049),
            .I(N_38_i_i));
    InMux I__1763 (
            .O(N__19046),
            .I(N__19039));
    InMux I__1762 (
            .O(N__19045),
            .I(N__19039));
    InMux I__1761 (
            .O(N__19044),
            .I(N__19036));
    LocalMux I__1760 (
            .O(N__19039),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    LocalMux I__1759 (
            .O(N__19036),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    InMux I__1758 (
            .O(N__19031),
            .I(N__19028));
    LocalMux I__1757 (
            .O(N__19028),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ));
    InMux I__1756 (
            .O(N__19025),
            .I(N__19021));
    InMux I__1755 (
            .O(N__19024),
            .I(N__19018));
    LocalMux I__1754 (
            .O(N__19021),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    LocalMux I__1753 (
            .O(N__19018),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    InMux I__1752 (
            .O(N__19013),
            .I(N__19007));
    InMux I__1751 (
            .O(N__19012),
            .I(N__19007));
    LocalMux I__1750 (
            .O(N__19007),
            .I(N__19004));
    Span4Mux_h I__1749 (
            .O(N__19004),
            .I(N__19001));
    Odrv4 I__1748 (
            .O(N__19001),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__1747 (
            .O(N__18998),
            .I(N__18995));
    LocalMux I__1746 (
            .O(N__18995),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ));
    CascadeMux I__1745 (
            .O(N__18992),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_ ));
    InMux I__1744 (
            .O(N__18989),
            .I(N__18986));
    LocalMux I__1743 (
            .O(N__18986),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ));
    InMux I__1742 (
            .O(N__18983),
            .I(N__18978));
    InMux I__1741 (
            .O(N__18982),
            .I(N__18975));
    InMux I__1740 (
            .O(N__18981),
            .I(N__18972));
    LocalMux I__1739 (
            .O(N__18978),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    LocalMux I__1738 (
            .O(N__18975),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    LocalMux I__1737 (
            .O(N__18972),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    InMux I__1736 (
            .O(N__18965),
            .I(N__18962));
    LocalMux I__1735 (
            .O(N__18962),
            .I(N__18959));
    Span4Mux_v I__1734 (
            .O(N__18959),
            .I(N__18956));
    Odrv4 I__1733 (
            .O(N__18956),
            .I(\pwm_generator_inst.un2_threshold_acc_2_9 ));
    CascadeMux I__1732 (
            .O(N__18953),
            .I(N__18950));
    InMux I__1731 (
            .O(N__18950),
            .I(N__18947));
    LocalMux I__1730 (
            .O(N__18947),
            .I(N__18944));
    Odrv4 I__1729 (
            .O(N__18944),
            .I(\pwm_generator_inst.un2_threshold_acc_1_24 ));
    InMux I__1728 (
            .O(N__18941),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ));
    InMux I__1727 (
            .O(N__18938),
            .I(N__18935));
    LocalMux I__1726 (
            .O(N__18935),
            .I(N__18932));
    Span4Mux_v I__1725 (
            .O(N__18932),
            .I(N__18929));
    Odrv4 I__1724 (
            .O(N__18929),
            .I(\pwm_generator_inst.un2_threshold_acc_2_10 ));
    InMux I__1723 (
            .O(N__18926),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ));
    CascadeMux I__1722 (
            .O(N__18923),
            .I(N__18920));
    InMux I__1721 (
            .O(N__18920),
            .I(N__18917));
    LocalMux I__1720 (
            .O(N__18917),
            .I(N__18914));
    Span4Mux_v I__1719 (
            .O(N__18914),
            .I(N__18911));
    Odrv4 I__1718 (
            .O(N__18911),
            .I(\pwm_generator_inst.un2_threshold_acc_2_11 ));
    InMux I__1717 (
            .O(N__18908),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ));
    InMux I__1716 (
            .O(N__18905),
            .I(N__18902));
    LocalMux I__1715 (
            .O(N__18902),
            .I(N__18899));
    Span4Mux_v I__1714 (
            .O(N__18899),
            .I(N__18896));
    Odrv4 I__1713 (
            .O(N__18896),
            .I(\pwm_generator_inst.un2_threshold_acc_2_12 ));
    InMux I__1712 (
            .O(N__18893),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ));
    CascadeMux I__1711 (
            .O(N__18890),
            .I(N__18887));
    InMux I__1710 (
            .O(N__18887),
            .I(N__18884));
    LocalMux I__1709 (
            .O(N__18884),
            .I(N__18881));
    Span4Mux_v I__1708 (
            .O(N__18881),
            .I(N__18878));
    Odrv4 I__1707 (
            .O(N__18878),
            .I(\pwm_generator_inst.un2_threshold_acc_2_13 ));
    InMux I__1706 (
            .O(N__18875),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ));
    InMux I__1705 (
            .O(N__18872),
            .I(N__18869));
    LocalMux I__1704 (
            .O(N__18869),
            .I(N__18866));
    Span4Mux_v I__1703 (
            .O(N__18866),
            .I(N__18863));
    Odrv4 I__1702 (
            .O(N__18863),
            .I(\pwm_generator_inst.un2_threshold_acc_2_14 ));
    InMux I__1701 (
            .O(N__18860),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ));
    CascadeMux I__1700 (
            .O(N__18857),
            .I(N__18854));
    InMux I__1699 (
            .O(N__18854),
            .I(N__18851));
    LocalMux I__1698 (
            .O(N__18851),
            .I(N__18848));
    Odrv12 I__1697 (
            .O(N__18848),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ));
    InMux I__1696 (
            .O(N__18845),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ));
    InMux I__1695 (
            .O(N__18842),
            .I(bfn_1_12_0_));
    InMux I__1694 (
            .O(N__18839),
            .I(N__18836));
    LocalMux I__1693 (
            .O(N__18836),
            .I(N__18833));
    Span4Mux_v I__1692 (
            .O(N__18833),
            .I(N__18830));
    Odrv4 I__1691 (
            .O(N__18830),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1 ));
    CascadeMux I__1690 (
            .O(N__18827),
            .I(N__18824));
    InMux I__1689 (
            .O(N__18824),
            .I(N__18821));
    LocalMux I__1688 (
            .O(N__18821),
            .I(N__18818));
    Odrv4 I__1687 (
            .O(N__18818),
            .I(\pwm_generator_inst.un2_threshold_acc_1_16 ));
    InMux I__1686 (
            .O(N__18815),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ));
    InMux I__1685 (
            .O(N__18812),
            .I(N__18809));
    LocalMux I__1684 (
            .O(N__18809),
            .I(N__18806));
    Span4Mux_v I__1683 (
            .O(N__18806),
            .I(N__18803));
    Odrv4 I__1682 (
            .O(N__18803),
            .I(\pwm_generator_inst.un2_threshold_acc_2_2 ));
    CascadeMux I__1681 (
            .O(N__18800),
            .I(N__18797));
    InMux I__1680 (
            .O(N__18797),
            .I(N__18794));
    LocalMux I__1679 (
            .O(N__18794),
            .I(N__18791));
    Odrv4 I__1678 (
            .O(N__18791),
            .I(\pwm_generator_inst.un2_threshold_acc_1_17 ));
    InMux I__1677 (
            .O(N__18788),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ));
    InMux I__1676 (
            .O(N__18785),
            .I(N__18782));
    LocalMux I__1675 (
            .O(N__18782),
            .I(N__18779));
    Span4Mux_v I__1674 (
            .O(N__18779),
            .I(N__18776));
    Odrv4 I__1673 (
            .O(N__18776),
            .I(\pwm_generator_inst.un2_threshold_acc_2_3 ));
    CascadeMux I__1672 (
            .O(N__18773),
            .I(N__18770));
    InMux I__1671 (
            .O(N__18770),
            .I(N__18767));
    LocalMux I__1670 (
            .O(N__18767),
            .I(N__18764));
    Odrv4 I__1669 (
            .O(N__18764),
            .I(\pwm_generator_inst.un2_threshold_acc_1_18 ));
    InMux I__1668 (
            .O(N__18761),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ));
    InMux I__1667 (
            .O(N__18758),
            .I(N__18755));
    LocalMux I__1666 (
            .O(N__18755),
            .I(N__18752));
    Span4Mux_v I__1665 (
            .O(N__18752),
            .I(N__18749));
    Odrv4 I__1664 (
            .O(N__18749),
            .I(\pwm_generator_inst.un2_threshold_acc_1_19 ));
    CascadeMux I__1663 (
            .O(N__18746),
            .I(N__18743));
    InMux I__1662 (
            .O(N__18743),
            .I(N__18740));
    LocalMux I__1661 (
            .O(N__18740),
            .I(N__18737));
    Span4Mux_v I__1660 (
            .O(N__18737),
            .I(N__18734));
    Span4Mux_v I__1659 (
            .O(N__18734),
            .I(N__18731));
    Odrv4 I__1658 (
            .O(N__18731),
            .I(\pwm_generator_inst.un2_threshold_acc_2_4 ));
    InMux I__1657 (
            .O(N__18728),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ));
    InMux I__1656 (
            .O(N__18725),
            .I(N__18722));
    LocalMux I__1655 (
            .O(N__18722),
            .I(N__18719));
    Span4Mux_v I__1654 (
            .O(N__18719),
            .I(N__18716));
    Odrv4 I__1653 (
            .O(N__18716),
            .I(\pwm_generator_inst.un2_threshold_acc_2_5 ));
    CascadeMux I__1652 (
            .O(N__18713),
            .I(N__18710));
    InMux I__1651 (
            .O(N__18710),
            .I(N__18707));
    LocalMux I__1650 (
            .O(N__18707),
            .I(N__18704));
    Span4Mux_h I__1649 (
            .O(N__18704),
            .I(N__18701));
    Odrv4 I__1648 (
            .O(N__18701),
            .I(\pwm_generator_inst.un2_threshold_acc_1_20 ));
    InMux I__1647 (
            .O(N__18698),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ));
    InMux I__1646 (
            .O(N__18695),
            .I(N__18692));
    LocalMux I__1645 (
            .O(N__18692),
            .I(N__18689));
    Span4Mux_v I__1644 (
            .O(N__18689),
            .I(N__18686));
    Odrv4 I__1643 (
            .O(N__18686),
            .I(\pwm_generator_inst.un2_threshold_acc_2_6 ));
    CascadeMux I__1642 (
            .O(N__18683),
            .I(N__18680));
    InMux I__1641 (
            .O(N__18680),
            .I(N__18677));
    LocalMux I__1640 (
            .O(N__18677),
            .I(N__18674));
    Span4Mux_h I__1639 (
            .O(N__18674),
            .I(N__18671));
    Odrv4 I__1638 (
            .O(N__18671),
            .I(\pwm_generator_inst.un2_threshold_acc_1_21 ));
    InMux I__1637 (
            .O(N__18668),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ));
    InMux I__1636 (
            .O(N__18665),
            .I(N__18662));
    LocalMux I__1635 (
            .O(N__18662),
            .I(N__18659));
    Span4Mux_v I__1634 (
            .O(N__18659),
            .I(N__18656));
    Odrv4 I__1633 (
            .O(N__18656),
            .I(\pwm_generator_inst.un2_threshold_acc_2_7 ));
    CascadeMux I__1632 (
            .O(N__18653),
            .I(N__18650));
    InMux I__1631 (
            .O(N__18650),
            .I(N__18647));
    LocalMux I__1630 (
            .O(N__18647),
            .I(N__18644));
    Span4Mux_h I__1629 (
            .O(N__18644),
            .I(N__18641));
    Odrv4 I__1628 (
            .O(N__18641),
            .I(\pwm_generator_inst.un2_threshold_acc_1_22 ));
    InMux I__1627 (
            .O(N__18638),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ));
    InMux I__1626 (
            .O(N__18635),
            .I(N__18632));
    LocalMux I__1625 (
            .O(N__18632),
            .I(N__18629));
    Span4Mux_v I__1624 (
            .O(N__18629),
            .I(N__18626));
    Odrv4 I__1623 (
            .O(N__18626),
            .I(\pwm_generator_inst.un2_threshold_acc_2_8 ));
    CascadeMux I__1622 (
            .O(N__18623),
            .I(N__18620));
    InMux I__1621 (
            .O(N__18620),
            .I(N__18617));
    LocalMux I__1620 (
            .O(N__18617),
            .I(\pwm_generator_inst.un2_threshold_acc_1_23 ));
    InMux I__1619 (
            .O(N__18614),
            .I(bfn_1_11_0_));
    InMux I__1618 (
            .O(N__18611),
            .I(bfn_1_9_0_));
    InMux I__1617 (
            .O(N__18608),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ));
    InMux I__1616 (
            .O(N__18605),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ));
    InMux I__1615 (
            .O(N__18602),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ));
    InMux I__1614 (
            .O(N__18599),
            .I(N__18596));
    LocalMux I__1613 (
            .O(N__18596),
            .I(N__18593));
    Span4Mux_v I__1612 (
            .O(N__18593),
            .I(N__18590));
    Odrv4 I__1611 (
            .O(N__18590),
            .I(\pwm_generator_inst.un2_threshold_acc_2_0 ));
    CascadeMux I__1610 (
            .O(N__18587),
            .I(N__18584));
    InMux I__1609 (
            .O(N__18584),
            .I(N__18581));
    LocalMux I__1608 (
            .O(N__18581),
            .I(\pwm_generator_inst.un2_threshold_acc_1_15 ));
    InMux I__1607 (
            .O(N__18578),
            .I(N__18575));
    LocalMux I__1606 (
            .O(N__18575),
            .I(N__18572));
    Span4Mux_h I__1605 (
            .O(N__18572),
            .I(N__18569));
    Odrv4 I__1604 (
            .O(N__18569),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__1603 (
            .O(N__18566),
            .I(N__18563));
    LocalMux I__1602 (
            .O(N__18563),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ));
    InMux I__1601 (
            .O(N__18560),
            .I(N__18557));
    LocalMux I__1600 (
            .O(N__18557),
            .I(N__18554));
    Odrv4 I__1599 (
            .O(N__18554),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__1598 (
            .O(N__18551),
            .I(N__18548));
    LocalMux I__1597 (
            .O(N__18548),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ));
    InMux I__1596 (
            .O(N__18545),
            .I(N__18542));
    LocalMux I__1595 (
            .O(N__18542),
            .I(N__18539));
    Odrv4 I__1594 (
            .O(N__18539),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__1593 (
            .O(N__18536),
            .I(N__18533));
    LocalMux I__1592 (
            .O(N__18533),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ));
    InMux I__1591 (
            .O(N__18530),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ));
    InMux I__1590 (
            .O(N__18527),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ));
    InMux I__1589 (
            .O(N__18524),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ));
    InMux I__1588 (
            .O(N__18521),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ));
    InMux I__1587 (
            .O(N__18518),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ));
    InMux I__1586 (
            .O(N__18515),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ));
    InMux I__1585 (
            .O(N__18512),
            .I(N__18509));
    LocalMux I__1584 (
            .O(N__18509),
            .I(N__18506));
    Odrv4 I__1583 (
            .O(N__18506),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1582 (
            .O(N__18503),
            .I(N__18500));
    LocalMux I__1581 (
            .O(N__18500),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ));
    InMux I__1580 (
            .O(N__18497),
            .I(N__18494));
    LocalMux I__1579 (
            .O(N__18494),
            .I(N__18491));
    Odrv4 I__1578 (
            .O(N__18491),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1577 (
            .O(N__18488),
            .I(N__18485));
    LocalMux I__1576 (
            .O(N__18485),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ));
    InMux I__1575 (
            .O(N__18482),
            .I(N__18479));
    LocalMux I__1574 (
            .O(N__18479),
            .I(N__18476));
    Odrv4 I__1573 (
            .O(N__18476),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1572 (
            .O(N__18473),
            .I(N__18470));
    LocalMux I__1571 (
            .O(N__18470),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ));
    InMux I__1570 (
            .O(N__18467),
            .I(N__18464));
    LocalMux I__1569 (
            .O(N__18464),
            .I(N__18461));
    Odrv4 I__1568 (
            .O(N__18461),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1567 (
            .O(N__18458),
            .I(N__18455));
    LocalMux I__1566 (
            .O(N__18455),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ));
    InMux I__1565 (
            .O(N__18452),
            .I(N__18449));
    LocalMux I__1564 (
            .O(N__18449),
            .I(N__18446));
    Odrv4 I__1563 (
            .O(N__18446),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1562 (
            .O(N__18443),
            .I(N__18440));
    LocalMux I__1561 (
            .O(N__18440),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ));
    InMux I__1560 (
            .O(N__18437),
            .I(N__18434));
    LocalMux I__1559 (
            .O(N__18434),
            .I(N__18431));
    Odrv4 I__1558 (
            .O(N__18431),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1557 (
            .O(N__18428),
            .I(N__18425));
    LocalMux I__1556 (
            .O(N__18425),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ));
    InMux I__1555 (
            .O(N__18422),
            .I(N__18419));
    LocalMux I__1554 (
            .O(N__18419),
            .I(N__18416));
    Span4Mux_h I__1553 (
            .O(N__18416),
            .I(N__18413));
    Odrv4 I__1552 (
            .O(N__18413),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1551 (
            .O(N__18410),
            .I(N__18407));
    LocalMux I__1550 (
            .O(N__18407),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ));
    IoInMux I__1549 (
            .O(N__18404),
            .I(N__18401));
    LocalMux I__1548 (
            .O(N__18401),
            .I(N__18398));
    Span4Mux_s3_v I__1547 (
            .O(N__18398),
            .I(N__18395));
    Span4Mux_h I__1546 (
            .O(N__18395),
            .I(N__18392));
    Sp12to4 I__1545 (
            .O(N__18392),
            .I(N__18389));
    Span12Mux_s9_v I__1544 (
            .O(N__18389),
            .I(N__18386));
    Span12Mux_v I__1543 (
            .O(N__18386),
            .I(N__18383));
    Odrv12 I__1542 (
            .O(N__18383),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1541 (
            .O(N__18380),
            .I(N__18377));
    LocalMux I__1540 (
            .O(N__18377),
            .I(N__18374));
    IoSpan4Mux I__1539 (
            .O(N__18374),
            .I(N__18371));
    IoSpan4Mux I__1538 (
            .O(N__18371),
            .I(N__18368));
    Odrv4 I__1537 (
            .O(N__18368),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_13_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_10_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_24_0_));
    defparam IN_MUX_bfv_10_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_25_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_10_25_0_));
    defparam IN_MUX_bfv_10_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_26_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_10_26_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_16_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_16_18_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_16_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_20_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_16_20_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .carryinitout(bfn_1_8_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_3_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_8_0_));
    defparam IN_MUX_bfv_3_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_9_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .carryinitout(bfn_3_9_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un6_running_cry_8 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un6_running_cry_16 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un6_running_cry_8 ),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_10_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_23_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un6_running_cry_16 ),
            .carryinitout(bfn_10_23_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un6_running_cry_8 ),
            .carryinitout(bfn_15_12_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un6_running_cry_16 ),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un6_running_cry_8 ),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un6_running_cry_16 ),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_15_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_5_0_));
    defparam IN_MUX_bfv_15_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_6_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_15_6_0_));
    defparam IN_MUX_bfv_15_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_7_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_15_7_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_12_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_12_21_0_));
    defparam IN_MUX_bfv_12_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_12_22_0_));
    defparam IN_MUX_bfv_12_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_23_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_12_23_0_));
    defparam IN_MUX_bfv_13_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_21_0_));
    defparam IN_MUX_bfv_13_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_13_22_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_16_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_22_0_));
    defparam IN_MUX_bfv_16_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_23_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_16_23_0_));
    defparam IN_MUX_bfv_16_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_24_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_16_24_0_));
    defparam IN_MUX_bfv_16_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_25_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_16_25_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_7 ),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_7_16_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__18404),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__18380),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__32402),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_166_i_g ));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0  (
            .USERSIGNALTOGLOBALBUFFER(N__33677),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_434_i_g ));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__21743),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_432_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__37811),
            .CLKHFEN(N__37813),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__37812),
            .RGB2PWM(N__19052),
            .RGB1(rgb_g),
            .CURREN(N__37879),
            .RGB2(rgb_b),
            .RGB1PWM(N__19058),
            .RGB0PWM(N__45728),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21278),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46118),
            .ce(),
            .sr(N__45590));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_6_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_6_7  (
            .in0(N__19127),
            .in1(N__19138),
            .in2(_gnd_net_),
            .in3(N__20004),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__18503),
            .in2(_gnd_net_),
            .in3(N__18512),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1  (
            .in0(N__18497),
            .in1(N__18488),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2  (
            .in0(_gnd_net_),
            .in1(N__18473),
            .in2(_gnd_net_),
            .in3(N__18482),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3  (
            .in0(_gnd_net_),
            .in1(N__18458),
            .in2(_gnd_net_),
            .in3(N__18467),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4  (
            .in0(N__18452),
            .in1(N__18443),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(N__18428),
            .in2(_gnd_net_),
            .in3(N__18437),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6  (
            .in0(_gnd_net_),
            .in1(N__18410),
            .in2(_gnd_net_),
            .in3(N__18422),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7  (
            .in0(_gnd_net_),
            .in1(N__18566),
            .in2(_gnd_net_),
            .in3(N__18578),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(N__18551),
            .in2(_gnd_net_),
            .in3(N__18560),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ),
            .ltout(),
            .carryin(bfn_1_8_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1  (
            .in0(_gnd_net_),
            .in1(N__18536),
            .in2(_gnd_net_),
            .in3(N__18545),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(N__19024),
            .in2(_gnd_net_),
            .in3(N__18530),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3  (
            .in0(N__19726),
            .in1(N__19169),
            .in2(_gnd_net_),
            .in3(N__18527),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(N__19203),
            .in2(_gnd_net_),
            .in3(N__18524),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5  (
            .in0(_gnd_net_),
            .in1(N__19252),
            .in2(_gnd_net_),
            .in3(N__18521),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6  (
            .in0(_gnd_net_),
            .in1(N__19269),
            .in2(_gnd_net_),
            .in3(N__18518),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7  (
            .in0(_gnd_net_),
            .in1(N__18981),
            .in2(_gnd_net_),
            .in3(N__18515),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(N__19231),
            .in2(_gnd_net_),
            .in3(N__18611),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(N__19182),
            .in2(_gnd_net_),
            .in3(N__18608),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__19045),
            .in2(_gnd_net_),
            .in3(N__18605),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18602),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_1_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_1_9_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(N__19300),
            .in2(_gnd_net_),
            .in3(N__19046),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_1_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_1_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(N__19183),
            .in2(_gnd_net_),
            .in3(N__19327),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_1_9_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_1_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_1_9_6  (
            .in0(N__19369),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18983),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_9_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_9_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(N__19396),
            .in2(_gnd_net_),
            .in3(N__19271),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__18599),
            .in2(N__18587),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__18839),
            .in2(N__18827),
            .in3(N__18815),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_10_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__18812),
            .in2(N__18800),
            .in3(N__18788),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_10_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__18785),
            .in2(N__18773),
            .in3(N__18761),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_10_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__18758),
            .in2(N__18746),
            .in3(N__18728),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_10_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__18725),
            .in2(N__18713),
            .in3(N__18698),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_10_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(N__18695),
            .in2(N__18683),
            .in3(N__18668),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_10_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(N__18665),
            .in2(N__18653),
            .in3(N__18638),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__18635),
            .in2(N__18623),
            .in3(N__18614),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__18965),
            .in2(N__18953),
            .in3(N__18941),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__18938),
            .in2(N__19124),
            .in3(N__18926),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__19112),
            .in2(N__18923),
            .in3(N__18908),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__18905),
            .in2(N__19125),
            .in3(N__18893),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__19116),
            .in2(N__18890),
            .in3(N__18875),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__18872),
            .in2(N__19126),
            .in3(N__18860),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__19120),
            .in2(N__18857),
            .in3(N__18845),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_12_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_12_0  (
            .in0(N__19517),
            .in1(N__19064),
            .in2(_gnd_net_),
            .in3(N__18842),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_12_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_12_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_12_1  (
            .in0(N__19145),
            .in1(N__19105),
            .in2(N__20069),
            .in3(N__19076),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_13_0 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_13_0  (
            .in0(N__20667),
            .in1(N__21264),
            .in2(N__20813),
            .in3(N__20520),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46103),
            .ce(),
            .sr(N__45641));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_13_1 .LUT_INIT=16'b1101010111000100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_13_1  (
            .in0(N__21265),
            .in1(N__20759),
            .in2(N__20522),
            .in3(N__20668),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46103),
            .ce(),
            .sr(N__45641));
    defparam rgb_drv_RNO_LC_1_29_4.C_ON=1'b0;
    defparam rgb_drv_RNO_LC_1_29_4.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_LC_1_29_4.LUT_INIT=16'b0101010100000000;
    LogicCell40 rgb_drv_RNO_LC_1_29_4 (
            .in0(N__45726),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40576),
            .lcout(rgb_drv_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_0_LC_1_30_5.C_ON=1'b0;
    defparam rgb_drv_RNO_0_LC_1_30_5.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_0_LC_1_30_5.LUT_INIT=16'b1010101001010101;
    LogicCell40 rgb_drv_RNO_0_LC_1_30_5 (
            .in0(N__45727),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40580),
            .lcout(N_38_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_8_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_8_4 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_8_4  (
            .in0(N__19044),
            .in1(N__19304),
            .in2(N__19760),
            .in3(N__19031),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_8_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_8_5  (
            .in0(N__19025),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19012),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_8_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_8_6 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_8_6  (
            .in0(N__19013),
            .in1(N__18998),
            .in2(N__18992),
            .in3(N__19748),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_8_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_8_7 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_8_7  (
            .in0(N__19749),
            .in1(N__18989),
            .in2(N__19376),
            .in3(N__18982),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0  (
            .in0(N__19277),
            .in1(N__19270),
            .in2(N__19400),
            .in3(N__19719),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_1  (
            .in0(N__19253),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19423),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_2 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_2  (
            .in0(N__19424),
            .in1(N__19241),
            .in2(N__19235),
            .in3(N__19718),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_9_3  (
            .in0(N__19205),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19447),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__19345),
            .in2(_gnd_net_),
            .in3(N__19232),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_5 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_5  (
            .in0(N__19346),
            .in1(N__19220),
            .in2(N__19214),
            .in3(N__19754),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_6 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_6  (
            .in0(N__19211),
            .in1(N__19204),
            .in2(N__19451),
            .in3(N__19717),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_7 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_7  (
            .in0(N__19190),
            .in1(N__19184),
            .in2(N__19744),
            .in3(N__19328),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__19168),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__19463),
            .in2(_gnd_net_),
            .in3(N__19439),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_10_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(N__19436),
            .in2(_gnd_net_),
            .in3(N__19415),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_10_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__19412),
            .in2(_gnd_net_),
            .in3(N__19385),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_10_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__19382),
            .in2(_gnd_net_),
            .in3(N__19358),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_10_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_10_5  (
            .in0(_gnd_net_),
            .in1(N__37669),
            .in2(N__19355),
            .in3(N__19337),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_10_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(N__19334),
            .in2(N__37722),
            .in3(N__19316),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_10_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(N__37673),
            .in2(N__19313),
            .in3(N__19289),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__19286),
            .in2(_gnd_net_),
            .in3(N__19280),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__19511),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__19505),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__19499),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__19493),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__19487),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__19481),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__19475),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__19469),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__19538),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__19532),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__19526),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_12_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19520),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_2_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_2_14_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__21032),
            .in2(_gnd_net_),
            .in3(N__21053),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_5_LC_3_6_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_5_LC_3_6_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_5_LC_3_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_5_LC_3_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19640),
            .lcout(\pwm_generator_inst.thresholdZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46117),
            .ce(),
            .sr(N__45579));
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_7_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_7_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_7_1 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_2_LC_3_7_1  (
            .in0(N__20123),
            .in1(N__20064),
            .in2(N__19592),
            .in3(N__20270),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46115),
            .ce(),
            .sr(N__45584));
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_7_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_7_2 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_3_7_2 .LUT_INIT=16'b1111111101010011;
    LogicCell40 \pwm_generator_inst.threshold_ACC_6_LC_3_7_2  (
            .in0(N__20273),
            .in1(N__20126),
            .in2(N__20077),
            .in3(N__19805),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46115),
            .ce(),
            .sr(N__45584));
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_7_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_7_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_7_3 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_0_LC_3_7_3  (
            .in0(N__20121),
            .in1(N__20062),
            .in2(N__19628),
            .in3(N__20268),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46115),
            .ce(),
            .sr(N__45584));
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_7_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_7_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_7_5 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_3_LC_3_7_5  (
            .in0(N__20124),
            .in1(N__20065),
            .in2(N__19574),
            .in3(N__20271),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46115),
            .ce(),
            .sr(N__45584));
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_7_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_7_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_7_6 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_5_LC_3_7_6  (
            .in0(N__20272),
            .in1(N__20125),
            .in2(N__20076),
            .in3(N__19547),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46115),
            .ce(),
            .sr(N__45584));
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_7_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_7_7 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_7_7 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_1_LC_3_7_7  (
            .in0(N__20122),
            .in1(N__20063),
            .in2(N__19610),
            .in3(N__20269),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46115),
            .ce(),
            .sr(N__45584));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0  (
            .in0(_gnd_net_),
            .in1(N__19634),
            .in2(N__19759),
            .in3(N__19753),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_3_8_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1  (
            .in0(_gnd_net_),
            .in1(N__19619),
            .in2(_gnd_net_),
            .in3(N__19601),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2  (
            .in0(_gnd_net_),
            .in1(N__19598),
            .in2(_gnd_net_),
            .in3(N__19583),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3  (
            .in0(_gnd_net_),
            .in1(N__19580),
            .in2(_gnd_net_),
            .in3(N__19565),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4  (
            .in0(_gnd_net_),
            .in1(N__19562),
            .in2(_gnd_net_),
            .in3(N__19556),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5  (
            .in0(_gnd_net_),
            .in1(N__19553),
            .in2(_gnd_net_),
            .in3(N__19541),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6  (
            .in0(_gnd_net_),
            .in1(N__19811),
            .in2(_gnd_net_),
            .in3(N__19799),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7  (
            .in0(_gnd_net_),
            .in1(N__19796),
            .in2(_gnd_net_),
            .in3(N__19790),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0  (
            .in0(_gnd_net_),
            .in1(N__19787),
            .in2(_gnd_net_),
            .in3(N__19781),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_3_9_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1  (
            .in0(N__19778),
            .in1(N__19769),
            .in2(N__19758),
            .in3(N__19667),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_3_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_3_9_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_3_9_3  (
            .in0(N__19654),
            .in1(N__19882),
            .in2(_gnd_net_),
            .in3(N__19909),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_duty_inputlt3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_9_4 .LUT_INIT=16'b1010101011111011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_3_9_4  (
            .in0(N__19865),
            .in1(N__20349),
            .in2(N__19664),
            .in3(N__20329),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_3_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_3_9_7 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_3_9_7  (
            .in0(N__21277),
            .in1(N__20848),
            .in2(_gnd_net_),
            .in3(N__20196),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_3_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_3_10_1 .LUT_INIT=16'b0011000000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_3_10_1  (
            .in0(N__19921),
            .in1(N__20869),
            .in2(N__19853),
            .in3(N__20661),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_3_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_3_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_3_10_2 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_3_10_2  (
            .in0(N__19849),
            .in1(N__20579),
            .in2(N__19661),
            .in3(N__19821),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46109),
            .ce(),
            .sr(N__45602));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_3_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_3_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_3_10_5 .LUT_INIT=16'b1100111111001101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_3_10_5  (
            .in0(N__19922),
            .in1(N__20870),
            .in2(N__19855),
            .in3(N__20662),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46109),
            .ce(),
            .sr(N__45602));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_3_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_3_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_3_10_6 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_3_10_6  (
            .in0(N__19894),
            .in1(N__20558),
            .in2(N__19856),
            .in3(N__19823),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46109),
            .ce(),
            .sr(N__45602));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_3_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_3_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_3_10_7 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_3_10_7  (
            .in0(N__19822),
            .in1(N__20570),
            .in2(N__19854),
            .in3(N__19895),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46109),
            .ce(),
            .sr(N__45602));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_11_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_11_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_3_11_3  (
            .in0(_gnd_net_),
            .in1(N__20428),
            .in2(_gnd_net_),
            .in3(N__20296),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_11_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_11_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_11_4  (
            .in0(N__20373),
            .in1(N__20451),
            .in2(N__19868),
            .in3(N__20397),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_11_5 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_11_5  (
            .in0(N__21269),
            .in1(N__20227),
            .in2(N__20216),
            .in3(N__20495),
            .lcout(\current_shift_inst.PI_CTRL.N_153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_11_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_11_6  (
            .in0(N__20669),
            .in1(N__21270),
            .in2(_gnd_net_),
            .in3(N__20206),
            .lcout(\current_shift_inst.PI_CTRL.N_154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_3_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_3_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_3_12_1 .LUT_INIT=16'b0100010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_3_12_1  (
            .in0(N__20183),
            .in1(N__20849),
            .in2(N__20231),
            .in3(N__20506),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46099),
            .ce(),
            .sr(N__45624));
    defparam \pwm_generator_inst.threshold_7_LC_4_6_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_7_LC_4_6_6 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_7_LC_4_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_7_LC_4_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20147),
            .lcout(\pwm_generator_inst.thresholdZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46116),
            .ce(),
            .sr(N__45574));
    defparam \pwm_generator_inst.threshold_2_LC_4_6_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_2_LC_4_6_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_2_LC_4_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_2_LC_4_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20177),
            .lcout(\pwm_generator_inst.thresholdZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46116),
            .ce(),
            .sr(N__45574));
    defparam \pwm_generator_inst.threshold_8_LC_4_7_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_8_LC_4_7_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_8_LC_4_7_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pwm_generator_inst.threshold_8_LC_4_7_0  (
            .in0(N__20132),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.thresholdZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46113),
            .ce(),
            .sr(N__45580));
    defparam \pwm_generator_inst.threshold_3_LC_4_7_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_3_LC_4_7_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_3_LC_4_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_3_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20171),
            .lcout(\pwm_generator_inst.thresholdZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46113),
            .ce(),
            .sr(N__45580));
    defparam \pwm_generator_inst.threshold_ACC_4_LC_4_8_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_4_8_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_4_8_2 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_4_LC_4_8_2  (
            .in0(N__20117),
            .in1(N__20074),
            .in2(N__20165),
            .in3(N__20264),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46112),
            .ce(),
            .sr(N__45585));
    defparam \pwm_generator_inst.threshold_ACC_7_LC_4_8_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_4_8_4 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_4_8_4 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_7_LC_4_8_4  (
            .in0(N__20118),
            .in1(N__20075),
            .in2(N__20156),
            .in3(N__20265),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46112),
            .ce(),
            .sr(N__45585));
    defparam \pwm_generator_inst.threshold_ACC_8_LC_4_8_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_4_8_5 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_4_8_5 .LUT_INIT=16'b1111111101010011;
    LogicCell40 \pwm_generator_inst.threshold_ACC_8_LC_4_8_5  (
            .in0(N__20266),
            .in1(N__20119),
            .in2(N__20078),
            .in3(N__20138),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46112),
            .ce(),
            .sr(N__45585));
    defparam \pwm_generator_inst.threshold_ACC_9_LC_4_8_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_4_8_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_4_8_6 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_9_LC_4_8_6  (
            .in0(N__20120),
            .in1(N__20267),
            .in2(N__20087),
            .in3(N__20073),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46112),
            .ce(),
            .sr(N__45585));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_4_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_4_9_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(N__20704),
            .in2(_gnd_net_),
            .in3(N__20802),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_9_7 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_4_9_7  (
            .in0(N__20731),
            .in1(N__20752),
            .in2(N__19925),
            .in3(N__20779),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_4_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_4_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_4_10_0 .LUT_INIT=16'b1111010001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_4_10_0  (
            .in0(N__21271),
            .in1(N__20665),
            .in2(N__20783),
            .in3(N__20515),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46104),
            .ce(),
            .sr(N__45596));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_4_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_4_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_4_10_1 .LUT_INIT=16'b1111001100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_4_10_1  (
            .in0(N__20664),
            .in1(N__21273),
            .in2(N__20521),
            .in3(N__20705),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46104),
            .ce(),
            .sr(N__45596));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_4_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_4_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_4_10_2 .LUT_INIT=16'b1111010001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_4_10_2  (
            .in0(N__21272),
            .in1(N__20666),
            .in2(N__20732),
            .in3(N__20516),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46104),
            .ce(),
            .sr(N__45596));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_10_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_10_3  (
            .in0(N__20452),
            .in1(N__20432),
            .in2(N__20404),
            .in3(N__20374),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_10_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_10_4 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_10_4  (
            .in0(N__20350),
            .in1(N__20330),
            .in2(N__20303),
            .in3(N__20300),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_4_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_4_11_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(N__20697),
            .in2(_gnd_net_),
            .in3(N__20778),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_4_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_4_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_4_11_3  (
            .in0(N__20803),
            .in1(N__20751),
            .in2(N__20234),
            .in3(N__20727),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_4_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_4_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(N__20834),
            .in2(_gnd_net_),
            .in3(N__20863),
            .lcout(\current_shift_inst.PI_CTRL.N_155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_4_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_4_11_6 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_4_11_6  (
            .in0(N__21253),
            .in1(N__20835),
            .in2(N__20207),
            .in3(N__20663),
            .lcout(\current_shift_inst.PI_CTRL.N_149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_12_0  (
            .in0(N__21139),
            .in1(N__20615),
            .in2(N__21314),
            .in3(N__20546),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_12_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_12_2  (
            .in0(N__20987),
            .in1(N__20975),
            .in2(N__20888),
            .in3(N__21065),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(N__21121),
            .in2(_gnd_net_),
            .in3(N__21169),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(N__21202),
            .in2(_gnd_net_),
            .in3(N__21187),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_12_5  (
            .in0(N__20974),
            .in1(N__20986),
            .in2(N__20540),
            .in3(N__21025),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_12_6  (
            .in0(N__20938),
            .in1(N__20887),
            .in2(N__20921),
            .in3(N__21064),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_4_12_7  (
            .in0(N__20477),
            .in1(N__20537),
            .in2(N__20531),
            .in3(N__20528),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_13_0  (
            .in0(N__20962),
            .in1(N__21082),
            .in2(N__21104),
            .in3(N__21292),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_13_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_13_3  (
            .in0(N__21293),
            .in1(N__20963),
            .in2(N__20471),
            .in3(N__21313),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_13_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_13_4  (
            .in0(N__20678),
            .in1(N__20609),
            .in2(N__20672),
            .in3(N__21110),
            .lcout(\current_shift_inst.PI_CTRL.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_13_5  (
            .in0(N__20998),
            .in1(N__21010),
            .in2(N__21158),
            .in3(N__21046),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_13_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_13_6  (
            .in0(N__21011),
            .in1(N__20999),
            .in2(N__20945),
            .in3(N__20920),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_4_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_4_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_4_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_4_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23664),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21385),
            .ce(),
            .sr(N__45654));
    defparam \pwm_generator_inst.threshold_1_LC_5_6_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_1_LC_5_6_1 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_1_LC_5_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_1_LC_5_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20603),
            .lcout(\pwm_generator_inst.thresholdZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46114),
            .ce(),
            .sr(N__45568));
    defparam \pwm_generator_inst.threshold_0_LC_5_6_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_0_LC_5_6_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_0_LC_5_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_0_LC_5_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20591),
            .lcout(\pwm_generator_inst.thresholdZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46114),
            .ce(),
            .sr(N__45568));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__21416),
            .in2(N__24125),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .clk(N__46100),
            .ce(),
            .sr(N__45591));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__21407),
            .in2(N__26414),
            .in3(N__20561),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(N__46100),
            .ce(),
            .sr(N__45591));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__21584),
            .in2(N__24053),
            .in3(N__20549),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__46100),
            .ce(),
            .sr(N__45591));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__21791),
            .in2(N__23981),
            .in3(N__20852),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__46100),
            .ce(),
            .sr(N__45591));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__21575),
            .in2(N__22907),
            .in3(N__20816),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__46100),
            .ce(),
            .sr(N__45591));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(N__21566),
            .in2(N__26153),
            .in3(N__20786),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__46100),
            .ce(),
            .sr(N__45591));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(N__21539),
            .in2(N__27530),
            .in3(N__20762),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__46100),
            .ce(),
            .sr(N__45591));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(N__21593),
            .in2(N__22319),
            .in3(N__20735),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__46100),
            .ce(),
            .sr(N__45591));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__23882),
            .in2(N__21398),
            .in3(N__20708),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__46095),
            .ce(),
            .sr(N__45597));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__21425),
            .in2(N__24194),
            .in3(N__20684),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__46095),
            .ce(),
            .sr(N__45597));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__21548),
            .in2(N__26942),
            .in3(N__20681),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__46095),
            .ce(),
            .sr(N__45597));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__21557),
            .in2(N__22661),
            .in3(N__20951),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__46095),
            .ce(),
            .sr(N__45597));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__21447),
            .in2(N__22505),
            .in3(N__20948),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__46095),
            .ce(),
            .sr(N__45597));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(N__22742),
            .in2(N__21489),
            .in3(N__20924),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__46095),
            .ce(),
            .sr(N__45597));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__21451),
            .in2(N__26342),
            .in3(N__20903),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__46095),
            .ce(),
            .sr(N__45597));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__23144),
            .in2(N__21490),
            .in3(N__20900),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__46095),
            .ce(),
            .sr(N__45597));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(N__21491),
            .in2(N__23294),
            .in3(N__20897),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__46089),
            .ce(),
            .sr(N__45603));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__23234),
            .in2(N__21521),
            .in3(N__20894),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__46089),
            .ce(),
            .sr(N__45603));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__21495),
            .in2(N__22994),
            .in3(N__20891),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__46089),
            .ce(),
            .sr(N__45603));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__26288),
            .in2(N__21522),
            .in3(N__20873),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__46089),
            .ce(),
            .sr(N__45603));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__21499),
            .in2(N__26819),
            .in3(N__21056),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__46089),
            .ce(),
            .sr(N__45603));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(N__26563),
            .in2(N__21523),
            .in3(N__21035),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__46089),
            .ce(),
            .sr(N__45603));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__21503),
            .in2(N__26687),
            .in3(N__21014),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__46089),
            .ce(),
            .sr(N__45603));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__24882),
            .in2(N__21524),
            .in3(N__21002),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__46089),
            .ce(),
            .sr(N__45603));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__21507),
            .in2(N__23522),
            .in3(N__20990),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__46080),
            .ce(),
            .sr(N__45611));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__23428),
            .in2(N__21525),
            .in3(N__20978),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__46080),
            .ce(),
            .sr(N__45611));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(N__21511),
            .in2(N__23374),
            .in3(N__20966),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__46080),
            .ce(),
            .sr(N__45611));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(N__31408),
            .in2(N__21526),
            .in3(N__20954),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__46080),
            .ce(),
            .sr(N__45611));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__21515),
            .in2(N__31352),
            .in3(N__21299),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__46080),
            .ce(),
            .sr(N__45611));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(N__27464),
            .in2(N__21527),
            .in3(N__21296),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__46080),
            .ce(),
            .sr(N__45611));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(N__21519),
            .in2(N__31463),
            .in3(N__21284),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__46080),
            .ce(),
            .sr(N__45611));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_13_7  (
            .in0(N__21520),
            .in1(N__27404),
            .in2(_gnd_net_),
            .in3(N__21281),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46080),
            .ce(),
            .sr(N__45611));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_5_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_5_14_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_5_14_2  (
            .in0(N__21206),
            .in1(N__21191),
            .in2(N__21176),
            .in3(N__21157),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_5_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_5_14_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_5_14_3  (
            .in0(N__21143),
            .in1(N__21071),
            .in2(N__21128),
            .in3(N__21125),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_5_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_5_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24049),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_5_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_5_14_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(N__21100),
            .in2(_gnd_net_),
            .in3(N__21086),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_5_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_5_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_5_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36917),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46068),
            .ce(),
            .sr(N__45633));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_5_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_5_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_5_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21913),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46068),
            .ce(),
            .sr(N__45633));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21893),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46068),
            .ce(),
            .sr(N__45633));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_5_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_5_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_5_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_5_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22861),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46068),
            .ce(),
            .sr(N__45633));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_5_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_5_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_5_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31610),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46042),
            .ce(N__33768),
            .sr(N__45652));
    defparam \delay_measurement_inst.stop_timer_hc_LC_5_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_5_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_5_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_5_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23665),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21386),
            .ce(),
            .sr(N__45655));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_1.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_1.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21374),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_6_LC_7_6_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_6_LC_7_6_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_6_LC_7_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_6_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21347),
            .lcout(\pwm_generator_inst.thresholdZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46110),
            .ce(),
            .sr(N__45561));
    defparam \pwm_generator_inst.threshold_4_LC_7_7_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_4_LC_7_7_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_4_LC_7_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_4_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21335),
            .lcout(\pwm_generator_inst.thresholdZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46105),
            .ce(),
            .sr(N__45565));
    defparam \pwm_generator_inst.threshold_9_LC_7_8_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_9_LC_7_8_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_9_LC_7_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_9_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21323),
            .lcout(\pwm_generator_inst.thresholdZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46101),
            .ce(),
            .sr(N__45569));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_7_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_7_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_7_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26462),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46090),
            .ce(),
            .sr(N__45581));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21872),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46090),
            .ce(),
            .sr(N__45581));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26758),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46090),
            .ce(),
            .sr(N__45581));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_7_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_7_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_7_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22816),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46090),
            .ce(),
            .sr(N__45581));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_11_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__21815),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46081),
            .ce(),
            .sr(N__45586));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_7_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_7_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_7_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27587),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46081),
            .ce(),
            .sr(N__45586));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22444),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46081),
            .ce(),
            .sr(N__45586));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33047),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46081),
            .ce(),
            .sr(N__45586));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26212),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46081),
            .ce(),
            .sr(N__45586));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_7_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_7_12_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMMAM_28_LC_7_12_1  (
            .in0(N__23417),
            .in1(N__31391),
            .in2(N__31345),
            .in3(N__23361),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_7_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_7_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGC4P2_19_LC_7_12_2  (
            .in0(N__21605),
            .in1(N__22589),
            .in2(N__21608),
            .in3(N__21758),
            .lcout(\current_shift_inst.PI_CTRL.N_74_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_7_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_7_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIBA9M_19_LC_7_12_3  (
            .in0(N__26679),
            .in1(N__23511),
            .in2(N__26564),
            .in3(N__26283),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_7_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_7_12_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIBB5B_28_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__31338),
            .in2(_gnd_net_),
            .in3(N__23416),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_7_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_7_12_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI01LC1_30_LC_7_12_5  (
            .in0(N__31459),
            .in1(N__31390),
            .in2(N__21599),
            .in3(N__21614),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_12_6 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_12_6  (
            .in0(N__26149),
            .in1(N__22906),
            .in2(N__23980),
            .in3(N__22277),
            .lcout(\current_shift_inst.PI_CTRL.N_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23138),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_7_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_7_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDA7M_15_LC_7_13_0  (
            .in0(N__22975),
            .in1(N__23223),
            .in2(N__23139),
            .in3(N__26811),
            .lcout(\current_shift_inst.PI_CTRL.N_74_16 ),
            .ltout(\current_shift_inst.PI_CTRL.N_74_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_7_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_7_13_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_11_LC_7_13_1  (
            .in0(N__21625),
            .in1(N__21634),
            .in2(N__21596),
            .in3(N__22649),
            .lcout(\current_shift_inst.PI_CTRL.N_103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_7_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_7_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26138),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_7_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_7_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36899),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_7_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_7_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23501),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_7_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_7_13_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDAC11_11_LC_7_13_5  (
            .in0(N__27395),
            .in1(N__21641),
            .in2(_gnd_net_),
            .in3(N__22648),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_7_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_7_13_6 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIE7HME_11_LC_7_13_6  (
            .in0(N__21635),
            .in1(N__21626),
            .in2(N__21617),
            .in3(N__21770),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_7_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_7_13_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFE9M_19_LC_7_13_7  (
            .in0(N__23500),
            .in1(N__26273),
            .in2(N__26559),
            .in3(N__23347),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_7_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_7_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_7_14_1 .LUT_INIT=16'b0100111101000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_7_14_1  (
            .in0(N__27193),
            .in1(N__27398),
            .in2(N__24209),
            .in3(N__27035),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46062),
            .ce(),
            .sr(N__45604));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_7_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_7_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22638),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_14_4 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_7_14_4  (
            .in0(N__27396),
            .in1(N__27196),
            .in2(N__27090),
            .in3(N__24776),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46062),
            .ce(),
            .sr(N__45604));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_7_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_7_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_7_14_5 .LUT_INIT=16'b0100111101000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_7_14_5  (
            .in0(N__27194),
            .in1(N__27399),
            .in2(N__24737),
            .in3(N__27036),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46062),
            .ce(),
            .sr(N__45604));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_7_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_7_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_7_14_6 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_7_14_6  (
            .in0(N__27397),
            .in1(N__27197),
            .in2(N__27091),
            .in3(N__24698),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46062),
            .ce(),
            .sr(N__45604));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_7_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_7_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_7_14_7 .LUT_INIT=16'b0100111101000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_7_14_7  (
            .in0(N__27195),
            .in1(N__27400),
            .in2(N__24659),
            .in3(N__27037),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46062),
            .ce(),
            .sr(N__45604));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__21674),
            .in2(_gnd_net_),
            .in3(N__36916),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_7_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_7_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_7_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__21668),
            .in2(_gnd_net_),
            .in3(N__21659),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__46054),
            .ce(),
            .sr(N__45612));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_7_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_7_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_7_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__26228),
            .in2(_gnd_net_),
            .in3(N__21656),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__46054),
            .ce(),
            .sr(N__45612));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_7_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_7_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_7_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__26720),
            .in2(_gnd_net_),
            .in3(N__21653),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__46054),
            .ce(),
            .sr(N__45612));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_7_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_7_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_7_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__22073),
            .in2(_gnd_net_),
            .in3(N__21650),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__46054),
            .ce(),
            .sr(N__45612));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_7_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_7_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_7_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(N__23162),
            .in2(_gnd_net_),
            .in3(N__21647),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__46054),
            .ce(),
            .sr(N__45612));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_7_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_7_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_7_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(N__26828),
            .in2(_gnd_net_),
            .in3(N__21644),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__46054),
            .ce(),
            .sr(N__45612));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_7_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_7_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_7_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(N__21824),
            .in2(_gnd_net_),
            .in3(N__21692),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__46054),
            .ce(),
            .sr(N__45612));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_7_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_7_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_7_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__33158),
            .in2(_gnd_net_),
            .in3(N__21689),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__46048),
            .ce(),
            .sr(N__45625));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_7_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_7_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_7_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__47387),
            .in2(_gnd_net_),
            .in3(N__21686),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__46048),
            .ce(),
            .sr(N__45625));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_7_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_7_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_7_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(N__31628),
            .in2(_gnd_net_),
            .in3(N__21683),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__46048),
            .ce(),
            .sr(N__45625));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_7_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_7_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_7_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__36998),
            .in2(_gnd_net_),
            .in3(N__21680),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__46048),
            .ce(),
            .sr(N__45625));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_7_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_7_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_7_16_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(N__37037),
            .in2(_gnd_net_),
            .in3(N__21677),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46048),
            .ce(),
            .sr(N__45625));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_7_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_7_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22845),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_7_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_7_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26202),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_7_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_7_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27579),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_7_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_7_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__22525),
            .in2(_gnd_net_),
            .in3(N__32943),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_7_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_7_17_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_7_17_1  (
            .in0(N__32948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22939),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_7_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_7_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_7_17_2  (
            .in0(N__23092),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32946),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_7_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_7_17_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_7_17_3  (
            .in0(N__32944),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22705),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_7_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_7_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_7_17_4  (
            .in0(N__23479),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32950),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_7_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_7_17_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_7_17_5  (
            .in0(N__32945),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22558),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_7_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_7_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_7_17_6  (
            .in0(N__24826),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32949),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_7_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_7_17_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_7_17_7  (
            .in0(N__32947),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23314),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_7_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_7_18_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_7_18_2  (
            .in0(N__23813),
            .in1(N__23599),
            .in2(N__28494),
            .in3(N__22046),
            .lcout(\phase_controller_inst1.stoper_hc.N_337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_7_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_7_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_7_18_6 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_7_18_6  (
            .in0(N__28242),
            .in1(N__23576),
            .in2(N__27878),
            .in3(N__23600),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46036),
            .ce(N__28873),
            .sr(N__45637));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_7_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_7_19_1 .LUT_INIT=16'b1111110011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5LMJQ_9_LC_7_19_1  (
            .in0(N__23605),
            .in1(N__30202),
            .in2(N__30485),
            .in3(N__41565),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_7_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_7_19_3 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILKVDQ_18_LC_7_19_3  (
            .in0(N__23769),
            .in1(N__41567),
            .in2(N__30701),
            .in3(N__30204),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_7_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_7_19_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI51CED1_18_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21746),
            .in3(N__30270),
            .lcout(elapsed_time_ns_1_RNI51CED1_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_7_19_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_7_19_7 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHGVDQ_14_LC_7_19_7  (
            .in0(N__23827),
            .in1(N__41566),
            .in2(N__30347),
            .in3(N__30203),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_7_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_7_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_7_20_4  (
            .in0(N__23031),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33046),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_7_22_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_7_22_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_7_22_2 .LUT_INIT=16'b1111111111100100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMLVDQ_19_LC_7_22_2  (
            .in0(N__41569),
            .in1(N__23712),
            .in2(N__30665),
            .in3(N__30206),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_25_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_25_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_25_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_25_4  (
            .in0(_gnd_net_),
            .in1(N__28685),
            .in2(_gnd_net_),
            .in3(N__23640),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_432_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_0.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_8_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21728),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46111),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_8_6_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_8_6_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_8_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_8_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21719),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46106),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_9_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_9_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_9_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_8_9_4 (
            .in0(N__21704),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46091),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_8_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_8_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_8_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21851),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46082),
            .ce(),
            .sr(N__45575));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_8_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_8_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21814),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_8_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_8_12_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID9B11_22_LC_8_12_0  (
            .in0(N__22650),
            .in1(N__26680),
            .in2(_gnd_net_),
            .in3(N__21752),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_8_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_8_12_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_12_LC_8_12_1  (
            .in0(N__22397),
            .in1(N__22403),
            .in2(N__21782),
            .in3(N__21779),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_8_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_8_12_2 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIC35V7_4_LC_8_12_2  (
            .in0(N__21764),
            .in1(N__22895),
            .in2(N__21773),
            .in3(N__22409),
            .lcout(\current_shift_inst.PI_CTRL.N_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_8_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_8_12_3 .LUT_INIT=16'b0000000111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIQB1L1_0_LC_8_12_3  (
            .in0(N__24048),
            .in1(N__26410),
            .in2(N__24124),
            .in3(N__23973),
            .lcout(\current_shift_inst.PI_CTRL.N_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_8_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_8_12_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_8_12_4  (
            .in0(N__23360),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_8_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_8_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_29_LC_8_12_6  (
            .in0(N__24881),
            .in1(N__27459),
            .in2(N__23289),
            .in3(N__26937),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_8_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_8_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_8_12_7  (
            .in0(N__22770),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33048),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_8_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_8_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDA7M_0_15_LC_8_13_0  (
            .in0(N__26803),
            .in1(N__23221),
            .in2(N__22985),
            .in3(N__23128),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_8_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_8_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22440),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37097),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_8_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_8_13_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_8_13_3  (
            .in0(N__33084),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26637),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_8_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_8_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23266),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_8_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_8_13_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__23959),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_8_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_8_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24111),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_8_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_8_14_0 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIGQQ01_11_LC_8_14_0  (
            .in0(N__22298),
            .in1(N__21813),
            .in2(N__33131),
            .in3(N__21932),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIGQQ01Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22297),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_14_2 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_8_14_2  (
            .in0(N__27200),
            .in1(N__27391),
            .in2(N__27094),
            .in3(N__24320),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46055),
            .ce(),
            .sr(N__45598));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_8_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_8_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_8_14_3 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_8_14_3  (
            .in0(N__27387),
            .in1(N__27201),
            .in2(N__24515),
            .in3(N__27047),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46055),
            .ce(),
            .sr(N__45598));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_8_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_8_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_8_14_4 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_8_14_4  (
            .in0(N__27198),
            .in1(N__27389),
            .in2(N__27092),
            .in3(N__24470),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46055),
            .ce(),
            .sr(N__45598));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_14_5 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_8_14_5  (
            .in0(N__27388),
            .in1(N__27202),
            .in2(N__24440),
            .in3(N__27048),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46055),
            .ce(),
            .sr(N__45598));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_14_6 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_8_14_6  (
            .in0(N__27199),
            .in1(N__27390),
            .in2(N__27093),
            .in3(N__24398),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46055),
            .ce(),
            .sr(N__45598));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_8_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_8_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__21899),
            .in2(_gnd_net_),
            .in3(N__21914),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_8_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_8_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__21878),
            .in2(_gnd_net_),
            .in3(N__21889),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_8_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_8_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__21857),
            .in2(_gnd_net_),
            .in3(N__21868),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_8_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_8_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__21833),
            .in2(_gnd_net_),
            .in3(N__21844),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_8_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_8_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__26729),
            .in2(_gnd_net_),
            .in3(N__21827),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_8_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_8_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__22787),
            .in2(_gnd_net_),
            .in3(N__21986),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_8_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_8_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__21983),
            .in2(_gnd_net_),
            .in3(N__21974),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_8_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_8_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(N__26426),
            .in2(_gnd_net_),
            .in3(N__21971),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_8_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_8_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__21968),
            .in2(_gnd_net_),
            .in3(N__21962),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_8 ),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_8_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_8_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(N__21959),
            .in2(_gnd_net_),
            .in3(N__21953),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_8_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_8_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_8_16_2  (
            .in0(_gnd_net_),
            .in1(N__21950),
            .in2(_gnd_net_),
            .in3(N__21944),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_8_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_8_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_8_16_3  (
            .in0(_gnd_net_),
            .in1(N__21941),
            .in2(_gnd_net_),
            .in3(N__21923),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_8_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_8_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_LUT4_0_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(N__23061),
            .in2(_gnd_net_),
            .in3(N__21920),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_8_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_8_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_LUT4_0_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(N__23010),
            .in2(_gnd_net_),
            .in3(N__21917),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_8_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_8_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_8_16_6  (
            .in0(_gnd_net_),
            .in1(N__22771),
            .in2(_gnd_net_),
            .in3(N__22013),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_8_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_8_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_8_16_7  (
            .in0(_gnd_net_),
            .in1(N__22672),
            .in2(_gnd_net_),
            .in3(N__22010),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_8_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_8_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__22521),
            .in2(_gnd_net_),
            .in3(N__22007),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_8_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_8_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(N__22695),
            .in2(_gnd_net_),
            .in3(N__22004),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_8_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_8_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_8_17_2  (
            .in0(_gnd_net_),
            .in1(N__22554),
            .in2(_gnd_net_),
            .in3(N__22001),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_8_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_8_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(N__23088),
            .in2(_gnd_net_),
            .in3(N__21998),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_8_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_8_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_8_17_4  (
            .in0(_gnd_net_),
            .in1(N__23310),
            .in2(_gnd_net_),
            .in3(N__21995),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_8_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_8_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(N__23194),
            .in2(_gnd_net_),
            .in3(N__21992),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_8_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_8_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__22935),
            .in2(_gnd_net_),
            .in3(N__21989),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_8_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_8_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(N__26710),
            .in2(_gnd_net_),
            .in3(N__22040),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_8_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_8_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__23032),
            .in2(_gnd_net_),
            .in3(N__22037),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_8_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_8_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__26593),
            .in2(_gnd_net_),
            .in3(N__22034),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_8_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_8_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__26638),
            .in2(_gnd_net_),
            .in3(N__22031),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_8_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_8_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__24822),
            .in2(_gnd_net_),
            .in3(N__22028),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_8_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_8_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__23475),
            .in2(_gnd_net_),
            .in3(N__22025),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_8_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_8_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(N__23452),
            .in2(_gnd_net_),
            .in3(N__22022),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_8_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_8_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_8_18_6  (
            .in0(_gnd_net_),
            .in1(N__23386),
            .in2(_gnd_net_),
            .in3(N__22019),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_8_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_8_18_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54K_LC_8_18_7  (
            .in0(N__33111),
            .in1(N__31409),
            .in2(_gnd_net_),
            .in3(N__22016),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNIG54KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_8_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_8_19_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL13KD1_9_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__22079),
            .in2(_gnd_net_),
            .in3(N__30265),
            .lcout(elapsed_time_ns_1_RNIL13KD1_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37148),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_8_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_8_19_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1TBED1_14_LC_8_19_2  (
            .in0(N__22061),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30266),
            .lcout(elapsed_time_ns_1_RNI1TBED1_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_8_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_8_19_3 .LUT_INIT=16'b1111110111101100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJIVDQ_16_LC_8_19_3  (
            .in0(N__41545),
            .in1(N__30200),
            .in2(N__30767),
            .in3(N__23549),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_8_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_8_19_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3VBED1_16_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22055),
            .in3(N__30264),
            .lcout(elapsed_time_ns_1_RNI3VBED1_0_16),
            .ltout(elapsed_time_ns_1_RNI3VBED1_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_8_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_8_19_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_8_19_5  (
            .in0(N__28339),
            .in1(N__23732),
            .in2(N__22052),
            .in3(N__28086),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_8_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_8_19_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(N__23708),
            .in2(N__22049),
            .in3(N__23762),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_8_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_8_19_7 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_8_19_7  (
            .in0(N__23763),
            .in1(N__23550),
            .in2(N__23714),
            .in3(N__23742),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_8_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_8_20_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI40CED1_17_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(N__22130),
            .in2(_gnd_net_),
            .in3(N__30263),
            .lcout(elapsed_time_ns_1_RNI40CED1_0_17),
            .ltout(elapsed_time_ns_1_RNI40CED1_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_8_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_8_20_1 .LUT_INIT=16'b1111111010111010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKJVDQ_17_LC_8_20_1  (
            .in0(N__30205),
            .in1(N__41568),
            .in2(N__22133),
            .in3(N__30731),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_14_LC_8_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_14_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_14_LC_8_20_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_14_LC_8_20_2  (
            .in0(_gnd_net_),
            .in1(N__28481),
            .in2(_gnd_net_),
            .in3(N__27752),
            .lcout(\phase_controller_inst1.stoper_hc.N_287 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_8_20_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_8_20_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3PJ05_15_LC_8_20_3  (
            .in0(N__45723),
            .in1(N__27992),
            .in2(N__28564),
            .in3(N__29900),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_a3_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_8_20_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_8_20_4 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9_24_LC_8_20_4  (
            .in0(N__28603),
            .in1(_gnd_net_),
            .in2(N__22124),
            .in3(N__29930),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBF1F9Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_8_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_8_20_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719_21_LC_8_20_5  (
            .in0(N__45722),
            .in1(N__28604),
            .in2(N__28565),
            .in3(N__29876),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI05719Z0Z_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_8_20_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_8_20_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGCC0J_31_LC_8_20_6  (
            .in0(N__45724),
            .in1(N__30850),
            .in2(N__22121),
            .in3(N__22118),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_8_20_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_8_20_7 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62CED1_19_LC_8_20_7  (
            .in0(N__22112),
            .in1(_gnd_net_),
            .in2(N__22103),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNI62CED1_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_8_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_8_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_8_21_3 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_8_21_3  (
            .in0(N__28489),
            .in1(N__23828),
            .in2(_gnd_net_),
            .in3(N__27751),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_8_25_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_8_25_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_8_25_2 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_8_25_2  (
            .in0(N__28690),
            .in1(N__23678),
            .in2(_gnd_net_),
            .in3(N__23644),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46008),
            .ce(),
            .sr(N__45657));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_6_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__22100),
            .in2(N__22091),
            .in3(N__25682),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_6_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__22268),
            .in2(N__22259),
            .in3(N__26075),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_6_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__22250),
            .in2(N__22241),
            .in3(N__26048),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_6_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(N__22232),
            .in2(N__22217),
            .in3(N__26024),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_6_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_6_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_6_4  (
            .in0(N__25997),
            .in1(N__22208),
            .in2(N__22196),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_6_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_6_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_6_5  (
            .in0(N__25973),
            .in1(N__22187),
            .in2(N__22178),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_6_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__22157),
            .in2(N__22169),
            .in3(N__25949),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_6_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(N__22139),
            .in2(N__22151),
            .in3(N__25922),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_7_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__22391),
            .in2(N__22382),
            .in3(N__25898),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_7_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__22373),
            .in2(N__22361),
            .in3(N__25832),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_9_7_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_9_7_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_9_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22352),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46096),
            .ce(),
            .sr(N__45557));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_10_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_10_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_9_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22328),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46074),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_9_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_9_11_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__22308),
            .in2(_gnd_net_),
            .in3(N__26142),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_9_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_9_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23427),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22990),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_9_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_9_12_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_9_12_1  (
            .in0(N__22318),
            .in1(N__23867),
            .in2(N__27528),
            .in3(N__24179),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_9_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_9_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22731),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_9_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_9_12_3 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_9_12_3  (
            .in0(N__22415),
            .in1(N__23868),
            .in2(N__27529),
            .in3(N__24180),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_9_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_9_12_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_29_LC_9_12_4  (
            .in0(N__24880),
            .in1(N__23279),
            .in2(N__26938),
            .in3(N__27458),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_9_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_9_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22486),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_9_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_9_12_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_9_12_6  (
            .in0(N__33050),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26586),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_9_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_9_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_9_12_7  (
            .in0(N__23187),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33049),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22888),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_9_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_9_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_9_13_2 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_9_13_2  (
            .in0(N__27378),
            .in1(N__27224),
            .in2(N__27114),
            .in3(N__24371),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46056),
            .ce(),
            .sr(N__45587));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_9_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_9_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_9_13_3 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_9_13_3  (
            .in0(N__27221),
            .in1(N__27379),
            .in2(N__27115),
            .in3(N__24593),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46056),
            .ce(),
            .sr(N__45587));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_13_4 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_9_13_4  (
            .in0(N__27376),
            .in1(N__27222),
            .in2(N__27112),
            .in3(N__24566),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46056),
            .ce(),
            .sr(N__45587));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_9_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_9_13_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI428M_12_LC_9_13_5  (
            .in0(N__26327),
            .in1(N__22729),
            .in2(N__22498),
            .in3(N__27375),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_9_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_9_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_9_13_6 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_9_13_6  (
            .in0(N__27377),
            .in1(N__27223),
            .in2(N__27113),
            .in3(N__24548),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46056),
            .ce(),
            .sr(N__45587));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_9_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_9_13_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI318M_30_LC_9_13_7  (
            .in0(N__26326),
            .in1(N__22730),
            .in2(N__22497),
            .in3(N__31455),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_9_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_9_14_0 .LUT_INIT=16'b1010000010101111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIVJ2U_4_LC_9_14_0  (
            .in0(N__22577),
            .in1(N__24148),
            .in2(N__33128),
            .in3(N__26759),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIVJ2UZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_9_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_9_14_1 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI3P3U_5_LC_9_14_1  (
            .in0(N__22571),
            .in1(N__26400),
            .in2(N__22820),
            .in3(N__33088),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI3P3UZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_9_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_9_14_2 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84I_LC_9_14_2  (
            .in0(N__22565),
            .in1(N__26331),
            .in2(N__33130),
            .in3(N__22538),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIH84IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_9_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_9_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23222),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_9_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_9_14_4 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22I_LC_9_14_4  (
            .in0(N__22529),
            .in1(N__22496),
            .in2(N__33129),
            .in3(N__22463),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNID22IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_9_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_9_14_5 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI7U4U_6_LC_9_14_5  (
            .in0(N__24038),
            .in1(N__22454),
            .in2(N__22448),
            .in3(N__33089),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI7U4UZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_9_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_9_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27460),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_9_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_9_14_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIF87U_8_LC_9_14_7  (
            .in0(N__22896),
            .in1(N__33090),
            .in2(N__22862),
            .in3(N__22829),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIF87UZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_9_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_9_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22812),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_9_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_9_15_1 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MP_LC_9_15_1  (
            .in0(N__24190),
            .in1(N__23011),
            .in2(N__33126),
            .in3(N__22781),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNI00MPZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_9_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_9_15_2 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVH_LC_9_15_2  (
            .in0(N__26930),
            .in1(N__33076),
            .in2(N__22775),
            .in3(N__22748),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNI9SVHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_9_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_9_15_3 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53I_LC_9_15_3  (
            .in0(N__22741),
            .in1(N__22706),
            .in2(N__33127),
            .in3(N__22682),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIF53IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_9_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_9_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__22673),
            .in2(_gnd_net_),
            .in3(N__33073),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_9_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_9_15_5 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0I_LC_9_15_5  (
            .in0(N__33080),
            .in1(N__22660),
            .in2(N__22616),
            .in3(N__22613),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIBV0IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_9_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_9_15_6 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIB36U_7_LC_9_15_6  (
            .in0(N__26461),
            .in1(N__23969),
            .in2(N__22607),
            .in3(N__33074),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIB36UZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_9_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_9_15_7 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKP_LC_9_15_7  (
            .in0(N__33075),
            .in1(N__23878),
            .in2(N__23066),
            .in3(N__22595),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNIUSKPZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_9_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_9_16_0 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00J_LC_9_16_0  (
            .in0(N__23233),
            .in1(N__23195),
            .in2(N__33066),
            .in3(N__23171),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIE00JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37127),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_9_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_9_16_2 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62J_LC_9_16_2  (
            .in0(N__26287),
            .in1(N__26711),
            .in2(N__33067),
            .in3(N__23150),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNII62JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_9_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_9_16_3 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5I_LC_9_16_3  (
            .in0(N__23143),
            .in1(N__32978),
            .in2(N__23099),
            .in3(N__23072),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIJB5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_9_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_9_16_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_inv_LC_9_16_4  (
            .in0(N__32974),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23065),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_9_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_9_16_5 .LUT_INIT=16'b0110111101101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14J_LC_9_16_5  (
            .in0(N__23045),
            .in1(N__23036),
            .in2(N__33132),
            .in3(N__26815),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIB14JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_9_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_9_16_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_inv_LC_9_16_6  (
            .in0(N__23012),
            .in1(_gnd_net_),
            .in2(N__33065),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_9_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_9_16_7 .LUT_INIT=16'b0011110011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31J_LC_9_16_7  (
            .in0(N__22989),
            .in1(N__22943),
            .in2(N__22919),
            .in3(N__32982),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIG31JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_9_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_9_17_0 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8J_LC_9_17_0  (
            .in0(N__23521),
            .in1(N__23480),
            .in2(N__33133),
            .in3(N__23459),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIJD8JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_9_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_9_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_9_17_1  (
            .in0(N__23453),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33103),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_9_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_9_17_2 .LUT_INIT=16'b0111110101111101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9J_LC_9_17_2  (
            .in0(N__33110),
            .in1(N__23441),
            .in2(N__23432),
            .in3(N__23429),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNILG9JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_9_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_9_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_9_17_3  (
            .in0(N__23387),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33104),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_9_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_9_17_4 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJ_LC_9_17_4  (
            .in0(N__33109),
            .in1(N__23375),
            .in2(N__23324),
            .in3(N__23321),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNINJAJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.N_266_i_1_LC_9_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.N_266_i_1_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.N_266_i_1_LC_9_17_5 .LUT_INIT=16'b0101000101010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.N_266_i_1_LC_9_17_5  (
            .in0(N__27753),
            .in1(N__24977),
            .in2(N__28496),
            .in3(N__23829),
            .lcout(\phase_controller_inst1.stoper_hc.N_266_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_9_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_9_17_7 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6I_LC_9_17_7  (
            .in0(N__23315),
            .in1(N__23290),
            .in2(N__23246),
            .in3(N__33105),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNILE6IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_9_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_9_18_2 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_9_18_2  (
            .in0(N__23814),
            .in1(N__23601),
            .in2(_gnd_net_),
            .in3(N__24975),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.N_275_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_9_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_9_18_3 .LUT_INIT=16'b0011001100010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_9_18_3  (
            .in0(N__28485),
            .in1(N__27810),
            .in2(N__23237),
            .in3(N__27744),
            .lcout(\phase_controller_inst1.stoper_hc.N_325 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_9_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_9_18_4 .LUT_INIT=16'b1100110011111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__28173),
            .in2(N__23531),
            .in3(N__27628),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_9_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_9_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_9_18_5 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_9_18_5  (
            .in0(N__27629),
            .in1(N__28064),
            .in2(N__23528),
            .in3(N__27599),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46031),
            .ce(N__28872),
            .sr(N__45626));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_9_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_9_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_9_18_6 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_9_18_6  (
            .in0(N__28063),
            .in1(N__28175),
            .in2(N__28310),
            .in3(N__30233),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46031),
            .ce(N__28872),
            .sr(N__45626));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_9_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_9_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_9_18_7 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_9_18_7  (
            .in0(N__28174),
            .in1(N__28065),
            .in2(N__28361),
            .in3(N__28298),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46031),
            .ce(N__28872),
            .sr(N__45626));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_19_0 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_9_19_0  (
            .in0(N__28290),
            .in1(N__28068),
            .in2(N__28343),
            .in3(N__28228),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46027),
            .ce(N__28871),
            .sr(N__45634));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_9_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_9_19_1 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB4DJ11_5_LC_9_19_1  (
            .in0(N__41711),
            .in1(N__41544),
            .in2(N__30083),
            .in3(N__28090),
            .lcout(elapsed_time_ns_1_RNIB4DJ11_0_5),
            .ltout(elapsed_time_ns_1_RNIB4DJ11_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_9_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_9_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_9_19_2 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_9_19_2  (
            .in0(N__28291),
            .in1(N__28069),
            .in2(N__23525),
            .in3(N__28229),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46027),
            .ce(N__28871),
            .sr(N__45634));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_9_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_9_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_9_19_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_9_19_4  (
            .in0(N__28292),
            .in1(N__28227),
            .in2(_gnd_net_),
            .in3(N__27707),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46027),
            .ce(N__28871),
            .sr(N__45634));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_9_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_9_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_9_19_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_9_19_5  (
            .in0(N__28226),
            .in1(N__27680),
            .in2(_gnd_net_),
            .in3(N__28294),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46027),
            .ce(N__28871),
            .sr(N__45634));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_9_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_9_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_9_19_7 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_9_19_7  (
            .in0(N__28067),
            .in1(N__28649),
            .in2(N__27650),
            .in3(N__28293),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46027),
            .ce(N__28871),
            .sr(N__45634));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_9_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_9_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_9_20_1 .LUT_INIT=16'b0101010101010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_9_20_1  (
            .in0(N__28233),
            .in1(N__23845),
            .in2(N__23833),
            .in3(N__27855),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46023),
            .ce(N__29308),
            .sr(N__45638));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_9_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_9_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_9_20_2 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_9_20_2  (
            .in0(N__23707),
            .in1(N__27856),
            .in2(_gnd_net_),
            .in3(N__28236),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46023),
            .ce(N__29308),
            .sr(N__45638));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_20_3 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_9_20_3  (
            .in0(N__28231),
            .in1(N__23776),
            .in2(_gnd_net_),
            .in3(N__27853),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46023),
            .ce(N__29308),
            .sr(N__45638));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_20_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_9_20_4  (
            .in0(N__27850),
            .in1(N__28234),
            .in2(_gnd_net_),
            .in3(N__23744),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46023),
            .ce(N__29308),
            .sr(N__45638));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_20_5 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_9_20_5  (
            .in0(N__28230),
            .in1(N__27852),
            .in2(_gnd_net_),
            .in3(N__23554),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46023),
            .ce(N__29308),
            .sr(N__45638));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_20_6 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_9_20_6  (
            .in0(N__27851),
            .in1(N__28235),
            .in2(N__23606),
            .in3(N__23572),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46023),
            .ce(N__29308),
            .sr(N__45638));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_9_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_9_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_9_20_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_9_20_7  (
            .in0(N__28232),
            .in1(N__25038),
            .in2(N__27957),
            .in3(N__27854),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46023),
            .ce(N__29308),
            .sr(N__45638));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_9_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_9_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_9_21_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_9_21_0  (
            .in0(N__28243),
            .in1(N__27939),
            .in2(N__25046),
            .in3(N__27864),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46020),
            .ce(N__28874),
            .sr(N__45642));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_9_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_9_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_9_21_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_9_21_1  (
            .in0(N__27861),
            .in1(N__28246),
            .in2(_gnd_net_),
            .in3(N__23555),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46020),
            .ce(N__28874),
            .sr(N__45642));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_9_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_9_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_9_21_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_9_21_3  (
            .in0(N__27862),
            .in1(N__28247),
            .in2(N__27761),
            .in3(N__28490),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46020),
            .ce(N__28874),
            .sr(N__45642));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_9_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_9_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_9_21_4 .LUT_INIT=16'b0101010101010001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_9_21_4  (
            .in0(N__28245),
            .in1(N__23846),
            .in2(N__23834),
            .in3(N__27865),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46020),
            .ce(N__28874),
            .sr(N__45642));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_9_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_9_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_9_21_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_9_21_6  (
            .in0(N__28244),
            .in1(N__27863),
            .in2(N__27964),
            .in3(N__26890),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46020),
            .ce(N__28874),
            .sr(N__45642));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_9_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_9_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_9_22_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_9_22_0  (
            .in0(N__27868),
            .in1(N__28241),
            .in2(N__26864),
            .in3(N__27946),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46016),
            .ce(N__28862),
            .sr(N__45649));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_9_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_9_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_9_22_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_9_22_3  (
            .in0(N__28238),
            .in1(N__27908),
            .in2(N__27958),
            .in3(N__27870),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46016),
            .ce(N__28862),
            .sr(N__45649));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_9_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_9_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_9_22_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_9_22_4  (
            .in0(N__27866),
            .in1(N__28239),
            .in2(_gnd_net_),
            .in3(N__23777),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46016),
            .ce(N__28862),
            .sr(N__45649));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_9_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_9_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_9_22_5 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_9_22_5  (
            .in0(N__28237),
            .in1(N__27869),
            .in2(_gnd_net_),
            .in3(N__23743),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46016),
            .ce(N__28862),
            .sr(N__45649));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_9_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_9_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_9_22_6 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_9_22_6  (
            .in0(N__27867),
            .in1(N__28240),
            .in2(_gnd_net_),
            .in3(N__23713),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46016),
            .ce(N__28862),
            .sr(N__45649));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_25_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_25_6 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_25_6  (
            .in0(N__28689),
            .in1(N__23677),
            .in2(_gnd_net_),
            .in3(N__23645),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_433_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S1_LC_9_28_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_9_28_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_9_28_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_9_28_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41982),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45992),
            .ce(),
            .sr(N__45662));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_10_6_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_10_6_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_10_6_3  (
            .in0(N__25827),
            .in1(N__25893),
            .in2(_gnd_net_),
            .in3(N__25920),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_10_6_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_10_6_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_10_6_4  (
            .in0(_gnd_net_),
            .in1(N__26043),
            .in2(_gnd_net_),
            .in3(N__25677),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_10_6_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_10_6_5 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_10_6_5  (
            .in0(N__25995),
            .in1(N__26019),
            .in2(N__23912),
            .in3(N__26073),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_10_6_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_10_6_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_10_6_6  (
            .in0(N__23909),
            .in1(N__25944),
            .in2(N__23903),
            .in3(N__25972),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_10_9_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_10_9_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_10_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_10_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23900),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46069),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_10_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_10_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_10_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_10_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23888),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46064),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__31074),
            .in2(_gnd_net_),
            .in3(N__29097),
            .lcout(\phase_controller_inst1.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_10_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_10_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23866),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_10_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_10_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_10_12_4 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_10_12_4  (
            .in0(N__27238),
            .in1(N__27403),
            .in2(N__27116),
            .in3(N__24290),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46050),
            .ce(),
            .sr(N__45570));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_10_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_10_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_10_12_5 .LUT_INIT=16'b0000110111011101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_10_12_5  (
            .in0(N__27402),
            .in1(N__27240),
            .in2(N__24257),
            .in3(N__27099),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46050),
            .ce(),
            .sr(N__45570));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_10_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_10_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24167),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_10_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_10_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_10_12_7 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_10_12_7  (
            .in0(N__27401),
            .in1(N__27239),
            .in2(N__24626),
            .in3(N__27098),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46050),
            .ce(),
            .sr(N__45570));
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_10_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_10_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(N__26353),
            .in2(N__26357),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_10_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_10_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_10_13_1 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_0_LC_10_13_1  (
            .in0(N__27088),
            .in1(N__24149),
            .in2(N__24134),
            .in3(N__24089),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .clk(N__46044),
            .ce(),
            .sr(N__45576));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_10_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_10_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_10_13_2 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_10_13_2  (
            .in0(N__27069),
            .in1(N__24086),
            .in2(N__26372),
            .in3(N__24080),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .clk(N__46044),
            .ce(),
            .sr(N__45576));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_10_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_10_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_10_13_3 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_10_13_3  (
            .in0(N__27089),
            .in1(N__24077),
            .in2(N__24062),
            .in3(N__24005),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .clk(N__46044),
            .ce(),
            .sr(N__45576));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_10_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_10_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_10_13_4 .LUT_INIT=16'b0111110111010111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_10_13_4  (
            .in0(N__27070),
            .in1(N__24002),
            .in2(N__23993),
            .in3(N__23930),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .clk(N__46044),
            .ce(),
            .sr(N__45576));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_10_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_10_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(N__23927),
            .in2(N__23921),
            .in3(N__24365),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_10_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_10_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(N__24362),
            .in2(N__26174),
            .in3(N__24350),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_10_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_10_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__26237),
            .in2(N__27554),
            .in3(N__24347),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_10_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_10_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__24344),
            .in2(N__24335),
            .in3(N__24311),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_10_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_10_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__24308),
            .in2(N__24299),
            .in3(N__24281),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_10_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_10_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__24278),
            .in2(N__24266),
            .in3(N__24245),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_10_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_10_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(N__26834),
            .in2(N__24242),
            .in3(N__24230),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_10_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_10_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__24227),
            .in2(N__24218),
            .in3(N__24197),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_10_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_10_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__24611),
            .in2(N__24602),
            .in3(N__24587),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_10_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_10_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__24584),
            .in2(N__24575),
            .in3(N__24560),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_10_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_10_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__26300),
            .in2(N__24557),
            .in3(N__24542),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_10_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_10_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__24539),
            .in2(N__24527),
            .in3(N__24500),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_10_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_10_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__24497),
            .in2(N__24485),
            .in3(N__24458),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_10_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_10_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__24455),
            .in2(N__24449),
            .in3(N__24422),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_10_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_10_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__24419),
            .in2(N__24407),
            .in3(N__24386),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_10_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_10_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__26243),
            .in2(N__24383),
            .in3(N__24374),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_10_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_10_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__26768),
            .in2(N__24794),
            .in3(N__24785),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_10_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_10_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__26363),
            .in2(N__26495),
            .in3(N__24782),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_10_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_10_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__26294),
            .in2(N__26603),
            .in3(N__24779),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_10_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_10_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__24890),
            .in2(N__24806),
            .in3(N__24764),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_10_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_10_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__24761),
            .in2(N__24749),
            .in3(N__24722),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_10_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_10_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(N__24719),
            .in2(N__24707),
            .in3(N__24686),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_10_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_10_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__24683),
            .in2(N__24671),
            .in3(N__24644),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_10_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_10_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(N__31361),
            .in2(N__24641),
            .in3(N__24614),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_10_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_10_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(N__31307),
            .in2(N__32857),
            .in3(N__24914),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_10_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_10_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__32853),
            .in2(N__24911),
            .in3(N__24899),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_10_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_10_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(N__31418),
            .in2(N__32858),
            .in3(N__24896),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_10_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_10_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_10_17_0  (
            .in0(N__33136),
            .in1(N__27310),
            .in2(_gnd_net_),
            .in3(N__24893),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_17_1 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE7DJ11_8_LC_10_17_1  (
            .in0(N__41716),
            .in1(N__41575),
            .in2(N__30512),
            .in3(N__27678),
            .lcout(elapsed_time_ns_1_RNIE7DJ11_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24883),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_17_3 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_17_3  (
            .in0(N__47048),
            .in1(N__47337),
            .in2(N__46397),
            .in3(N__47002),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_10_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_10_17_4 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7J_LC_10_17_4  (
            .in0(N__33135),
            .in1(N__24884),
            .in2(N__24842),
            .in3(N__24827),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIHA7JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_10_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_10_17_6 .LUT_INIT=16'b0111001100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_10_17_6  (
            .in0(N__28644),
            .in1(N__41387),
            .in2(N__24944),
            .in3(N__24959),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_10_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_10_17_7 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNID6DJ11_7_LC_10_17_7  (
            .in0(N__41715),
            .in1(N__41574),
            .in2(N__30539),
            .in3(N__27706),
            .lcout(elapsed_time_ns_1_RNID6DJ11_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_10_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_10_18_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_10_18_0  (
            .in0(N__27701),
            .in1(N__24976),
            .in2(N__27679),
            .in3(N__30232),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_10_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_10_18_1 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_10_18_1  (
            .in0(N__28480),
            .in1(_gnd_net_),
            .in2(N__24983),
            .in3(N__27811),
            .lcout(\phase_controller_inst1.stoper_hc.N_327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_10_18_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_10_18_2 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ2MD11_13_LC_10_18_2  (
            .in0(N__41519),
            .in1(N__41702),
            .in2(N__30371),
            .in3(N__27897),
            .lcout(elapsed_time_ns_1_RNIQ2MD11_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_10_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_10_18_3 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP1MD11_12_LC_10_18_3  (
            .in0(N__26847),
            .in1(N__41518),
            .in2(N__30395),
            .in3(N__41700),
            .lcout(elapsed_time_ns_1_RNIP1MD11_0_12),
            .ltout(elapsed_time_ns_1_RNIP1MD11_0_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_10_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_10_18_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_10_18_4  (
            .in0(N__25031),
            .in1(N__27896),
            .in2(N__24980),
            .in3(N__26882),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_10_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_10_18_5 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_10_18_5  (
            .in0(N__24958),
            .in1(N__28176),
            .in2(N__24943),
            .in3(N__27815),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_10_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_10_18_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_10_18_6  (
            .in0(N__28613),
            .in1(N__24957),
            .in2(N__27857),
            .in3(N__24939),
            .lcout(\phase_controller_inst1.stoper_hc.N_307 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_10_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_10_18_7 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO0MD11_11_LC_10_18_7  (
            .in0(N__26883),
            .in1(N__41701),
            .in2(N__30419),
            .in3(N__41520),
            .lcout(elapsed_time_ns_1_RNIO0MD11_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_10_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_10_19_0 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVLD11_10_LC_10_19_0  (
            .in0(N__41497),
            .in1(N__41692),
            .in2(N__30446),
            .in3(N__25042),
            .lcout(elapsed_time_ns_1_RNINVLD11_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_10_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_10_19_1 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA3DJ11_4_LC_10_19_1  (
            .in0(N__41689),
            .in1(N__41496),
            .in2(N__30107),
            .in3(N__28338),
            .lcout(elapsed_time_ns_1_RNIA3DJ11_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_10_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_10_19_2 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP2ND11_21_LC_10_19_2  (
            .in0(N__41498),
            .in1(N__25013),
            .in2(N__30608),
            .in3(N__41691),
            .lcout(elapsed_time_ns_1_RNIP2ND11_0_21),
            .ltout(elapsed_time_ns_1_RNIP2ND11_0_21_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_10_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_10_19_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_10_19_3  (
            .in0(N__25000),
            .in1(N__28507),
            .in2(N__25007),
            .in3(N__28393),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_19_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_19_4  (
            .in0(N__25124),
            .in1(N__25142),
            .in2(N__25004),
            .in3(N__25108),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_10_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_10_19_5 .LUT_INIT=16'b0000000011101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIURK5B_31_LC_10_19_5  (
            .in0(N__28007),
            .in1(N__29929),
            .in2(N__27991),
            .in3(N__30854),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_10_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_10_19_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU7ND11_26_LC_10_19_6  (
            .in0(N__41499),
            .in1(N__41693),
            .in2(N__30971),
            .in3(N__25001),
            .lcout(elapsed_time_ns_1_RNIU7ND11_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_10_19_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_10_19_7 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0AND11_28_LC_10_19_7  (
            .in0(N__41690),
            .in1(N__25136),
            .in2(N__41550),
            .in3(N__30926),
            .lcout(elapsed_time_ns_1_RNI0AND11_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_10_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_10_20_0 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIR4ND11_23_LC_10_20_0  (
            .in0(N__24992),
            .in1(N__41688),
            .in2(N__30566),
            .in3(N__41500),
            .lcout(elapsed_time_ns_1_RNIR4ND11_0_23),
            .ltout(elapsed_time_ns_1_RNIR4ND11_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_20_1  (
            .in0(N__28018),
            .in1(N__28519),
            .in2(N__24986),
            .in3(N__25117),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_20_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__25135),
            .in2(_gnd_net_),
            .in3(N__25093),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_10_20_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_10_20_3 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1BND11_29_LC_10_20_3  (
            .in0(N__41504),
            .in1(N__41695),
            .in2(N__30905),
            .in3(N__25118),
            .lcout(elapsed_time_ns_1_RNI1BND11_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_10_20_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_10_20_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO1ND11_20_LC_10_20_4  (
            .in0(N__41696),
            .in1(N__25109),
            .in2(N__41563),
            .in3(N__30629),
            .lcout(elapsed_time_ns_1_RNIO1ND11_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_10_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_10_20_5 .LUT_INIT=16'b1110101011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6_15_LC_10_20_5  (
            .in0(N__28594),
            .in1(N__28580),
            .in2(N__28412),
            .in3(N__28552),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJO4K6Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_10_20_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_10_20_6 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09_31_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__30841),
            .in2(N__25097),
            .in3(N__27984),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTG09Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_10_20_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_10_20_7 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV8ND11_27_LC_10_20_7  (
            .in0(N__25094),
            .in1(N__41694),
            .in2(N__41549),
            .in3(N__30947),
            .lcout(elapsed_time_ns_1_RNIV8ND11_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_1_c_inv_LC_10_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_1_c_inv_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_1_c_inv_LC_10_21_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_1_c_inv_LC_10_21_0  (
            .in0(N__28897),
            .in1(N__25073),
            .in2(N__25085),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_2_c_inv_LC_10_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_2_c_inv_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_2_c_inv_LC_10_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_2_c_inv_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__25067),
            .in2(N__25058),
            .in3(N__25487),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_3_c_inv_LC_10_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_3_c_inv_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_3_c_inv_LC_10_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_3_c_inv_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__25304),
            .in2(N__25295),
            .in3(N__25460),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_4_c_inv_LC_10_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_4_c_inv_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_4_c_inv_LC_10_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_4_c_inv_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__25286),
            .in2(N__25277),
            .in3(N__25442),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_5_c_inv_LC_10_21_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_5_c_inv_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_5_c_inv_LC_10_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_5_c_inv_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__25265),
            .in2(N__25256),
            .in3(N__25658),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_6_c_inv_LC_10_21_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_6_c_inv_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_6_c_inv_LC_10_21_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_6_c_inv_LC_10_21_5  (
            .in0(N__25640),
            .in1(N__25247),
            .in2(N__25238),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_7_c_inv_LC_10_21_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_7_c_inv_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_7_c_inv_LC_10_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_7_c_inv_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__25226),
            .in2(N__25217),
            .in3(N__25622),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_8_c_inv_LC_10_21_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_8_c_inv_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_8_c_inv_LC_10_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_8_c_inv_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(N__25193),
            .in2(N__25205),
            .in3(N__25604),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_9_c_inv_LC_10_22_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_9_c_inv_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_9_c_inv_LC_10_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_9_c_inv_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__25187),
            .in2(N__25172),
            .in3(N__25586),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_10_c_inv_LC_10_22_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_10_c_inv_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_10_c_inv_LC_10_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_10_c_inv_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__25160),
            .in2(N__25154),
            .in3(N__25568),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_11_c_inv_LC_10_22_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_11_c_inv_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_11_c_inv_LC_10_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_11_c_inv_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(N__25424),
            .in2(N__25418),
            .in3(N__25550),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_12_c_inv_LC_10_22_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_12_c_inv_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_12_c_inv_LC_10_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_12_c_inv_LC_10_22_3  (
            .in0(_gnd_net_),
            .in1(N__25400),
            .in2(N__25409),
            .in3(N__25532),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_13_c_inv_LC_10_22_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_13_c_inv_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_13_c_inv_LC_10_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_13_c_inv_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(N__25394),
            .in2(N__25388),
            .in3(N__25811),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_14_c_inv_LC_10_22_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_14_c_inv_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_14_c_inv_LC_10_22_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_14_c_inv_LC_10_22_5  (
            .in0(N__25793),
            .in1(N__25379),
            .in2(N__25373),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_15_c_inv_LC_10_22_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_15_c_inv_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_15_c_inv_LC_10_22_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_15_c_inv_LC_10_22_6  (
            .in0(_gnd_net_),
            .in1(N__25364),
            .in2(N__25358),
            .in3(N__25775),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_16_c_inv_LC_10_22_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_16_c_inv_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_16_c_inv_LC_10_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_16_c_inv_LC_10_22_7  (
            .in0(_gnd_net_),
            .in1(N__25349),
            .in2(N__25343),
            .in3(N__25754),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_17_c_inv_LC_10_23_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_17_c_inv_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_17_c_inv_LC_10_23_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_17_c_inv_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(N__25325),
            .in2(N__25334),
            .in3(N__25736),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_10_23_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_18_c_inv_LC_10_23_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_18_c_inv_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_18_c_inv_LC_10_23_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_18_c_inv_LC_10_23_1  (
            .in0(_gnd_net_),
            .in1(N__25319),
            .in2(N__25313),
            .in3(N__25718),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_inv_LC_10_23_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_inv_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_inv_LC_10_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_inv_LC_10_23_2  (
            .in0(_gnd_net_),
            .in1(N__25514),
            .in2(N__25508),
            .in3(N__25697),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_10_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_10_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_10_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25499),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNIV5S7_LC_10_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNIV5S7_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNIV5S7_LC_10_23_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNIV5S7_LC_10_23_5  (
            .in0(_gnd_net_),
            .in1(N__30800),
            .in2(_gnd_net_),
            .in3(N__28926),
            .lcout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_23_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_10_23_6  (
            .in0(N__28711),
            .in1(_gnd_net_),
            .in2(N__25496),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJB21_LC_10_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJB21_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJB21_LC_10_23_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJB21_LC_10_23_7  (
            .in0(_gnd_net_),
            .in1(N__28712),
            .in2(_gnd_net_),
            .in3(N__28912),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_19_c_RNINJBZ0Z21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_10_24_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_10_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_10_24_0  (
            .in0(_gnd_net_),
            .in1(N__25493),
            .in2(N__28901),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_24_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_10_24_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_10_24_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_10_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_10_24_1  (
            .in0(N__28813),
            .in1(N__25486),
            .in2(_gnd_net_),
            .in3(N__25472),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__45999),
            .ce(),
            .sr(N__45650));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_10_24_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_10_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_10_24_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_10_24_2  (
            .in0(N__28822),
            .in1(N__25459),
            .in2(N__25469),
            .in3(N__25445),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__45999),
            .ce(),
            .sr(N__45650));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_10_24_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_10_24_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_10_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_10_24_3  (
            .in0(N__28814),
            .in1(N__25441),
            .in2(_gnd_net_),
            .in3(N__25427),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__45999),
            .ce(),
            .sr(N__45650));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_10_24_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_10_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_10_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_10_24_4  (
            .in0(N__28823),
            .in1(N__25657),
            .in2(_gnd_net_),
            .in3(N__25643),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__45999),
            .ce(),
            .sr(N__45650));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_10_24_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_10_24_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_10_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_10_24_5  (
            .in0(N__28815),
            .in1(N__25639),
            .in2(_gnd_net_),
            .in3(N__25625),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__45999),
            .ce(),
            .sr(N__45650));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_10_24_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_10_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_10_24_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_10_24_6  (
            .in0(N__28824),
            .in1(N__25621),
            .in2(_gnd_net_),
            .in3(N__25607),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__45999),
            .ce(),
            .sr(N__45650));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_10_24_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_10_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_10_24_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_10_24_7  (
            .in0(N__28816),
            .in1(N__25603),
            .in2(_gnd_net_),
            .in3(N__25589),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__45999),
            .ce(),
            .sr(N__45650));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_10_25_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_10_25_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_10_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_10_25_0  (
            .in0(N__28870),
            .in1(N__25585),
            .in2(_gnd_net_),
            .in3(N__25571),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_10_25_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__45996),
            .ce(),
            .sr(N__45653));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_10_25_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_10_25_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_10_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_10_25_1  (
            .in0(N__28817),
            .in1(N__25567),
            .in2(_gnd_net_),
            .in3(N__25553),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__45996),
            .ce(),
            .sr(N__45653));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_10_25_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_10_25_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_10_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_10_25_2  (
            .in0(N__28867),
            .in1(N__25549),
            .in2(_gnd_net_),
            .in3(N__25535),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__45996),
            .ce(),
            .sr(N__45653));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_10_25_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_10_25_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_10_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_10_25_3  (
            .in0(N__28818),
            .in1(N__25531),
            .in2(_gnd_net_),
            .in3(N__25517),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__45996),
            .ce(),
            .sr(N__45653));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_10_25_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_10_25_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_10_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_10_25_4  (
            .in0(N__28868),
            .in1(N__25810),
            .in2(_gnd_net_),
            .in3(N__25796),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__45996),
            .ce(),
            .sr(N__45653));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_10_25_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_10_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_10_25_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_10_25_5  (
            .in0(N__28819),
            .in1(N__25792),
            .in2(_gnd_net_),
            .in3(N__25778),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__45996),
            .ce(),
            .sr(N__45653));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_10_25_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_10_25_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_10_25_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_10_25_6  (
            .in0(N__28869),
            .in1(N__25771),
            .in2(_gnd_net_),
            .in3(N__25757),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__45996),
            .ce(),
            .sr(N__45653));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_10_25_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_10_25_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_10_25_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_10_25_7  (
            .in0(N__28820),
            .in1(N__25753),
            .in2(_gnd_net_),
            .in3(N__25739),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__45996),
            .ce(),
            .sr(N__45653));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_10_26_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_10_26_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_10_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_10_26_0  (
            .in0(N__28866),
            .in1(N__25735),
            .in2(_gnd_net_),
            .in3(N__25721),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_10_26_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__45994),
            .ce(),
            .sr(N__45656));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_10_26_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_10_26_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_10_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_10_26_1  (
            .in0(N__28828),
            .in1(N__25717),
            .in2(_gnd_net_),
            .in3(N__25703),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__45994),
            .ce(),
            .sr(N__45656));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_10_26_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_10_26_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_10_26_2 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_10_26_2  (
            .in0(N__25696),
            .in1(N__28829),
            .in2(_gnd_net_),
            .in3(N__25700),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45994),
            .ce(),
            .sr(N__45656));
    defparam \pwm_generator_inst.counter_0_LC_11_6_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_11_6_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_11_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_11_6_0  (
            .in0(N__25871),
            .in1(N__25681),
            .in2(_gnd_net_),
            .in3(N__25661),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__46083),
            .ce(),
            .sr(N__45540));
    defparam \pwm_generator_inst.counter_1_LC_11_6_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_11_6_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_11_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_11_6_1  (
            .in0(N__25865),
            .in1(N__26074),
            .in2(_gnd_net_),
            .in3(N__26051),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__46083),
            .ce(),
            .sr(N__45540));
    defparam \pwm_generator_inst.counter_2_LC_11_6_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_11_6_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_11_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_11_6_2  (
            .in0(N__25872),
            .in1(N__26047),
            .in2(_gnd_net_),
            .in3(N__26027),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__46083),
            .ce(),
            .sr(N__45540));
    defparam \pwm_generator_inst.counter_3_LC_11_6_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_11_6_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_11_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_11_6_3  (
            .in0(N__25866),
            .in1(N__26020),
            .in2(_gnd_net_),
            .in3(N__26000),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__46083),
            .ce(),
            .sr(N__45540));
    defparam \pwm_generator_inst.counter_4_LC_11_6_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_11_6_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_11_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_11_6_4  (
            .in0(N__25873),
            .in1(N__25996),
            .in2(_gnd_net_),
            .in3(N__25976),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__46083),
            .ce(),
            .sr(N__45540));
    defparam \pwm_generator_inst.counter_5_LC_11_6_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_11_6_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_11_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_11_6_5  (
            .in0(N__25867),
            .in1(N__25971),
            .in2(_gnd_net_),
            .in3(N__25952),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__46083),
            .ce(),
            .sr(N__45540));
    defparam \pwm_generator_inst.counter_6_LC_11_6_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_11_6_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_11_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_11_6_6  (
            .in0(N__25874),
            .in1(N__25948),
            .in2(_gnd_net_),
            .in3(N__25925),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__46083),
            .ce(),
            .sr(N__45540));
    defparam \pwm_generator_inst.counter_7_LC_11_6_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_11_6_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_11_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_11_6_7  (
            .in0(N__25868),
            .in1(N__25921),
            .in2(_gnd_net_),
            .in3(N__25901),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__46083),
            .ce(),
            .sr(N__45540));
    defparam \pwm_generator_inst.counter_8_LC_11_7_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_11_7_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_11_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_11_7_0  (
            .in0(N__25870),
            .in1(N__25897),
            .in2(_gnd_net_),
            .in3(N__25877),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__46075),
            .ce(),
            .sr(N__45545));
    defparam \pwm_generator_inst.counter_9_LC_11_7_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_11_7_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_11_7_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_11_7_1  (
            .in0(N__25831),
            .in1(N__25869),
            .in2(_gnd_net_),
            .in3(N__25835),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46075),
            .ce(),
            .sr(N__45545));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__28983),
            .in2(_gnd_net_),
            .in3(N__28964),
            .lcout(\phase_controller_inst1.N_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_11_10_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_10_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_10_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_11_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_11_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27510),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_11_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_11_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__31294),
            .in2(_gnd_net_),
            .in3(N__29083),
            .lcout(\phase_controller_inst1.N_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36878),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_11_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_11_13_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIJD8U_9_LC_11_13_0  (
            .in0(N__33116),
            .in1(N__26134),
            .in2(N__26216),
            .in3(N__26186),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIJD8UZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_11_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_11_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_11_13_2 .LUT_INIT=16'b0101111100010011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_11_13_2  (
            .in0(N__27082),
            .in1(N__27374),
            .in2(N__26162),
            .in3(N__27249),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46037),
            .ce(),
            .sr(N__45571));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_11_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_11_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_11_13_3 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_11_13_3  (
            .in0(N__27370),
            .in1(N__27083),
            .in2(N__27256),
            .in3(N__26096),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46037),
            .ce(),
            .sr(N__45571));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_11_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_11_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_11_13_4 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_11_13_4  (
            .in0(N__27080),
            .in1(N__27372),
            .in2(N__26087),
            .in3(N__27247),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46037),
            .ce(),
            .sr(N__45571));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_11_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_11_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_11_13_5 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_11_13_5  (
            .in0(N__27371),
            .in1(N__27084),
            .in2(N__27257),
            .in3(N__26483),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46037),
            .ce(),
            .sr(N__45571));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_11_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_11_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_11_13_6 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_11_13_6  (
            .in0(N__27081),
            .in1(N__27373),
            .in2(N__26474),
            .in3(N__27248),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46037),
            .ce(),
            .sr(N__45571));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_11_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_11_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26460),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_11_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_11_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26393),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_11_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_11_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26533),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_11_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_11_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_0_12_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33112),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_11_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_11_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26338),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_11_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_11_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26668),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_11_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_11_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26272),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_11_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_11_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26902),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37109),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_11_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_11_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26804),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_11_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_11_15_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__26754),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37166),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_15_5  (
            .in0(N__26703),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33068),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_11_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_11_15_6 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76J_LC_11_15_6  (
            .in0(N__26678),
            .in1(N__26645),
            .in2(N__33125),
            .in3(N__26615),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIF76JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_11_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_11_15_7 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45J_LC_11_15_7  (
            .in0(N__26594),
            .in1(N__26549),
            .in2(N__26510),
            .in3(N__33069),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNID45JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_16_0 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI5R941_10_LC_11_16_0  (
            .in0(N__27509),
            .in1(N__27586),
            .in2(N__33134),
            .in3(N__27563),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI5R941Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_11_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_11_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_11_16_2 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_11_16_2  (
            .in0(N__27252),
            .in1(N__27327),
            .in2(N__27119),
            .in3(N__27539),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46029),
            .ce(),
            .sr(N__45588));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_11_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_11_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_11_16_3 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_11_16_3  (
            .in0(N__27323),
            .in1(N__27254),
            .in2(N__27479),
            .in3(N__27110),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46029),
            .ce(),
            .sr(N__45588));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_11_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_11_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_11_16_4 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_11_16_4  (
            .in0(N__27250),
            .in1(N__27325),
            .in2(N__27117),
            .in3(N__27470),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46029),
            .ce(),
            .sr(N__45588));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_11_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_11_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_11_16_5 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_11_16_5  (
            .in0(N__27324),
            .in1(N__27255),
            .in2(N__27419),
            .in3(N__27111),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46029),
            .ce(),
            .sr(N__45588));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_11_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_11_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_11_16_6 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_11_16_6  (
            .in0(N__27251),
            .in1(N__27326),
            .in2(N__27118),
            .in3(N__27410),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46029),
            .ce(),
            .sr(N__45588));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_11_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_11_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_11_16_7 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_11_16_7  (
            .in0(N__27322),
            .in1(N__27253),
            .in2(N__27134),
            .in3(N__27109),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46029),
            .ce(),
            .sr(N__45588));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_11_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_11_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_11_17_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_11_17_0  (
            .in0(N__28168),
            .in1(N__27959),
            .in2(N__26891),
            .in3(N__27873),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46024),
            .ce(N__29309),
            .sr(N__45592));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_11_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_11_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_11_17_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_11_17_1  (
            .in0(N__27871),
            .in1(N__28171),
            .in2(N__27965),
            .in3(N__26863),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46024),
            .ce(N__29309),
            .sr(N__45592));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_17_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_11_17_2  (
            .in0(N__28169),
            .in1(N__27960),
            .in2(N__27907),
            .in3(N__27874),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46024),
            .ce(N__29309),
            .sr(N__45592));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_17_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_11_17_3  (
            .in0(N__27872),
            .in1(N__28172),
            .in2(N__28495),
            .in3(N__27760),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46024),
            .ce(N__29309),
            .sr(N__45592));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_11_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_11_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_11_17_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_11_17_4  (
            .in0(N__28167),
            .in1(N__27702),
            .in2(_gnd_net_),
            .in3(N__28313),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46024),
            .ce(N__29309),
            .sr(N__45592));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_11_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_11_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_11_17_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_11_17_5  (
            .in0(N__28311),
            .in1(N__28170),
            .in2(_gnd_net_),
            .in3(N__27677),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46024),
            .ce(N__29309),
            .sr(N__45592));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_11_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_11_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_11_17_6 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_11_17_6  (
            .in0(N__28066),
            .in1(N__28645),
            .in2(N__27649),
            .in3(N__28312),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46024),
            .ce(N__29309),
            .sr(N__45592));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_17_7 .LUT_INIT=16'b0001110100011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_17_7  (
            .in0(N__33281),
            .in1(N__42191),
            .in2(N__33425),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_11_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_11_18_0 .LUT_INIT=16'b1111111101011100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITCMJQ_1_LC_11_18_0  (
            .in0(N__33800),
            .in1(N__27622),
            .in2(N__41564),
            .in3(N__30186),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_11_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_11_18_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDP2KD1_1_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27632),
            .in3(N__30281),
            .lcout(elapsed_time_ns_1_RNIDP2KD1_0_1),
            .ltout(elapsed_time_ns_1_RNIDP2KD1_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_11_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_11_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_11_18_2 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_11_18_2  (
            .in0(N__28056),
            .in1(N__27611),
            .in2(N__27602),
            .in3(N__27598),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46021),
            .ce(N__29304),
            .sr(N__45599));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_11_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_11_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_11_18_3 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_11_18_3  (
            .in0(N__28308),
            .in1(N__28061),
            .in2(N__30231),
            .in3(N__28166),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46021),
            .ce(N__29304),
            .sr(N__45599));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_11_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_11_18_4 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ4OD11_31_LC_11_18_4  (
            .in0(N__28163),
            .in1(N__41710),
            .in2(N__30857),
            .in3(N__41530),
            .lcout(elapsed_time_ns_1_RNIQ4OD11_0_31),
            .ltout(elapsed_time_ns_1_RNIQ4OD11_0_31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_11_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_11_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_11_18_5 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_11_18_5  (
            .in0(N__28306),
            .in1(N__28060),
            .in2(N__28364),
            .in3(N__28354),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46021),
            .ce(N__29304),
            .sr(N__45599));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_11_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_11_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_11_18_6 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_11_18_6  (
            .in0(N__28164),
            .in1(N__28337),
            .in2(N__28070),
            .in3(N__28309),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46021),
            .ce(N__29304),
            .sr(N__45599));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_11_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_11_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_11_18_7 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_11_18_7  (
            .in0(N__28307),
            .in1(N__28165),
            .in2(N__28097),
            .in3(N__28062),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46021),
            .ce(N__29304),
            .sr(N__45599));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_11_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_11_19_0 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP3OD11_30_LC_11_19_0  (
            .in0(N__28019),
            .in1(N__41697),
            .in2(N__41551),
            .in3(N__30881),
            .lcout(elapsed_time_ns_1_RNIP3OD11_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_11_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_11_19_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847_31_LC_11_19_1  (
            .in0(N__30856),
            .in1(N__45720),
            .in2(_gnd_net_),
            .in3(N__28006),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOG847Z0Z_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_11_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_11_19_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5I_31_LC_11_19_2  (
            .in0(N__29875),
            .in1(N__45718),
            .in2(N__27995),
            .in3(N__28529),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8FB5IZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_11_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_11_19_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642_6_LC_11_19_3  (
            .in0(N__30471),
            .in1(N__30057),
            .in2(N__28411),
            .in3(N__30336),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICM642Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_11_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_11_19_4 .LUT_INIT=16'b1011000010100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4_31_LC_11_19_4  (
            .in0(N__45719),
            .in1(N__30855),
            .in2(N__28532),
            .in3(N__29925),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIICEP4Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_11_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_11_19_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK670F_31_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__28378),
            .in2(_gnd_net_),
            .in3(N__29874),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_382_i ),
            .ltout(\delay_measurement_inst.delay_hc_timer.N_382_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_11_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_11_19_6 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS5ND11_24_LC_11_19_6  (
            .in0(N__31016),
            .in1(N__28520),
            .in2(N__28523),
            .in3(N__41698),
            .lcout(elapsed_time_ns_1_RNIS5ND11_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_11_19_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_11_19_7 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIT6ND11_25_LC_11_19_7  (
            .in0(N__41699),
            .in1(N__28508),
            .in2(N__30995),
            .in3(N__41511),
            .lcout(elapsed_time_ns_1_RNIT6ND11_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_11_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_11_20_0 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS4MD11_15_LC_11_20_0  (
            .in0(N__28461),
            .in1(N__41522),
            .in2(N__30305),
            .in3(N__41704),
            .lcout(elapsed_time_ns_1_RNIS4MD11_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_11_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_11_20_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_11_20_1  (
            .in0(N__30684),
            .in1(N__30720),
            .in2(N__30661),
            .in3(N__30750),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_11_20_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_11_20_2 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQ3ND11_22_LC_11_20_2  (
            .in0(N__28394),
            .in1(N__41703),
            .in2(N__41573),
            .in3(N__30584),
            .lcout(elapsed_time_ns_1_RNIQ3ND11_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_11_20_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_11_20_3 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58F_31_LC_11_20_3  (
            .in0(N__45721),
            .in1(_gnd_net_),
            .in2(N__28382),
            .in3(N__29870),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRF58FZ0Z_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_11_20_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_11_20_4 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIS27MU_3_LC_11_20_4  (
            .in0(N__28643),
            .in1(N__41523),
            .in2(N__28367),
            .in3(N__30122),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_11_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_11_20_5 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQURR91_3_LC_11_20_5  (
            .in0(N__30185),
            .in1(_gnd_net_),
            .in2(N__28652),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIQURR91_0_3),
            .ltout(elapsed_time_ns_1_RNIQURR91_0_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_11_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_11_20_6 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_11_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28616),
            .in3(N__41386),
            .lcout(\phase_controller_inst1.stoper_hc.N_283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_11_21_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_11_21_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992_24_LC_11_21_0  (
            .in0(N__30985),
            .in1(N__28538),
            .in2(N__31015),
            .in3(N__28934),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7O992Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_11_21_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_11_21_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91_7_LC_11_21_1  (
            .in0(N__30529),
            .in1(N__30470),
            .in2(_gnd_net_),
            .in3(N__30502),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMKF91Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_11_21_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_11_21_2 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2_15_LC_11_21_2  (
            .in0(N__30301),
            .in1(N__28574),
            .in2(N__28583),
            .in3(N__30335),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7V3Q2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_11_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_11_21_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_11_21_3  (
            .in0(N__30385),
            .in1(N__30409),
            .in2(N__30439),
            .in3(N__30361),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_11_21_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_11_21_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542_15_LC_11_21_4  (
            .in0(N__30501),
            .in1(N__30528),
            .in2(N__28568),
            .in3(N__30300),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU542Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_11_21_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_11_21_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_11_21_7  (
            .in0(N__30598),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30580),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lt31_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_11_22_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_11_22_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9PDO_26_LC_11_22_1  (
            .in0(N__30919),
            .in1(N__30940),
            .in2(_gnd_net_),
            .in3(N__30961),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_11_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_11_22_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITTI01_20_LC_11_22_5  (
            .in0(N__30895),
            .in1(N__30622),
            .in2(N__30559),
            .in3(N__30874),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_0_sqmuxa_0_o2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_2_LC_11_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_11_23_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_11_23_4 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst2.state_2_LC_11_23_4  (
            .in0(N__33722),
            .in1(N__41830),
            .in2(N__41987),
            .in3(N__41879),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46000),
            .ce(),
            .sr(N__45639));
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_23_5 .LUT_INIT=16'b1100111001001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_11_23_5  (
            .in0(N__28713),
            .in1(N__28733),
            .in2(N__30799),
            .in3(N__28927),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46000),
            .ce(),
            .sr(N__45639));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_23_6 .LUT_INIT=16'b1101110000001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_11_23_6  (
            .in0(N__28928),
            .in1(N__41880),
            .in2(N__28721),
            .in3(N__30795),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46000),
            .ce(),
            .sr(N__45639));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_23_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_23_7 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_23_7  (
            .in0(N__28821),
            .in1(N__28913),
            .in2(N__28720),
            .in3(N__28896),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46000),
            .ce(),
            .sr(N__45639));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_11_24_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_11_24_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_11_24_5  (
            .in0(N__33747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30791),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_24_6 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_11_24_6  (
            .in0(N__30790),
            .in1(N__33746),
            .in2(_gnd_net_),
            .in3(N__28732),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_11_25_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_11_25_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_11_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28691),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S2_LC_11_29_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_11_29_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_11_29_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_11_29_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46243),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45990),
            .ce(),
            .sr(N__45658));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_12_8_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_12_8_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_12_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_12_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29018),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46063),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_9_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__43846),
            .in2(_gnd_net_),
            .in3(N__43925),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_12_9_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_12_9_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_12_9_1.LUT_INIT=16'b1100110011001100;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_12_9_1 (
            .in0(_gnd_net_),
            .in1(N__29006),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46057),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__31238),
            .in2(_gnd_net_),
            .in3(N__29064),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_LC_12_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_12_10_2 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_12_10_2  (
            .in0(N__28997),
            .in1(N__28991),
            .in2(N__43678),
            .in3(N__43926),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46049),
            .ce(),
            .sr(N__45553));
    defparam \phase_controller_inst1.state_1_LC_12_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_12_10_3 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst1.state_1_LC_12_10_3  (
            .in0(N__28985),
            .in1(N__31073),
            .in2(N__28970),
            .in3(N__29104),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46049),
            .ce(),
            .sr(N__45553));
    defparam \phase_controller_inst1.state_2_LC_12_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_12_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_12_10_6 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_inst1.state_2_LC_12_10_6  (
            .in0(N__29072),
            .in1(N__28969),
            .in2(N__31252),
            .in3(N__28984),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46049),
            .ce(),
            .sr(N__45553));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_12_11_1 .LUT_INIT=16'b1010001011100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_12_11_1  (
            .in0(N__28965),
            .in1(N__43897),
            .in2(N__43850),
            .in3(N__43792),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46043),
            .ce(),
            .sr(N__45558));
    defparam \phase_controller_inst1.start_timer_tr_LC_12_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_12_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_12_11_2 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_12_11_2  (
            .in0(N__43663),
            .in1(N__29050),
            .in2(N__32735),
            .in3(N__28946),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46043),
            .ce(),
            .sr(N__45558));
    defparam \phase_controller_inst1.state_0_LC_12_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_12_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_12_11_3 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \phase_controller_inst1.state_0_LC_12_11_3  (
            .in0(N__29108),
            .in1(N__31078),
            .in2(N__31298),
            .in3(N__29084),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46043),
            .ce(),
            .sr(N__45558));
    defparam \phase_controller_inst1.state_3_LC_12_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_12_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_12_11_4 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \phase_controller_inst1.state_3_LC_12_11_4  (
            .in0(N__40517),
            .in1(N__29071),
            .in2(N__31256),
            .in3(N__29051),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46043),
            .ce(),
            .sr(N__45558));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__43895),
            .in2(_gnd_net_),
            .in3(N__29320),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNITEL9_LC_12_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNITEL9_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNITEL9_LC_12_12_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNITEL9_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__43845),
            .in2(_gnd_net_),
            .in3(N__43782),
            .lcout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNII3D41_LC_12_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNII3D41_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNII3D41_LC_12_12_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNII3D41_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29042),
            .in3(N__43896),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_19_c_RNII3DZ0Z41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_12_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_12_12_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_12_12_5  (
            .in0(N__32720),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33245),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__29167),
            .in2(N__29039),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_12_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_12_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_12_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_12_13_1  (
            .in0(N__29273),
            .in1(N__29566),
            .in2(_gnd_net_),
            .in3(N__29030),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__46034),
            .ce(),
            .sr(N__45566));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_12_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_12_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_12_13_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_12_13_2  (
            .in0(N__29277),
            .in1(N__29027),
            .in2(N__29537),
            .in3(N__29021),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__46034),
            .ce(),
            .sr(N__45566));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_13_3  (
            .in0(N__29274),
            .in1(N__29509),
            .in2(_gnd_net_),
            .in3(N__29135),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__46034),
            .ce(),
            .sr(N__45566));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_13_4  (
            .in0(N__29278),
            .in1(N__29467),
            .in2(_gnd_net_),
            .in3(N__29132),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__46034),
            .ce(),
            .sr(N__45566));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_12_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_12_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_12_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_12_13_5  (
            .in0(N__29275),
            .in1(N__29434),
            .in2(_gnd_net_),
            .in3(N__29129),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__46034),
            .ce(),
            .sr(N__45566));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_13_6  (
            .in0(N__29279),
            .in1(N__29407),
            .in2(_gnd_net_),
            .in3(N__29126),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__46034),
            .ce(),
            .sr(N__45566));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_12_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_12_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_12_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_12_13_7  (
            .in0(N__29276),
            .in1(N__29368),
            .in2(_gnd_net_),
            .in3(N__29123),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__46034),
            .ce(),
            .sr(N__45566));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_14_0  (
            .in0(N__29287),
            .in1(N__29833),
            .in2(_gnd_net_),
            .in3(N__29120),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__46032),
            .ce(),
            .sr(N__45572));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_12_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_12_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_12_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_12_14_1  (
            .in0(N__29280),
            .in1(N__29794),
            .in2(_gnd_net_),
            .in3(N__29117),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__46032),
            .ce(),
            .sr(N__45572));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_14_2  (
            .in0(N__29284),
            .in1(N__29764),
            .in2(_gnd_net_),
            .in3(N__29114),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__46032),
            .ce(),
            .sr(N__45572));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_12_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_12_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_12_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_12_14_3  (
            .in0(N__29281),
            .in1(N__29734),
            .in2(_gnd_net_),
            .in3(N__29111),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__46032),
            .ce(),
            .sr(N__45572));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_12_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_12_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_12_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_12_14_4  (
            .in0(N__29285),
            .in1(N__29704),
            .in2(_gnd_net_),
            .in3(N__29345),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__46032),
            .ce(),
            .sr(N__45572));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_12_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_12_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_12_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_12_14_5  (
            .in0(N__29282),
            .in1(N__29671),
            .in2(_gnd_net_),
            .in3(N__29342),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__46032),
            .ce(),
            .sr(N__45572));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_12_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_12_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_12_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_12_14_6  (
            .in0(N__29286),
            .in1(N__29647),
            .in2(_gnd_net_),
            .in3(N__29339),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__46032),
            .ce(),
            .sr(N__45572));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_12_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_12_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_12_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_12_14_7  (
            .in0(N__29283),
            .in1(N__29602),
            .in2(_gnd_net_),
            .in3(N__29336),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__46032),
            .ce(),
            .sr(N__45572));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_12_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_12_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_12_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_12_15_0  (
            .in0(N__29297),
            .in1(N__30028),
            .in2(_gnd_net_),
            .in3(N__29333),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__46028),
            .ce(),
            .sr(N__45577));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_12_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_12_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_12_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_12_15_1  (
            .in0(N__29299),
            .in1(N__29992),
            .in2(_gnd_net_),
            .in3(N__29330),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__46028),
            .ce(),
            .sr(N__45577));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_12_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_12_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_12_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_12_15_2  (
            .in0(N__29298),
            .in1(N__29956),
            .in2(_gnd_net_),
            .in3(N__29327),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46028),
            .ce(),
            .sr(N__45577));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_15_4 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_15_4  (
            .in0(N__43901),
            .in1(N__29324),
            .in2(N__29168),
            .in3(N__29300),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46028),
            .ce(),
            .sr(N__45577));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_1_c_inv_LC_12_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_1_c_inv_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_1_c_inv_LC_12_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_1_c_inv_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__29183),
            .in2(N__29144),
            .in3(N__29160),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_2_c_inv_LC_12_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_2_c_inv_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_2_c_inv_LC_12_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_2_c_inv_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__29579),
            .in2(N__29552),
            .in3(N__29570),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_3_c_inv_LC_12_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_3_c_inv_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_3_c_inv_LC_12_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_3_c_inv_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__29543),
            .in2(N__29519),
            .in3(N__29536),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_4_c_inv_LC_12_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_4_c_inv_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_4_c_inv_LC_12_16_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_4_c_inv_LC_12_16_3  (
            .in0(N__29510),
            .in1(N__29495),
            .in2(N__29486),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_5_c_inv_LC_12_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_5_c_inv_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_5_c_inv_LC_12_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_5_c_inv_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__29477),
            .in2(N__29453),
            .in3(N__29468),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_6_c_inv_LC_12_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_6_c_inv_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_6_c_inv_LC_12_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_6_c_inv_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__29444),
            .in2(N__29420),
            .in3(N__29435),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_7_c_inv_LC_12_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_7_c_inv_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_7_c_inv_LC_12_16_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_7_c_inv_LC_12_16_6  (
            .in0(N__29408),
            .in1(N__29384),
            .in2(N__29393),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_8_c_inv_LC_12_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_8_c_inv_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_8_c_inv_LC_12_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_8_c_inv_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(N__29354),
            .in2(N__29378),
            .in3(N__29369),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_9_c_inv_LC_12_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_9_c_inv_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_9_c_inv_LC_12_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_9_c_inv_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__29846),
            .in2(N__29819),
            .in3(N__29834),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_10_c_inv_LC_12_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_10_c_inv_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_10_c_inv_LC_12_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_10_c_inv_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__29780),
            .in2(N__29810),
            .in3(N__29795),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_11_c_inv_LC_12_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_11_c_inv_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_11_c_inv_LC_12_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_11_c_inv_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__29750),
            .in2(N__29774),
            .in3(N__29765),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_12_c_inv_LC_12_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_12_c_inv_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_12_c_inv_LC_12_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_12_c_inv_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__29720),
            .in2(N__29744),
            .in3(N__29735),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_13_c_inv_LC_12_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_13_c_inv_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_13_c_inv_LC_12_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_13_c_inv_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(N__29690),
            .in2(N__29714),
            .in3(N__29705),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_14_c_inv_LC_12_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_14_c_inv_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_14_c_inv_LC_12_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_14_c_inv_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(N__29684),
            .in2(N__29657),
            .in3(N__29672),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_15_c_inv_LC_12_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_15_c_inv_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_15_c_inv_LC_12_17_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_15_c_inv_LC_12_17_6  (
            .in0(N__29648),
            .in1(N__29633),
            .in2(N__29627),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_16_c_inv_LC_12_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_16_c_inv_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_16_c_inv_LC_12_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_16_c_inv_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__29615),
            .in2(N__29588),
            .in3(N__29603),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_17_c_inv_LC_12_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_17_c_inv_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_17_c_inv_LC_12_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_17_c_inv_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__30041),
            .in2(N__30014),
            .in3(N__30029),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_18_c_inv_LC_12_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_18_c_inv_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_18_c_inv_LC_12_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_18_c_inv_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(N__30005),
            .in2(N__29978),
            .in3(N__29993),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_inv_LC_12_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_inv_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_inv_LC_12_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_19_c_inv_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__29969),
            .in2(N__29942),
            .in3(N__29957),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_12_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_12_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_LUT4_0_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29933),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_12_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_12_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352_1_LC_12_19_0  (
            .in0(N__30121),
            .in1(N__33796),
            .in2(N__41605),
            .in3(N__30131),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1U352Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_12_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_12_19_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKR_2_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(N__30120),
            .in2(_gnd_net_),
            .in3(N__41601),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPNKRZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_12_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_12_19_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU4A94_9_LC_12_19_2  (
            .in0(N__30472),
            .in1(N__30130),
            .in2(N__29903),
            .in3(N__29896),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_12_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_12_19_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_17_LC_12_19_3  (
            .in0(N__30137),
            .in1(N__30657),
            .in2(N__29879),
            .in3(N__30727),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_12_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_12_19_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIU2KD1_6_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(N__30143),
            .in2(_gnd_net_),
            .in3(N__30280),
            .lcout(elapsed_time_ns_1_RNIIU2KD1_0_6),
            .ltout(elapsed_time_ns_1_RNIIU2KD1_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_12_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_12_19_5 .LUT_INIT=16'b1110111011111010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2IMJQ_6_LC_12_19_5  (
            .in0(N__30201),
            .in1(N__30059),
            .in2(N__30146),
            .in3(N__41521),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_12_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_12_19_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJV461_16_LC_12_19_6  (
            .in0(N__30058),
            .in1(N__30691),
            .in2(N__30763),
            .in3(N__30340),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_i_0_a2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_12_19_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_12_19_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_4_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(N__30073),
            .in2(_gnd_net_),
            .in3(N__30097),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKRZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_12_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_12_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_12_20_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__31572),
            .in2(N__33823),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__46009),
            .ce(N__33773),
            .sr(N__45605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_12_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_12_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_12_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(N__31548),
            .in2(N__31603),
            .in3(N__30086),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__46009),
            .ce(N__33773),
            .sr(N__45605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_12_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_12_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_12_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(N__31524),
            .in2(N__31577),
            .in3(N__30062),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__46009),
            .ce(N__33773),
            .sr(N__45605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_12_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_12_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_12_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(N__31815),
            .in2(N__31553),
            .in3(N__30044),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__46009),
            .ce(N__33773),
            .sr(N__45605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_12_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_12_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_12_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(N__31794),
            .in2(N__31529),
            .in3(N__30515),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__46009),
            .ce(N__33773),
            .sr(N__45605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_12_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_12_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_12_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(N__31776),
            .in2(N__31820),
            .in3(N__30488),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__46009),
            .ce(N__33773),
            .sr(N__45605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_12_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_12_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_12_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(N__31795),
            .in2(N__31760),
            .in3(N__30449),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__46009),
            .ce(N__33773),
            .sr(N__45605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_12_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_12_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_12_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(N__31777),
            .in2(N__31730),
            .in3(N__30422),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__46009),
            .ce(N__33773),
            .sr(N__45605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_12_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_12_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_12_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(N__31695),
            .in2(N__31759),
            .in3(N__30398),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_12_21_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__46003),
            .ce(N__33771),
            .sr(N__45619));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_12_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_12_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_12_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(N__31671),
            .in2(N__31729),
            .in3(N__30374),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__46003),
            .ce(N__33771),
            .sr(N__45619));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_12_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_12_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_12_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(N__31647),
            .in2(N__31700),
            .in3(N__30350),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__46003),
            .ce(N__33771),
            .sr(N__45619));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_12_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_12_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_12_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_12_21_3  (
            .in0(_gnd_net_),
            .in1(N__32019),
            .in2(N__31676),
            .in3(N__30308),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__46003),
            .ce(N__33771),
            .sr(N__45619));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_12_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_12_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_12_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_12_21_4  (
            .in0(_gnd_net_),
            .in1(N__31998),
            .in2(N__31652),
            .in3(N__30284),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc5lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__46003),
            .ce(N__33771),
            .sr(N__45619));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_12_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_12_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_12_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(N__31980),
            .in2(N__32024),
            .in3(N__30734),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__46003),
            .ce(N__33771),
            .sr(N__45619));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_12_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_12_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_12_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_12_21_6  (
            .in0(_gnd_net_),
            .in1(N__31999),
            .in2(N__31964),
            .in3(N__30704),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__46003),
            .ce(N__33771),
            .sr(N__45619));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_12_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_12_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_12_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(N__31981),
            .in2(N__31931),
            .in3(N__30668),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__46003),
            .ce(N__33771),
            .sr(N__45619));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_12_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_12_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_12_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(N__31901),
            .in2(N__31960),
            .in3(N__30632),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_12_22_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__45998),
            .ce(N__33770),
            .sr(N__45630));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_12_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_12_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_12_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_12_22_1  (
            .in0(_gnd_net_),
            .in1(N__31866),
            .in2(N__31930),
            .in3(N__30611),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__45998),
            .ce(N__33770),
            .sr(N__45630));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_12_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_12_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_12_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(N__31842),
            .in2(N__31900),
            .in3(N__30587),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__45998),
            .ce(N__33770),
            .sr(N__45630));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_12_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_12_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_12_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_12_22_3  (
            .in0(_gnd_net_),
            .in1(N__32346),
            .in2(N__31871),
            .in3(N__30569),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__45998),
            .ce(N__33770),
            .sr(N__45630));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_12_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_12_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_12_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(N__32325),
            .in2(N__31847),
            .in3(N__30542),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__45998),
            .ce(N__33770),
            .sr(N__45630));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_12_22_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_12_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_12_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_12_22_5  (
            .in0(_gnd_net_),
            .in1(N__32307),
            .in2(N__32351),
            .in3(N__30998),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__45998),
            .ce(N__33770),
            .sr(N__45630));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_12_22_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_12_22_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_12_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_12_22_6  (
            .in0(_gnd_net_),
            .in1(N__32326),
            .in2(N__32291),
            .in3(N__30974),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__45998),
            .ce(N__33770),
            .sr(N__45630));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_12_22_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_12_22_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_12_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_12_22_7  (
            .in0(_gnd_net_),
            .in1(N__32308),
            .in2(N__32261),
            .in3(N__30950),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__45998),
            .ce(N__33770),
            .sr(N__45630));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_12_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_12_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_12_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_12_23_0  (
            .in0(_gnd_net_),
            .in1(N__32226),
            .in2(N__32290),
            .in3(N__30929),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_12_23_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__45995),
            .ce(N__33769),
            .sr(N__45635));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_12_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_12_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_12_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_12_23_1  (
            .in0(_gnd_net_),
            .in1(N__32202),
            .in2(N__32260),
            .in3(N__30908),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__45995),
            .ce(N__33769),
            .sr(N__45635));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_12_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_12_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_12_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_12_23_2  (
            .in0(_gnd_net_),
            .in1(N__32182),
            .in2(N__32231),
            .in3(N__30884),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__45995),
            .ce(N__33769),
            .sr(N__45635));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_12_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_12_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_12_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_12_23_3  (
            .in0(_gnd_net_),
            .in1(N__32035),
            .in2(N__32207),
            .in3(N__30863),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__45995),
            .ce(N__33769),
            .sr(N__45635));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_12_23_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_12_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_12_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_12_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30860),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45995),
            .ce(N__33769),
            .sr(N__45635));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_12_24_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_12_24_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_12_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_12_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33748),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45993),
            .ce(),
            .sr(N__45640));
    defparam \phase_controller_inst1.S2_LC_12_26_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_12_26_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_12_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_12_26_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31079),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45991),
            .ce(),
            .sr(N__45651));
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_0 .C_ON=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_0 .SEQ_MODE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_0  (
            .in0(N__45725),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pll_inst.red_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_13_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_13_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_13_7_0 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_13_7_0  (
            .in0(N__39895),
            .in1(N__32494),
            .in2(N__32577),
            .in3(N__33997),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46076),
            .ce(N__44290),
            .sr(N__45536));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_13_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_13_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_13_7_1 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_13_7_1  (
            .in0(N__33995),
            .in1(N__39371),
            .in2(N__32576),
            .in3(N__39896),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46076),
            .ce(N__44290),
            .sr(N__45536));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_13_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_13_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_13_7_2 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_13_7_2  (
            .in0(N__38592),
            .in1(N__32560),
            .in2(N__31127),
            .in3(N__33996),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46076),
            .ce(N__44290),
            .sr(N__45536));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_13_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_13_7_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__38591),
            .in2(_gnd_net_),
            .in3(N__35913),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_13_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_13_8_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_13_8_0  (
            .in0(N__32505),
            .in1(N__31103),
            .in2(N__39729),
            .in3(N__31022),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_13_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_13_8_1 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_13_8_1  (
            .in0(N__31102),
            .in1(N__38599),
            .in2(N__35924),
            .in3(N__32507),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_13_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_13_8_2 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_13_8_2  (
            .in0(N__32506),
            .in1(N__39888),
            .in2(N__39728),
            .in3(N__31101),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_13_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_13_8_3 .LUT_INIT=16'b1110111011111010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_13_8_3  (
            .in0(N__42737),
            .in1(N__39068),
            .in2(N__32386),
            .in3(N__43168),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_13_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_13_8_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUKL2M1_6_LC_13_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31109),
            .in3(N__39138),
            .lcout(elapsed_time_ns_1_RNIUKL2M1_0_6),
            .ltout(elapsed_time_ns_1_RNIUKL2M1_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_13_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_13_8_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_13_8_5  (
            .in0(N__39198),
            .in1(N__38966),
            .in2(N__31106),
            .in3(N__34049),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_13_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_13_8_6 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_13_8_6  (
            .in0(N__39673),
            .in1(_gnd_net_),
            .in2(N__31091),
            .in3(N__34177),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_13_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_13_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_13_8_7 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_13_8_7  (
            .in0(N__39889),
            .in1(N__32382),
            .in2(N__31088),
            .in3(N__34001),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46070),
            .ce(N__44293),
            .sr(N__45541));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_13_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_13_9_0 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_13_9_0  (
            .in0(N__39919),
            .in1(N__43152),
            .in2(N__36206),
            .in3(N__42741),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_13_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_13_9_1 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIJ4DM1_19_LC_13_9_1  (
            .in0(N__39136),
            .in1(_gnd_net_),
            .in2(N__31085),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIIJ4DM1_0_19),
            .ltout(elapsed_time_ns_1_RNIIJ4DM1_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_13_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_13_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_13_9_2 .LUT_INIT=16'b0011001100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__39882),
            .in2(N__31082),
            .in3(N__39731),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46065),
            .ce(N__44291),
            .sr(N__45546));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_13_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_13_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_13_9_3 .LUT_INIT=16'b0000000011111010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_13_9_3  (
            .in0(N__39730),
            .in1(_gnd_net_),
            .in2(N__32675),
            .in3(N__39886),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46065),
            .ce(N__44291),
            .sr(N__45546));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_13_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_13_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_13_9_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_13_9_4  (
            .in0(N__34223),
            .in1(N__39884),
            .in2(N__34191),
            .in3(N__39732),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46065),
            .ce(N__44291),
            .sr(N__45546));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_13_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_13_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_13_9_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_13_9_5  (
            .in0(N__38976),
            .in1(N__39885),
            .in2(_gnd_net_),
            .in3(N__34000),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46065),
            .ce(N__44291),
            .sr(N__45546));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_13_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_13_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_13_9_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_13_9_6  (
            .in0(N__33998),
            .in1(N__39883),
            .in2(_gnd_net_),
            .in3(N__34051),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46065),
            .ce(N__44291),
            .sr(N__45546));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_13_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_13_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_13_9_7 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_13_9_7  (
            .in0(N__32362),
            .in1(N__33999),
            .in2(N__32579),
            .in3(N__39887),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46065),
            .ce(N__44291),
            .sr(N__45546));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_13_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_13_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_13_10_0 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_13_10_0  (
            .in0(N__32764),
            .in1(N__32771),
            .in2(N__40001),
            .in3(N__39734),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46058),
            .ce(N__39585),
            .sr(N__45549));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_13_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_13_10_1 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_13_10_1  (
            .in0(N__39873),
            .in1(N__39738),
            .in2(_gnd_net_),
            .in3(N__32823),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46058),
            .ce(N__39585),
            .sr(N__45549));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_13_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_13_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_13_10_2 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_13_10_2  (
            .in0(N__39739),
            .in1(N__39874),
            .in2(_gnd_net_),
            .in3(N__32674),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46058),
            .ce(N__39585),
            .sr(N__45549));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_13_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_13_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_13_10_5 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_13_10_5  (
            .in0(N__34007),
            .in1(N__31126),
            .in2(N__32578),
            .in3(N__38603),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46058),
            .ce(N__39585),
            .sr(N__45549));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_13_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_13_10_6 .LUT_INIT=16'b0001000000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_13_10_6  (
            .in0(N__32763),
            .in1(N__34192),
            .in2(N__39200),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_13_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_13_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__33209),
            .in2(N__34121),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_13_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_13_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_13_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_13_11_1  (
            .in0(N__39587),
            .in1(N__34072),
            .in2(_gnd_net_),
            .in3(N__31154),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__46051),
            .ce(),
            .sr(N__45554));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_13_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_13_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_13_11_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_13_11_2  (
            .in0(N__39551),
            .in1(N__34463),
            .in2(N__33167),
            .in3(N__31151),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__46051),
            .ce(),
            .sr(N__45554));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_13_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_13_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_13_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_13_11_3  (
            .in0(N__39588),
            .in1(N__34426),
            .in2(_gnd_net_),
            .in3(N__31148),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__46051),
            .ce(),
            .sr(N__45554));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_13_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_13_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_13_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_13_11_4  (
            .in0(N__39552),
            .in1(N__34403),
            .in2(_gnd_net_),
            .in3(N__31145),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__46051),
            .ce(),
            .sr(N__45554));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_13_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_13_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_13_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_13_11_5  (
            .in0(N__39589),
            .in1(N__34366),
            .in2(_gnd_net_),
            .in3(N__31142),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__46051),
            .ce(),
            .sr(N__45554));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_13_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_13_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_13_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_13_11_6  (
            .in0(N__39553),
            .in1(N__34318),
            .in2(_gnd_net_),
            .in3(N__31139),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__46051),
            .ce(),
            .sr(N__45554));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_13_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_13_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_13_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_13_11_7  (
            .in0(N__39590),
            .in1(N__34295),
            .in2(_gnd_net_),
            .in3(N__31136),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__46051),
            .ce(),
            .sr(N__45554));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_13_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_13_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_13_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_13_12_0  (
            .in0(N__39581),
            .in1(N__34249),
            .in2(_gnd_net_),
            .in3(N__31133),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__46045),
            .ce(),
            .sr(N__45559));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_13_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_13_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_13_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_13_12_1  (
            .in0(N__39544),
            .in1(N__34708),
            .in2(_gnd_net_),
            .in3(N__31130),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__46045),
            .ce(),
            .sr(N__45559));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_13_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_13_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_13_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_13_12_2  (
            .in0(N__39578),
            .in1(N__34676),
            .in2(_gnd_net_),
            .in3(N__31181),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__46045),
            .ce(),
            .sr(N__45559));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_13_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_13_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_13_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_13_12_3  (
            .in0(N__39545),
            .in1(N__34634),
            .in2(_gnd_net_),
            .in3(N__31178),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__46045),
            .ce(),
            .sr(N__45559));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_13_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_13_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_13_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_13_12_4  (
            .in0(N__39579),
            .in1(N__34612),
            .in2(_gnd_net_),
            .in3(N__31175),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__46045),
            .ce(),
            .sr(N__45559));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_13_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_13_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_13_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_13_12_5  (
            .in0(N__39546),
            .in1(N__34585),
            .in2(_gnd_net_),
            .in3(N__31172),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__46045),
            .ce(),
            .sr(N__45559));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_13_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_13_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_13_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_13_12_6  (
            .in0(N__39580),
            .in1(N__34558),
            .in2(_gnd_net_),
            .in3(N__31169),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__46045),
            .ce(),
            .sr(N__45559));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_13_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_13_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_13_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_13_12_7  (
            .in0(N__39547),
            .in1(N__34522),
            .in2(_gnd_net_),
            .in3(N__31166),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__46045),
            .ce(),
            .sr(N__45559));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_13_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_13_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_13_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_13_13_0  (
            .in0(N__39548),
            .in1(N__34855),
            .in2(_gnd_net_),
            .in3(N__31163),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__46038),
            .ce(),
            .sr(N__45562));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_13_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_13_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_13_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_13_13_1  (
            .in0(N__39550),
            .in1(N__34819),
            .in2(_gnd_net_),
            .in3(N__31160),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__46038),
            .ce(),
            .sr(N__45562));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_13_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_13_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_13_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_13_13_2  (
            .in0(N__39549),
            .in1(N__34798),
            .in2(_gnd_net_),
            .in3(N__31157),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46038),
            .ce(),
            .sr(N__45562));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_13_6 .LUT_INIT=16'b1000101011001010;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_13_13_6  (
            .in0(N__31287),
            .in1(N__33244),
            .in2(N__33203),
            .in3(N__34772),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46038),
            .ce(),
            .sr(N__45562));
    defparam \phase_controller_inst2.state_0_LC_13_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_13_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_13_14_0 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_inst2.state_0_LC_13_14_0  (
            .in0(N__43740),
            .in1(N__31270),
            .in2(N__46247),
            .in3(N__46152),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46035),
            .ce(),
            .sr(N__45567));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_13_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_13_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_13_14_1 .LUT_INIT=16'b1010001011100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_13_14_1  (
            .in0(N__31271),
            .in1(N__43508),
            .in2(N__43583),
            .in3(N__43616),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46035),
            .ce(),
            .sr(N__45567));
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_13_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_13_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_RNI9M3O_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(N__31269),
            .in2(_gnd_net_),
            .in3(N__46151),
            .lcout(\phase_controller_inst2.time_passed_RNI9M3O ),
            .ltout(\phase_controller_inst2.time_passed_RNI9M3O_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_3_LC_13_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_13_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_13_14_3 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \phase_controller_inst2.state_3_LC_13_14_3  (
            .in0(N__41946),
            .in1(N__40513),
            .in2(N__31259),
            .in3(N__33715),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46035),
            .ce(),
            .sr(N__45567));
    defparam \phase_controller_inst1.state_4_LC_13_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_13_14_5 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_13_14_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_13_14_5  (
            .in0(N__40564),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43650),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46035),
            .ce(),
            .sr(N__45567));
    defparam \current_shift_inst.stop_timer_s1_LC_13_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_13_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_13_15_0 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_13_15_0  (
            .in0(N__31253),
            .in1(N__31195),
            .in2(N__31507),
            .in3(N__32423),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46033),
            .ce(),
            .sr(N__45573));
    defparam \current_shift_inst.timer_s1.running_LC_13_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_13_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_13_15_2 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_13_15_2  (
            .in0(N__31502),
            .in1(N__35810),
            .in2(_gnd_net_),
            .in3(N__32424),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46033),
            .ce(),
            .sr(N__45573));
    defparam \current_shift_inst.start_timer_s1_LC_13_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_13_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_13_15_3 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_13_15_3  (
            .in0(N__31194),
            .in1(N__31503),
            .in2(_gnd_net_),
            .in3(N__31255),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46033),
            .ce(),
            .sr(N__45573));
    defparam \phase_controller_inst1.S1_LC_13_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_13_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_13_15_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.S1_LC_13_15_4  (
            .in0(N__31254),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46033),
            .ce(),
            .sr(N__45573));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31448),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_13_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_13_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31401),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_13_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_13_16_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_13_16_3  (
            .in0(N__31334),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33263),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37565),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46030),
            .ce(N__41021),
            .sr(N__45578));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_13_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_13_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35381),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_13_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_13_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35336),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_13_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_13_17_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_13_17_0  (
            .in0(N__47194),
            .in1(N__33385),
            .in2(N__44054),
            .in3(N__31480),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_13_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_13_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_13_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37532),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46025),
            .ce(N__41020),
            .sr(N__45582));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31475),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_3 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_3  (
            .in0(N__33386),
            .in1(N__47195),
            .in2(N__31481),
            .in3(N__44053),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_13_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_13_17_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_13_17_4  (
            .in0(N__42192),
            .in1(N__33384),
            .in2(_gnd_net_),
            .in3(N__31476),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_13_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_13_17_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__47196),
            .in2(_gnd_net_),
            .in3(N__33553),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_13_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_13_17_6 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_13_17_6  (
            .in0(N__47197),
            .in1(_gnd_net_),
            .in2(N__33557),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_0_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_13_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_13_18_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_13_18_0  (
            .in0(N__42241),
            .in1(N__36768),
            .in2(_gnd_net_),
            .in3(N__36726),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_13_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_13_18_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_13_18_1  (
            .in0(N__46975),
            .in1(N__47325),
            .in2(N__35344),
            .in3(N__33310),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_18_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_18_2  (
            .in0(N__42239),
            .in1(N__35382),
            .in2(_gnd_net_),
            .in3(N__33339),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_13_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_13_18_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_13_18_3  (
            .in0(N__46973),
            .in1(N__47327),
            .in2(N__35200),
            .in3(N__35473),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_13_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_13_18_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_13_18_4  (
            .in0(N__42238),
            .in1(N__33367),
            .in2(_gnd_net_),
            .in3(N__35436),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_13_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_13_18_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_13_18_5  (
            .in0(N__35337),
            .in1(N__42240),
            .in2(_gnd_net_),
            .in3(N__33309),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_13_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_13_18_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_13_18_6  (
            .in0(N__47326),
            .in1(N__46976),
            .in2(N__36773),
            .in3(N__36727),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_18_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_18_7  (
            .in0(N__46974),
            .in1(N__47328),
            .in2(N__35201),
            .in3(N__35474),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_19_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_13_19_0  (
            .in0(N__44917),
            .in1(N__47335),
            .in2(N__47003),
            .in3(N__44878),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_19_1 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_19_1  (
            .in0(N__31508),
            .in1(N__35817),
            .in2(_gnd_net_),
            .in3(N__32428),
            .lcout(\current_shift_inst.timer_s1.N_167_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_13_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_13_19_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_13_19_2  (
            .in0(N__44916),
            .in1(N__47334),
            .in2(_gnd_net_),
            .in3(N__44877),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_13_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_13_19_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_13_19_3  (
            .in0(N__47333),
            .in1(N__46992),
            .in2(N__47450),
            .in3(N__47470),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_13_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_13_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44915),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_13_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_13_19_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_13_19_7  (
            .in0(N__47332),
            .in1(N__41340),
            .in2(_gnd_net_),
            .in3(N__41292),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45228),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_13_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_13_20_1 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_13_20_1  (
            .in0(N__36981),
            .in1(N__42257),
            .in2(_gnd_net_),
            .in3(N__42387),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_20_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(N__37061),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35278),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45075),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_13_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_13_20_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_13_20_6  (
            .in0(N__47336),
            .in1(N__44680),
            .in2(N__47004),
            .in3(N__44698),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_13_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_13_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_13_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_13_21_0  (
            .in0(N__32143),
            .in1(N__33816),
            .in2(_gnd_net_),
            .in3(N__31613),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_21_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__46010),
            .ce(N__32471),
            .sr(N__45606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_13_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_13_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_13_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_13_21_1  (
            .in0(N__32139),
            .in1(N__31596),
            .in2(_gnd_net_),
            .in3(N__31580),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__46010),
            .ce(N__32471),
            .sr(N__45606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_13_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_13_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_13_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_13_21_2  (
            .in0(N__32144),
            .in1(N__31573),
            .in2(_gnd_net_),
            .in3(N__31556),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__46010),
            .ce(N__32471),
            .sr(N__45606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_13_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_13_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_13_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_13_21_3  (
            .in0(N__32140),
            .in1(N__31549),
            .in2(_gnd_net_),
            .in3(N__31532),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__46010),
            .ce(N__32471),
            .sr(N__45606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_13_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_13_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_13_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_13_21_4  (
            .in0(N__32145),
            .in1(N__31525),
            .in2(_gnd_net_),
            .in3(N__31823),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__46010),
            .ce(N__32471),
            .sr(N__45606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_13_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_13_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_13_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_13_21_5  (
            .in0(N__32141),
            .in1(N__31816),
            .in2(_gnd_net_),
            .in3(N__31799),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__46010),
            .ce(N__32471),
            .sr(N__45606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_13_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_13_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_13_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_13_21_6  (
            .in0(N__32146),
            .in1(N__31796),
            .in2(_gnd_net_),
            .in3(N__31781),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__46010),
            .ce(N__32471),
            .sr(N__45606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_13_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_13_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_13_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_13_21_7  (
            .in0(N__32142),
            .in1(N__31778),
            .in2(_gnd_net_),
            .in3(N__31763),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__46010),
            .ce(N__32471),
            .sr(N__45606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_13_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_13_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_13_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_13_22_0  (
            .in0(N__32150),
            .in1(N__31752),
            .in2(_gnd_net_),
            .in3(N__31733),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_22_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__46004),
            .ce(N__32469),
            .sr(N__45620));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_13_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_13_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_13_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_13_22_1  (
            .in0(N__32162),
            .in1(N__31722),
            .in2(_gnd_net_),
            .in3(N__31703),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__46004),
            .ce(N__32469),
            .sr(N__45620));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_13_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_13_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_13_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_13_22_2  (
            .in0(N__32147),
            .in1(N__31696),
            .in2(_gnd_net_),
            .in3(N__31679),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__46004),
            .ce(N__32469),
            .sr(N__45620));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_13_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_13_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_13_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_13_22_3  (
            .in0(N__32159),
            .in1(N__31672),
            .in2(_gnd_net_),
            .in3(N__31655),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__46004),
            .ce(N__32469),
            .sr(N__45620));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_13_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_13_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_13_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_13_22_4  (
            .in0(N__32148),
            .in1(N__31648),
            .in2(_gnd_net_),
            .in3(N__31631),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__46004),
            .ce(N__32469),
            .sr(N__45620));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_13_22_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_13_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_13_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_13_22_5  (
            .in0(N__32160),
            .in1(N__32020),
            .in2(_gnd_net_),
            .in3(N__32003),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__46004),
            .ce(N__32469),
            .sr(N__45620));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_13_22_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_13_22_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_13_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_13_22_6  (
            .in0(N__32149),
            .in1(N__32000),
            .in2(_gnd_net_),
            .in3(N__31985),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__46004),
            .ce(N__32469),
            .sr(N__45620));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_13_22_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_13_22_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_13_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_13_22_7  (
            .in0(N__32161),
            .in1(N__31982),
            .in2(_gnd_net_),
            .in3(N__31967),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__46004),
            .ce(N__32469),
            .sr(N__45620));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_13_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_13_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_13_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_13_23_0  (
            .in0(N__32155),
            .in1(N__31953),
            .in2(_gnd_net_),
            .in3(N__31934),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__46001),
            .ce(N__32470),
            .sr(N__45631));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_13_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_13_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_13_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_13_23_1  (
            .in0(N__32165),
            .in1(N__31923),
            .in2(_gnd_net_),
            .in3(N__31904),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__46001),
            .ce(N__32470),
            .sr(N__45631));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_13_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_13_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_13_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_13_23_2  (
            .in0(N__32156),
            .in1(N__31893),
            .in2(_gnd_net_),
            .in3(N__31874),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__46001),
            .ce(N__32470),
            .sr(N__45631));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_13_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_13_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_13_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_13_23_3  (
            .in0(N__32166),
            .in1(N__31867),
            .in2(_gnd_net_),
            .in3(N__31850),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__46001),
            .ce(N__32470),
            .sr(N__45631));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_13_23_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_13_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_13_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_13_23_4  (
            .in0(N__32157),
            .in1(N__31843),
            .in2(_gnd_net_),
            .in3(N__31826),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__46001),
            .ce(N__32470),
            .sr(N__45631));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_13_23_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_13_23_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_13_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_13_23_5  (
            .in0(N__32167),
            .in1(N__32347),
            .in2(_gnd_net_),
            .in3(N__32330),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__46001),
            .ce(N__32470),
            .sr(N__45631));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_13_23_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_13_23_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_13_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_13_23_6  (
            .in0(N__32158),
            .in1(N__32327),
            .in2(_gnd_net_),
            .in3(N__32312),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__46001),
            .ce(N__32470),
            .sr(N__45631));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_13_23_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_13_23_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_13_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_13_23_7  (
            .in0(N__32168),
            .in1(N__32309),
            .in2(_gnd_net_),
            .in3(N__32294),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__46001),
            .ce(N__32470),
            .sr(N__45631));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_13_24_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_13_24_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_13_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_13_24_0  (
            .in0(N__32151),
            .in1(N__32283),
            .in2(_gnd_net_),
            .in3(N__32264),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__45997),
            .ce(N__32462),
            .sr(N__45636));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_13_24_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_13_24_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_13_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_13_24_1  (
            .in0(N__32163),
            .in1(N__32253),
            .in2(_gnd_net_),
            .in3(N__32234),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__45997),
            .ce(N__32462),
            .sr(N__45636));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_13_24_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_13_24_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_13_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_13_24_2  (
            .in0(N__32152),
            .in1(N__32227),
            .in2(_gnd_net_),
            .in3(N__32210),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__45997),
            .ce(N__32462),
            .sr(N__45636));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_13_24_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_13_24_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_13_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_13_24_3  (
            .in0(N__32164),
            .in1(N__32203),
            .in2(_gnd_net_),
            .in3(N__32186),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__45997),
            .ce(N__32462),
            .sr(N__45636));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_13_24_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_13_24_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_13_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_13_24_4  (
            .in0(N__32153),
            .in1(N__32183),
            .in2(_gnd_net_),
            .in3(N__32171),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__45997),
            .ce(N__32462),
            .sr(N__45636));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_13_24_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_13_24_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_13_24_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_13_24_5  (
            .in0(N__32036),
            .in1(N__32154),
            .in2(_gnd_net_),
            .in3(N__32039),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45997),
            .ce(N__32462),
            .sr(N__45636));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_26_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_26_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_26_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_13_26_1  (
            .in0(_gnd_net_),
            .in1(N__35818),
            .in2(_gnd_net_),
            .in3(N__32429),
            .lcout(\current_shift_inst.timer_s1.N_166_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_14_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_14_7_0 .LUT_INIT=16'b1010111011111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_14_7_0  (
            .in0(N__42733),
            .in1(N__32610),
            .in2(N__43172),
            .in3(N__38657),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_14_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_14_7_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPFL2M1_1_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32393),
            .in3(N__39133),
            .lcout(elapsed_time_ns_1_RNIPFL2M1_0_1),
            .ltout(elapsed_time_ns_1_RNIPFL2M1_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_14_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_14_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_14_7_2 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_14_7_2  (
            .in0(N__32551),
            .in1(N__32596),
            .in2(N__32390),
            .in3(N__32618),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46084),
            .ce(N__39598),
            .sr(N__45531));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_14_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_14_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_14_7_3 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_14_7_3  (
            .in0(N__33992),
            .in1(N__39894),
            .in2(N__32387),
            .in3(N__32559),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46084),
            .ce(N__39598),
            .sr(N__45531));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_14_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_14_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_14_7_4 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_14_7_4  (
            .in0(N__39891),
            .in1(N__32363),
            .in2(N__32574),
            .in3(N__33993),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46084),
            .ce(N__39598),
            .sr(N__45531));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_14_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_14_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_14_7_5 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_14_7_5  (
            .in0(N__33991),
            .in1(N__39893),
            .in2(N__32495),
            .in3(N__32558),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46084),
            .ce(N__39598),
            .sr(N__45531));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_14_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_14_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_14_7_6 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_14_7_6  (
            .in0(N__39892),
            .in1(N__39370),
            .in2(N__32575),
            .in3(N__33994),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46084),
            .ce(N__39598),
            .sr(N__45531));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_14_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_14_8_0 .LUT_INIT=16'b1111101111111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_14_8_0  (
            .in0(N__39017),
            .in1(N__43156),
            .in2(N__42745),
            .in3(N__32753),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_14_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_14_8_1 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_14_8_1  (
            .in0(N__42824),
            .in1(N__42971),
            .in2(N__43169),
            .in3(N__34169),
            .lcout(elapsed_time_ns_1_RNIUCHF91_0_15),
            .ltout(elapsed_time_ns_1_RNIUCHF91_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_14_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_14_8_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(N__40080),
            .in2(N__32636),
            .in3(N__32754),
            .lcout(\phase_controller_inst1.stoper_tr.N_251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_14_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_14_8_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1OL2M1_9_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__32633),
            .in2(_gnd_net_),
            .in3(N__39137),
            .lcout(elapsed_time_ns_1_RNI1OL2M1_0_9),
            .ltout(elapsed_time_ns_1_RNI1OL2M1_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_14_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_14_8_4 .LUT_INIT=16'b0011111100110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(N__40081),
            .in2(N__32627),
            .in3(N__39199),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.N_211_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_14_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_14_8_5 .LUT_INIT=16'b0000000010111010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_14_8_5  (
            .in0(N__34220),
            .in1(N__34170),
            .in2(N__32624),
            .in3(N__39677),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_14_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_14_8_6 .LUT_INIT=16'b1111111100110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(N__32611),
            .in2(N__32621),
            .in3(N__39890),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_14_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_14_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_14_8_7 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_14_8_7  (
            .in0(N__32612),
            .in1(N__32597),
            .in2(N__32582),
            .in3(N__32567),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46077),
            .ce(N__44294),
            .sr(N__45537));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_14_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_14_9_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_14_9_0  (
            .in0(N__32684),
            .in1(N__39918),
            .in2(N__32795),
            .in3(N__34026),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_14_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_14_9_1 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_14_9_1  (
            .in0(N__43146),
            .in1(N__32484),
            .in2(N__42994),
            .in3(N__35867),
            .lcout(elapsed_time_ns_1_RNICG2591_0_4),
            .ltout(elapsed_time_ns_1_RNICG2591_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_14_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_14_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_14_9_2  (
            .in0(N__32668),
            .in1(N__32822),
            .in2(N__32687),
            .in3(N__39356),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_14_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_14_9_3 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_14_9_3  (
            .in0(N__43148),
            .in1(N__36365),
            .in2(N__42746),
            .in3(N__32670),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_14_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_14_9_4 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFG4DM1_16_LC_14_9_4  (
            .in0(N__39135),
            .in1(_gnd_net_),
            .in2(N__32678),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIFG4DM1_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_14_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_14_9_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGH4DM1_17_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__32645),
            .in2(_gnd_net_),
            .in3(N__39134),
            .lcout(elapsed_time_ns_1_RNIGH4DM1_0_17),
            .ltout(elapsed_time_ns_1_RNIGH4DM1_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_14_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_14_9_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_14_9_6  (
            .in0(N__32669),
            .in1(N__39917),
            .in2(N__32648),
            .in3(N__34025),
            .lcout(\phase_controller_inst1.stoper_tr.N_214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_14_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_14_9_7 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_14_9_7  (
            .in0(N__43147),
            .in1(N__34052),
            .in2(N__42995),
            .in3(N__39044),
            .lcout(elapsed_time_ns_1_RNIGK2591_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_14_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_14_10_0 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_14_10_0  (
            .in0(N__36316),
            .in1(N__42735),
            .in2(N__32830),
            .in3(N__43157),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_10_1 .LUT_INIT=16'b1111111010101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_14_10_1  (
            .in0(N__42736),
            .in1(N__34027),
            .in2(N__43171),
            .in3(N__36257),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_14_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_14_10_2 .LUT_INIT=16'b0011000000110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHI4DM1_18_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(N__39140),
            .in2(N__32639),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIHI4DM1_0_18),
            .ltout(elapsed_time_ns_1_RNIHI4DM1_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_14_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_14_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_14_10_3 .LUT_INIT=16'b0000000011111010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_14_10_3  (
            .in0(N__39736),
            .in1(_gnd_net_),
            .in2(N__32834),
            .in3(N__39860),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46066),
            .ce(N__44289),
            .sr(N__45547));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_14_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_14_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_14_10_4 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_14_10_4  (
            .in0(N__39859),
            .in1(_gnd_net_),
            .in2(N__32831),
            .in3(N__39737),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46066),
            .ce(N__44289),
            .sr(N__45547));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_14_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_14_10_5 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_14_10_5  (
            .in0(N__43430),
            .in1(N__42990),
            .in2(N__43170),
            .in3(N__39858),
            .lcout(elapsed_time_ns_1_RNISCJF91_0_31),
            .ltout(elapsed_time_ns_1_RNISCJF91_0_31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_14_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_14_10_6 .LUT_INIT=16'b1111000011111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_14_10_6  (
            .in0(N__32801),
            .in1(N__32794),
            .in2(N__32774),
            .in3(N__39735),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_14_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_14_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_14_10_7 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_14_10_7  (
            .in0(N__32765),
            .in1(N__39733),
            .in2(N__32738),
            .in3(N__39993),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46066),
            .ce(N__44289),
            .sr(N__45547));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_14_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_14_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_14_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32730),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46059),
            .ce(),
            .sr(N__45550));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_11_5 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_11_5  (
            .in0(N__33199),
            .in1(N__33179),
            .in2(N__34120),
            .in3(N__39586),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46059),
            .ce(),
            .sr(N__45550));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_14_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_14_12_1 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_14_12_1  (
            .in0(N__33232),
            .in1(N__32695),
            .in2(_gnd_net_),
            .in3(N__32734),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(\phase_controller_inst1.stoper_tr.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_LC_14_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_14_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_14_12_2 .LUT_INIT=16'b1000101011111010;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_14_12_2  (
            .in0(N__32696),
            .in1(N__34771),
            .in2(N__32699),
            .in3(N__33234),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46052),
            .ce(),
            .sr(N__45555));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIJPMR_LC_14_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIJPMR_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIJPMR_LC_14_12_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIJPMR_LC_14_12_3  (
            .in0(N__33233),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34767),
            .lcout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_12_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33212),
            .in3(N__33197),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIP6N32_LC_14_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIP6N32_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIP6N32_LC_14_12_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIP6N32_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(N__33198),
            .in2(_gnd_net_),
            .in3(N__33178),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_19_c_RNIP6NZ0Z32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_14_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_14_13_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_14_13_0  (
            .in0(N__46613),
            .in1(N__47180),
            .in2(N__41353),
            .in3(N__41302),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_14_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_14_13_3 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_14_13_3  (
            .in0(N__47177),
            .in1(N__42395),
            .in2(N__36986),
            .in3(N__46617),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_14_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_14_13_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_14_13_4  (
            .in0(N__46618),
            .in1(N__47178),
            .in2(N__35294),
            .in3(N__35245),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37079),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_14_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_14_13_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_14_13_6  (
            .in0(N__35519),
            .in1(N__47179),
            .in2(N__46802),
            .in3(N__35135),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_14_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_14_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33143),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_14_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_14_14_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_14_14_1  (
            .in0(N__47046),
            .in1(N__47109),
            .in2(_gnd_net_),
            .in3(N__46389),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41053),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46039),
            .ce(N__41022),
            .sr(N__45563));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_14_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_14_14_3  (
            .in0(N__46605),
            .in1(N__47105),
            .in2(N__35441),
            .in3(N__33373),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_14_4 .LUT_INIT=16'b1010001110100011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_14_14_4  (
            .in0(N__33374),
            .in1(N__35437),
            .in2(N__47193),
            .in3(N__46606),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_14_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_14_14_5 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_14_14_5  (
            .in0(N__33277),
            .in1(N__33290),
            .in2(_gnd_net_),
            .in3(N__47104),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_14_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_14_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33421),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_14_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_14_14_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__47103),
            .in2(N__33284),
            .in3(N__33276),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_14_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_14_15_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_14_15_0  (
            .in0(N__45080),
            .in1(N__47204),
            .in2(N__46806),
            .in3(N__45036),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_15_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_15_1  (
            .in0(N__47198),
            .in1(N__42044),
            .in2(N__46805),
            .in3(N__42010),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_14_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_14_15_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_14_15_2  (
            .in0(N__46632),
            .in1(N__47199),
            .in2(N__35399),
            .in3(N__33344),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_14_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_14_15_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_14_15_3  (
            .in0(N__47205),
            .in1(N__35515),
            .in2(N__46804),
            .in3(N__35134),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_14_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_14_15_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_14_15_4  (
            .in0(N__46633),
            .in1(N__47200),
            .in2(N__35348),
            .in3(N__33314),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_14_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_14_15_5 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_14_15_5  (
            .in0(N__47203),
            .in1(N__46628),
            .in2(N__42445),
            .in3(N__42487),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_14_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_14_15_6 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_14_15_6  (
            .in0(N__35246),
            .in1(N__47201),
            .in2(N__46807),
            .in3(N__35293),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_14_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_14_15_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_14_15_7  (
            .in0(N__47202),
            .in1(N__35572),
            .in2(N__46803),
            .in3(N__35114),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_16_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_16_0  (
            .in0(N__47223),
            .in1(N__46879),
            .in2(N__35573),
            .in3(N__35113),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_14_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_14_16_1 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_14_16_1  (
            .in0(N__46881),
            .in1(N__47225),
            .in2(N__41749),
            .in3(N__41785),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_14_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_14_16_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_14_16_2  (
            .in0(N__47226),
            .in1(N__46882),
            .in2(N__45239),
            .in3(N__45190),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_16_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_16_3  (
            .in0(N__46883),
            .in1(N__47227),
            .in2(N__41231),
            .in3(N__41261),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_14_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_14_16_4 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_14_16_4  (
            .in0(N__47222),
            .in1(N__46885),
            .in2(N__42081),
            .in3(N__42121),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_14_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_14_16_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_14_16_5  (
            .in0(N__46880),
            .in1(N__47224),
            .in2(N__45154),
            .in3(N__45112),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_14_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_14_16_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_14_16_6  (
            .in0(N__47221),
            .in1(N__46884),
            .in2(N__35395),
            .in3(N__33340),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_16_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_14_16_7  (
            .in0(N__46878),
            .in1(N__47228),
            .in2(N__42341),
            .in3(N__42292),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_14_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_14_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__33431),
            .in2(N__33417),
            .in3(N__33410),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_14_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_14_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__35150),
            .in2(_gnd_net_),
            .in3(N__33356),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_14_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_14_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__35252),
            .in2(_gnd_net_),
            .in3(N__33353),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_14_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_14_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__33350),
            .in2(_gnd_net_),
            .in3(N__33323),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_14_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_14_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__33320),
            .in2(_gnd_net_),
            .in3(N__33296),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_14_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_14_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__35210),
            .in2(_gnd_net_),
            .in3(N__33293),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_14_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_14_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__42353),
            .in2(_gnd_net_),
            .in3(N__33482),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_14_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_14_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__33542),
            .in2(_gnd_net_),
            .in3(N__33479),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_14_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_14_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__33476),
            .in2(_gnd_net_),
            .in3(N__33461),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_14_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_14_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__33632),
            .in2(_gnd_net_),
            .in3(N__33458),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_14_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_14_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__33653),
            .in2(_gnd_net_),
            .in3(N__33455),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_14_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_14_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__33527),
            .in2(_gnd_net_),
            .in3(N__33452),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_14_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_14_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__33449),
            .in2(_gnd_net_),
            .in3(N__33440),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_14_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_14_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__33608),
            .in2(_gnd_net_),
            .in3(N__33437),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_14_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_14_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__33641),
            .in2(_gnd_net_),
            .in3(N__33434),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_14_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_14_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__33518),
            .in2(_gnd_net_),
            .in3(N__33509),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_14_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_14_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__33533),
            .in2(_gnd_net_),
            .in3(N__33506),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_14_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_14_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__33617),
            .in2(_gnd_net_),
            .in3(N__33503),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_14_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_14_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__33662),
            .in2(_gnd_net_),
            .in3(N__33500),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_14_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_14_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__33599),
            .in2(_gnd_net_),
            .in3(N__33497),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_14_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_14_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__33590),
            .in2(_gnd_net_),
            .in3(N__33494),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_14_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_14_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__37577),
            .in2(_gnd_net_),
            .in3(N__33491),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_14_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_14_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__33860),
            .in2(_gnd_net_),
            .in3(N__33488),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_14_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_14_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__33842),
            .in2(_gnd_net_),
            .in3(N__33485),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_14_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_14_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__33623),
            .in2(_gnd_net_),
            .in3(N__33581),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_14_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_14_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__33851),
            .in2(_gnd_net_),
            .in3(N__33578),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_14_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_14_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__33833),
            .in2(_gnd_net_),
            .in3(N__33575),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_14_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_14_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__35837),
            .in2(_gnd_net_),
            .in3(N__33572),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_14_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_14_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__33569),
            .in2(_gnd_net_),
            .in3(N__33563),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_14_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_14_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33560),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42101),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41211),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42467),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47429),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45131),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_14_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_14_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35499),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35550),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44978),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_14_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_14_21_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_14_21_6  (
            .in0(N__35457),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41768),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_14_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_14_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_14_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44663),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41101),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_14_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44756),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_14_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_14_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_14_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41321),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_14_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_14_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44840),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47027),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_14_23_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_14_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_14_23_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_14_23_0  (
            .in0(_gnd_net_),
            .in1(N__33824),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46005),
            .ce(N__33772),
            .sr(N__45621));
    defparam \phase_controller_inst2.start_timer_hc_LC_14_24_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_14_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_14_24_2 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_14_24_2  (
            .in0(N__43677),
            .in1(N__35825),
            .in2(N__33749),
            .in3(N__33683),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46002),
            .ce(),
            .sr(N__45632));
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_14_25_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_14_25_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_14_25_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_1_LC_14_25_7  (
            .in0(_gnd_net_),
            .in1(N__41962),
            .in2(_gnd_net_),
            .in3(N__33714),
            .lcout(\phase_controller_inst2.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_15_4_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_15_4_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_15_4_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_15_4_5  (
            .in0(_gnd_net_),
            .in1(N__35741),
            .in2(_gnd_net_),
            .in3(N__46355),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_434_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_15_5_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_15_5_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_15_5_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_15_5_0  (
            .in0(N__35696),
            .in1(N__38715),
            .in2(_gnd_net_),
            .in3(N__33665),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_5_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__46102),
            .ce(N__35785),
            .sr(N__45519));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_15_5_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_15_5_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_15_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_15_5_1  (
            .in0(N__35683),
            .in1(N__35886),
            .in2(_gnd_net_),
            .in3(N__33887),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__46102),
            .ce(N__35785),
            .sr(N__45519));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_15_5_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_15_5_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_15_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_15_5_2  (
            .in0(N__35697),
            .in1(N__36144),
            .in2(_gnd_net_),
            .in3(N__33884),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__46102),
            .ce(N__35785),
            .sr(N__45519));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_15_5_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_15_5_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_15_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_15_5_3  (
            .in0(N__35684),
            .in1(N__36123),
            .in2(_gnd_net_),
            .in3(N__33881),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__46102),
            .ce(N__35785),
            .sr(N__45519));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_15_5_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_15_5_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_15_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_15_5_4  (
            .in0(N__35698),
            .in1(N__36099),
            .in2(_gnd_net_),
            .in3(N__33878),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__46102),
            .ce(N__35785),
            .sr(N__45519));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_15_5_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_15_5_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_15_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_15_5_5  (
            .in0(N__35685),
            .in1(N__36072),
            .in2(_gnd_net_),
            .in3(N__33875),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__46102),
            .ce(N__35785),
            .sr(N__45519));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_15_5_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_15_5_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_15_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_15_5_6  (
            .in0(N__35699),
            .in1(N__36042),
            .in2(_gnd_net_),
            .in3(N__33872),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__46102),
            .ce(N__35785),
            .sr(N__45519));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_15_5_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_15_5_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_15_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_15_5_7  (
            .in0(N__35686),
            .in1(N__36015),
            .in2(_gnd_net_),
            .in3(N__33869),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__46102),
            .ce(N__35785),
            .sr(N__45519));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_15_6_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_15_6_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_15_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_15_6_0  (
            .in0(N__35717),
            .in1(N__35988),
            .in2(_gnd_net_),
            .in3(N__33866),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_15_6_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__46097),
            .ce(N__35777),
            .sr(N__45526));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_15_6_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_15_6_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_15_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_15_6_1  (
            .in0(N__35674),
            .in1(N__35955),
            .in2(_gnd_net_),
            .in3(N__33863),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__46097),
            .ce(N__35777),
            .sr(N__45526));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_15_6_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_15_6_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_15_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_15_6_2  (
            .in0(N__35714),
            .in1(N__36456),
            .in2(_gnd_net_),
            .in3(N__33914),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__46097),
            .ce(N__35777),
            .sr(N__45526));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_15_6_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_15_6_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_15_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_15_6_3  (
            .in0(N__35671),
            .in1(N__36432),
            .in2(_gnd_net_),
            .in3(N__33911),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__46097),
            .ce(N__35777),
            .sr(N__45526));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_15_6_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_15_6_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_15_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_15_6_4  (
            .in0(N__35715),
            .in1(N__36405),
            .in2(_gnd_net_),
            .in3(N__33908),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__46097),
            .ce(N__35777),
            .sr(N__45526));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_15_6_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_15_6_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_15_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_15_6_5  (
            .in0(N__35672),
            .in1(N__36381),
            .in2(_gnd_net_),
            .in3(N__33905),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__46097),
            .ce(N__35777),
            .sr(N__45526));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_15_6_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_15_6_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_15_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_15_6_6  (
            .in0(N__35716),
            .in1(N__36333),
            .in2(_gnd_net_),
            .in3(N__33902),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__46097),
            .ce(N__35777),
            .sr(N__45526));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_15_6_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_15_6_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_15_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_15_6_7  (
            .in0(N__35673),
            .in1(N__36271),
            .in2(_gnd_net_),
            .in3(N__33899),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__46097),
            .ce(N__35777),
            .sr(N__45526));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_15_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_15_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_15_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_15_7_0  (
            .in0(N__35675),
            .in1(N__36225),
            .in2(_gnd_net_),
            .in3(N__33896),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_15_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__46092),
            .ce(N__35786),
            .sr(N__45528));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_15_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_15_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_15_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_15_7_1  (
            .in0(N__35679),
            .in1(N__36168),
            .in2(_gnd_net_),
            .in3(N__33893),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__46092),
            .ce(N__35786),
            .sr(N__45528));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_15_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_15_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_15_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_15_7_2  (
            .in0(N__35676),
            .in1(N__36711),
            .in2(_gnd_net_),
            .in3(N__33890),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__46092),
            .ce(N__35786),
            .sr(N__45528));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_15_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_15_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_15_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_15_7_3  (
            .in0(N__35680),
            .in1(N__36690),
            .in2(_gnd_net_),
            .in3(N__33941),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__46092),
            .ce(N__35786),
            .sr(N__45528));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_15_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_15_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_15_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_15_7_4  (
            .in0(N__35677),
            .in1(N__36666),
            .in2(_gnd_net_),
            .in3(N__33938),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__46092),
            .ce(N__35786),
            .sr(N__45528));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_15_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_15_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_15_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_15_7_5  (
            .in0(N__35681),
            .in1(N__36639),
            .in2(_gnd_net_),
            .in3(N__33935),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__46092),
            .ce(N__35786),
            .sr(N__45528));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_15_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_15_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_15_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_15_7_6  (
            .in0(N__35678),
            .in1(N__36609),
            .in2(_gnd_net_),
            .in3(N__33932),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__46092),
            .ce(N__35786),
            .sr(N__45528));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_15_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_15_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_15_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_15_7_7  (
            .in0(N__35682),
            .in1(N__36582),
            .in2(_gnd_net_),
            .in3(N__33929),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__46092),
            .ce(N__35786),
            .sr(N__45528));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_15_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_15_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_15_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_15_8_0  (
            .in0(N__35718),
            .in1(N__36555),
            .in2(_gnd_net_),
            .in3(N__33926),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__46085),
            .ce(N__35784),
            .sr(N__45532));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_15_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_15_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_15_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_15_8_1  (
            .in0(N__35722),
            .in1(N__36522),
            .in2(_gnd_net_),
            .in3(N__33923),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__46085),
            .ce(N__35784),
            .sr(N__45532));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_15_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_15_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_15_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_15_8_2  (
            .in0(N__35719),
            .in1(N__36498),
            .in2(_gnd_net_),
            .in3(N__33920),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__46085),
            .ce(N__35784),
            .sr(N__45532));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_15_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_15_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_15_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_15_8_3  (
            .in0(N__35723),
            .in1(N__36834),
            .in2(_gnd_net_),
            .in3(N__33917),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__46085),
            .ce(N__35784),
            .sr(N__45532));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_15_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_15_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_15_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_15_8_4  (
            .in0(N__35720),
            .in1(N__36475),
            .in2(_gnd_net_),
            .in3(N__34058),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__46085),
            .ce(N__35784),
            .sr(N__45532));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_15_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_15_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_15_8_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_15_8_5  (
            .in0(N__36853),
            .in1(N__35721),
            .in2(_gnd_net_),
            .in3(N__34055),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46085),
            .ce(N__35784),
            .sr(N__45532));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_15_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_15_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_15_9_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_15_9_0  (
            .in0(N__39876),
            .in1(N__34050),
            .in2(_gnd_net_),
            .in3(N__34003),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46078),
            .ce(N__39599),
            .sr(N__45538));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_15_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_15_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_15_9_1 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_15_9_1  (
            .in0(N__34028),
            .in1(N__39879),
            .in2(_gnd_net_),
            .in3(N__39751),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46078),
            .ce(N__39599),
            .sr(N__45538));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_15_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_15_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_15_9_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_15_9_2  (
            .in0(N__39875),
            .in1(N__38977),
            .in2(_gnd_net_),
            .in3(N__34002),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46078),
            .ce(N__39599),
            .sr(N__45538));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_9_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_15_9_3  (
            .in0(N__39990),
            .in1(N__39880),
            .in2(N__39236),
            .in3(N__39752),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46078),
            .ce(N__39599),
            .sr(N__45538));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_9_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_15_9_4  (
            .in0(N__39877),
            .in1(N__39991),
            .in2(N__39754),
            .in3(N__43336),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46078),
            .ce(N__39599),
            .sr(N__45538));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_9_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_15_9_6  (
            .in0(N__39878),
            .in1(N__39992),
            .in2(N__39755),
            .in3(N__39262),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46078),
            .ce(N__39599),
            .sr(N__45538));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_9_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_15_9_7  (
            .in0(N__34222),
            .in1(N__39881),
            .in2(N__34190),
            .in3(N__39753),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46078),
            .ce(N__39599),
            .sr(N__45538));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_15_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_15_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_15_10_0 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_15_10_0  (
            .in0(N__39863),
            .in1(N__40076),
            .in2(N__40000),
            .in3(N__39744),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46071),
            .ce(N__44292),
            .sr(N__45542));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_15_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_15_10_1 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_15_10_1  (
            .in0(N__40075),
            .in1(N__43167),
            .in2(N__42789),
            .in3(N__42734),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_15_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_15_10_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDE4DM1_14_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34226),
            .in3(N__39139),
            .lcout(elapsed_time_ns_1_RNIDE4DM1_0_14),
            .ltout(elapsed_time_ns_1_RNIDE4DM1_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_15_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_15_10_3 .LUT_INIT=16'b0011001100110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__34221),
            .in2(N__34199),
            .in3(N__34196),
            .lcout(\phase_controller_inst1.stoper_tr.N_241 ),
            .ltout(\phase_controller_inst1.stoper_tr.N_241_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_15_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_15_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_15_10_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_15_10_4  (
            .in0(N__39861),
            .in1(N__43337),
            .in2(N__34136),
            .in3(N__39742),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46071),
            .ce(N__44292),
            .sr(N__45542));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_15_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_15_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_15_10_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_15_10_5  (
            .in0(N__39740),
            .in1(N__39864),
            .in2(N__39266),
            .in3(N__39988),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46071),
            .ce(N__44292),
            .sr(N__45542));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_15_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_15_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_15_10_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_15_10_6  (
            .in0(N__39862),
            .in1(N__39232),
            .in2(N__39999),
            .in3(N__39743),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46071),
            .ce(N__44292),
            .sr(N__45542));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_15_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_15_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_15_10_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_15_10_7  (
            .in0(N__39741),
            .in1(N__39865),
            .in2(N__40028),
            .in3(N__39989),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46071),
            .ce(N__44292),
            .sr(N__45542));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_1_c_inv_LC_15_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_1_c_inv_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_1_c_inv_LC_15_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_1_c_inv_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__34133),
            .in2(N__34094),
            .in3(N__34110),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_2_c_inv_LC_15_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_2_c_inv_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_2_c_inv_LC_15_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_2_c_inv_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__34085),
            .in2(N__34487),
            .in3(N__34073),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_3_c_inv_LC_15_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_3_c_inv_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_3_c_inv_LC_15_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_3_c_inv_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__34475),
            .in2(N__34448),
            .in3(N__34462),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_4_c_inv_LC_15_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_4_c_inv_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_4_c_inv_LC_15_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_4_c_inv_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__34439),
            .in2(N__34412),
            .in3(N__34427),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_5_c_inv_LC_15_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_5_c_inv_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_5_c_inv_LC_15_11_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_5_c_inv_LC_15_11_4  (
            .in0(N__34402),
            .in1(N__34388),
            .in2(N__34376),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_6_c_inv_LC_15_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_6_c_inv_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_6_c_inv_LC_15_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_6_c_inv_LC_15_11_5  (
            .in0(N__34367),
            .in1(N__34352),
            .in2(N__34340),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_7_c_inv_LC_15_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_7_c_inv_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_7_c_inv_LC_15_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_7_c_inv_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__34328),
            .in2(N__34304),
            .in3(N__34319),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_8_c_inv_LC_15_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_8_c_inv_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_8_c_inv_LC_15_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_8_c_inv_LC_15_11_7  (
            .in0(N__34294),
            .in1(N__34280),
            .in2(N__34271),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_9_c_inv_LC_15_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_9_c_inv_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_9_c_inv_LC_15_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_9_c_inv_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__34262),
            .in2(N__34235),
            .in3(N__34250),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_10_c_inv_LC_15_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_10_c_inv_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_10_c_inv_LC_15_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_10_c_inv_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__34718),
            .in2(N__34694),
            .in3(N__34709),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_11_c_inv_LC_15_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_11_c_inv_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_11_c_inv_LC_15_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_11_c_inv_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__34685),
            .in2(N__34661),
            .in3(N__34675),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_12_c_inv_LC_15_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_12_c_inv_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_12_c_inv_LC_15_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_12_c_inv_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(N__34619),
            .in2(N__34649),
            .in3(N__34633),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_13_c_inv_LC_15_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_13_c_inv_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_13_c_inv_LC_15_12_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_13_c_inv_LC_15_12_4  (
            .in0(N__34613),
            .in1(N__39938),
            .in2(N__34598),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_14_c_inv_LC_15_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_14_c_inv_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_14_c_inv_LC_15_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_14_c_inv_LC_15_12_5  (
            .in0(N__34586),
            .in1(N__40052),
            .in2(N__34571),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_15_c_inv_LC_15_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_15_c_inv_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_15_c_inv_LC_15_12_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_15_c_inv_LC_15_12_6  (
            .in0(N__34559),
            .in1(N__34544),
            .in2(N__34532),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_16_c_inv_LC_15_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_16_c_inv_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_16_c_inv_LC_15_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_16_c_inv_LC_15_12_7  (
            .in0(N__34523),
            .in1(N__34508),
            .in2(N__34496),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_17_c_inv_LC_15_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_17_c_inv_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_17_c_inv_LC_15_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_17_c_inv_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__34868),
            .in2(N__34841),
            .in3(N__34856),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_18_c_inv_LC_15_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_18_c_inv_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_18_c_inv_LC_15_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_18_c_inv_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__34805),
            .in2(N__34832),
            .in3(N__34820),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_inv_LC_15_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_inv_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_inv_LC_15_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_19_c_inv_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__39611),
            .in2(N__34784),
            .in3(N__34799),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_15_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_15_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34775),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_15_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_15_13_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_15_13_5  (
            .in0(N__43573),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43529),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__34751),
            .in2(N__44095),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__44040),
            .in2(N__34745),
            .in3(N__37215),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_14_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_14_2  (
            .in0(N__37216),
            .in1(N__46509),
            .in2(N__34730),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__34940),
            .in2(N__46648),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(N__46513),
            .in2(N__34934),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(N__34925),
            .in2(N__46649),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__46517),
            .in2(N__34919),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(N__34904),
            .in2(N__46650),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__46554),
            .in2(N__34898),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__34889),
            .in2(N__46756),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__46558),
            .in2(N__34883),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(N__34874),
            .in2(N__46757),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__46562),
            .in2(N__35012),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(N__35003),
            .in2(N__46758),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(N__46566),
            .in2(N__34997),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(N__34988),
            .in2(N__46759),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(N__46760),
            .in2(N__34982),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(N__34973),
            .in2(N__46911),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(N__46764),
            .in2(N__34967),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_16_3  (
            .in0(_gnd_net_),
            .in1(N__34952),
            .in2(N__46912),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__46768),
            .in2(N__35090),
            .in3(N__35075),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(N__41129),
            .in2(N__46913),
            .in3(N__35072),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(N__46772),
            .in2(N__35069),
            .in3(N__35060),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(N__35219),
            .in2(N__46914),
            .in3(N__35057),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__46776),
            .in2(N__35144),
            .in3(N__35054),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__35180),
            .in2(N__46915),
            .in3(N__35051),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__46780),
            .in2(N__35048),
            .in3(N__35033),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__35030),
            .in2(N__46916),
            .in3(N__35018),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__46784),
            .in2(N__40757),
            .in3(N__35015),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__35171),
            .in2(N__46917),
            .in3(N__35159),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_15_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_15_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__46788),
            .in2(N__44539),
            .in3(N__35156),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_0_11_LC_15_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_0_11_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_0_11_LC_15_17_7 .LUT_INIT=16'b1000110100100111;
    LogicCell40 \current_shift_inst.control_input_RNO_0_11_LC_15_17_7  (
            .in0(N__40937),
            .in1(N__41138),
            .in2(N__44498),
            .in3(N__35153),
            .lcout(\current_shift_inst.control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_15_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_15_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35427),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_18_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_18_1  (
            .in0(N__41778),
            .in1(N__42248),
            .in2(_gnd_net_),
            .in3(N__41733),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_18_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_18_2  (
            .in0(N__47352),
            .in1(N__46886),
            .in2(N__44857),
            .in3(N__44811),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_18_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_18_3  (
            .in0(N__42039),
            .in1(N__42245),
            .in2(_gnd_net_),
            .in3(N__42003),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_18_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_18_4  (
            .in0(N__42249),
            .in1(N__35508),
            .in2(_gnd_net_),
            .in3(N__35127),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_15_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_15_18_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_15_18_5  (
            .in0(N__35568),
            .in1(N__42246),
            .in2(_gnd_net_),
            .in3(N__35106),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42038),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_18_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_18_7  (
            .in0(N__45141),
            .in1(N__42247),
            .in2(_gnd_net_),
            .in3(N__45105),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_15_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_15_19_0 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_15_19_0  (
            .in0(N__42250),
            .in1(N__35274),
            .in2(N__35244),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_15_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_15_19_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_15_19_1  (
            .in0(N__45224),
            .in1(N__42251),
            .in2(_gnd_net_),
            .in3(N__45183),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_19_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_19_2  (
            .in0(N__46968),
            .in1(N__47350),
            .in2(N__44776),
            .in3(N__44733),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36750),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_15_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_15_19_4 .LUT_INIT=16'b1000110110001101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_15_19_4  (
            .in0(N__42252),
            .in1(N__35193),
            .in2(N__35472),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_19_5 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_19_5  (
            .in0(N__47351),
            .in1(N__46969),
            .in2(N__44952),
            .in3(N__44986),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_19_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_19_6  (
            .in0(N__42253),
            .in1(N__47439),
            .in2(_gnd_net_),
            .in3(N__47466),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_15_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_15_19_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_15_19_7  (
            .in0(N__44679),
            .in1(N__42254),
            .in2(_gnd_net_),
            .in3(N__44697),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_20_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(N__37558),
            .in2(N__37495),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__46022),
            .ce(N__41019),
            .sr(N__45589));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(N__38113),
            .in2(N__37528),
            .in3(N__35402),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__46022),
            .ce(N__41019),
            .sr(N__45589));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(N__38089),
            .in2(N__37496),
            .in3(N__35351),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__46022),
            .ce(N__41019),
            .sr(N__45589));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(N__38065),
            .in2(N__38117),
            .in3(N__35306),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__46022),
            .ce(N__41019),
            .sr(N__45589));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_20_4  (
            .in0(_gnd_net_),
            .in1(N__38090),
            .in2(N__38041),
            .in3(N__35303),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__46022),
            .ce(N__41019),
            .sr(N__45589));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(N__38014),
            .in2(N__38069),
            .in3(N__35300),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__46022),
            .ce(N__41019),
            .sr(N__45589));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__37990),
            .in2(N__38042),
            .in3(N__35297),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__46022),
            .ce(N__41019),
            .sr(N__45589));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_20_7  (
            .in0(_gnd_net_),
            .in1(N__38015),
            .in2(N__37966),
            .in3(N__35255),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__46022),
            .ce(N__41019),
            .sr(N__45589));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(N__37936),
            .in2(N__37994),
            .in3(N__35534),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__46017),
            .ce(N__41018),
            .sr(N__45593));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__38347),
            .in2(N__37967),
            .in3(N__35531),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__46017),
            .ce(N__41018),
            .sr(N__45593));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__37937),
            .in2(N__38324),
            .in3(N__35528),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__46017),
            .ce(N__41018),
            .sr(N__45593));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__38293),
            .in2(N__38351),
            .in3(N__35525),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__46017),
            .ce(N__41018),
            .sr(N__45593));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__38323),
            .in2(N__38269),
            .in3(N__35522),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__46017),
            .ce(N__41018),
            .sr(N__45593));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__38242),
            .in2(N__38297),
            .in3(N__35483),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__46017),
            .ce(N__41018),
            .sr(N__45593));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__38218),
            .in2(N__38270),
            .in3(N__35480),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__46017),
            .ce(N__41018),
            .sr(N__45593));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__38243),
            .in2(N__38195),
            .in3(N__35477),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__46017),
            .ce(N__41018),
            .sr(N__45593));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__38161),
            .in2(N__38222),
            .in3(N__35444),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__46014),
            .ce(N__41017),
            .sr(N__45600));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(N__38137),
            .in2(N__38194),
            .in3(N__35600),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__46014),
            .ce(N__41017),
            .sr(N__45600));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__38162),
            .in2(N__38558),
            .in3(N__35597),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__46014),
            .ce(N__41017),
            .sr(N__45600));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(N__38527),
            .in2(N__38141),
            .in3(N__35594),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__46014),
            .ce(N__41017),
            .sr(N__45600));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(N__38557),
            .in2(N__38503),
            .in3(N__35591),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__46014),
            .ce(N__41017),
            .sr(N__45600));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(N__38476),
            .in2(N__38531),
            .in3(N__35588),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__46014),
            .ce(N__41017),
            .sr(N__45600));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(N__38452),
            .in2(N__38504),
            .in3(N__35585),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__46014),
            .ce(N__41017),
            .sr(N__45600));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_22_7  (
            .in0(_gnd_net_),
            .in1(N__38477),
            .in2(N__38428),
            .in3(N__35582),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__46014),
            .ce(N__41017),
            .sr(N__45600));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__38398),
            .in2(N__38456),
            .in3(N__35579),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__46011),
            .ce(N__41016),
            .sr(N__45607));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(N__38374),
            .in2(N__38429),
            .in3(N__35576),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__46011),
            .ce(N__41016),
            .sr(N__45607));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(N__38399),
            .in2(N__38933),
            .in3(N__35846),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__46011),
            .ce(N__41016),
            .sr(N__45607));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__38783),
            .in2(N__38378),
            .in3(N__35843),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__46011),
            .ce(N__41016),
            .sr(N__45607));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35840),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_15_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_15_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_15_23_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_15_23_7  (
            .in0(N__41182),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_15_24_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_15_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_15_24_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(N__41850),
            .in2(_gnd_net_),
            .in3(N__41888),
            .lcout(\phase_controller_inst2.start_timer_hc_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_25_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_25_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_25_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35819),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_16_5_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_16_5_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_16_5_0 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_16_5_0  (
            .in0(N__35744),
            .in1(N__46286),
            .in2(_gnd_net_),
            .in3(N__46351),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46107),
            .ce(),
            .sr(N__45514));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_6_0 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_6_0  (
            .in0(N__35743),
            .in1(N__46285),
            .in2(_gnd_net_),
            .in3(N__46350),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_435_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_6_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_6_7  (
            .in0(_gnd_net_),
            .in1(N__35742),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_7_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_7_0  (
            .in0(N__39063),
            .in1(N__39012),
            .in2(N__42842),
            .in3(N__42785),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_7_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_7_1  (
            .in0(N__36252),
            .in1(N__36198),
            .in2(N__36317),
            .in3(N__36363),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_7_2 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_7_2  (
            .in0(N__36199),
            .in1(N__38623),
            .in2(N__38675),
            .in3(N__36253),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_16_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_16_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_16_7_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_16_LC_16_7_3  (
            .in0(N__35930),
            .in1(N__36364),
            .in2(N__35933),
            .in3(N__38636),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_380 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_7_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_7_4  (
            .in0(_gnd_net_),
            .in1(N__35860),
            .in2(_gnd_net_),
            .in3(N__39382),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_16_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_16_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGE841_17_LC_16_7_5  (
            .in0(N__39011),
            .in1(N__36309),
            .in2(N__42790),
            .in3(N__39062),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35890),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46098),
            .ce(N__38694),
            .sr(N__45527));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_16_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_16_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_16_7_7 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_16_7_7  (
            .in0(N__43102),
            .in1(N__38674),
            .in2(N__35923),
            .in3(N__42993),
            .lcout(elapsed_time_ns_1_RNIAE2591_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_8_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(N__36145),
            .in2(N__38726),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__46093),
            .ce(N__38696),
            .sr(N__45529));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__36124),
            .in2(N__35894),
            .in3(N__35849),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__46093),
            .ce(N__38696),
            .sr(N__45529));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_8_2  (
            .in0(_gnd_net_),
            .in1(N__36146),
            .in2(N__36104),
            .in3(N__36128),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__46093),
            .ce(N__38696),
            .sr(N__45529));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_8_3  (
            .in0(_gnd_net_),
            .in1(N__36125),
            .in2(N__36077),
            .in3(N__36107),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__46093),
            .ce(N__38696),
            .sr(N__45529));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__36103),
            .in2(N__36049),
            .in3(N__36080),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__46093),
            .ce(N__38696),
            .sr(N__45529));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_8_5  (
            .in0(_gnd_net_),
            .in1(N__36076),
            .in2(N__36022),
            .in3(N__36053),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__46093),
            .ce(N__38696),
            .sr(N__45529));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(N__35989),
            .in2(N__36050),
            .in3(N__36026),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__46093),
            .ce(N__38696),
            .sr(N__45529));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(N__35956),
            .in2(N__36023),
            .in3(N__35999),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__46093),
            .ce(N__38696),
            .sr(N__45529));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_9_0  (
            .in0(_gnd_net_),
            .in1(N__36457),
            .in2(N__35996),
            .in3(N__35966),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__46086),
            .ce(N__38697),
            .sr(N__45533));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_9_1  (
            .in0(_gnd_net_),
            .in1(N__36433),
            .in2(N__35963),
            .in3(N__35936),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__46086),
            .ce(N__38697),
            .sr(N__45533));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_9_2  (
            .in0(_gnd_net_),
            .in1(N__36458),
            .in2(N__36410),
            .in3(N__36440),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__46086),
            .ce(N__38697),
            .sr(N__45533));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__36382),
            .in2(N__36437),
            .in3(N__36413),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__46086),
            .ce(N__38697),
            .sr(N__45533));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_9_4  (
            .in0(_gnd_net_),
            .in1(N__36409),
            .in2(N__36340),
            .in3(N__36386),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__46086),
            .ce(N__38697),
            .sr(N__45533));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_9_5  (
            .in0(_gnd_net_),
            .in1(N__36383),
            .in2(N__36283),
            .in3(N__36344),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__46086),
            .ce(N__38697),
            .sr(N__45533));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__36226),
            .in2(N__36341),
            .in3(N__36287),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__46086),
            .ce(N__38697),
            .sr(N__45533));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(N__36169),
            .in2(N__36284),
            .in3(N__36236),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__46086),
            .ce(N__38697),
            .sr(N__45533));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__36712),
            .in2(N__36233),
            .in3(N__36179),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__46079),
            .ce(N__38698),
            .sr(N__45539));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(N__36691),
            .in2(N__36176),
            .in3(N__36149),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__46079),
            .ce(N__38698),
            .sr(N__45539));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(N__36713),
            .in2(N__36671),
            .in3(N__36695),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__46079),
            .ce(N__38698),
            .sr(N__45539));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__36692),
            .in2(N__36644),
            .in3(N__36674),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__46079),
            .ce(N__38698),
            .sr(N__45539));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(N__36670),
            .in2(N__36616),
            .in3(N__36647),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__46079),
            .ce(N__38698),
            .sr(N__45539));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(N__36643),
            .in2(N__36589),
            .in3(N__36620),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__46079),
            .ce(N__38698),
            .sr(N__45539));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(N__36556),
            .in2(N__36617),
            .in3(N__36593),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__46079),
            .ce(N__38698),
            .sr(N__45539));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_10_7  (
            .in0(_gnd_net_),
            .in1(N__36523),
            .in2(N__36590),
            .in3(N__36566),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__46079),
            .ce(N__38698),
            .sr(N__45539));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__36499),
            .in2(N__36563),
            .in3(N__36533),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__46072),
            .ce(N__38699),
            .sr(N__45543));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__36835),
            .in2(N__36530),
            .in3(N__36503),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__46072),
            .ce(N__38699),
            .sr(N__45543));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(N__36500),
            .in2(N__36482),
            .in3(N__36461),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__46072),
            .ce(N__38699),
            .sr(N__45543));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__36854),
            .in2(N__36839),
            .in3(N__36815),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__46072),
            .ce(N__38699),
            .sr(N__45543));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36812),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46072),
            .ce(N__38699),
            .sr(N__45543));
    defparam \phase_controller_inst2.T45_LC_16_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.T45_LC_16_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T45_LC_16_12_2 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_inst2.T45_LC_16_12_2  (
            .in0(N__36802),
            .in1(N__41972),
            .in2(_gnd_net_),
            .in3(N__46168),
            .lcout(T45_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46067),
            .ce(),
            .sr(N__45548));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_16_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_16_13_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_16_13_2  (
            .in0(N__37762),
            .in1(N__36788),
            .in2(_gnd_net_),
            .in3(N__37247),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_16_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_16_13_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_16_13_3  (
            .in0(N__44078),
            .in1(_gnd_net_),
            .in2(N__36791),
            .in3(N__37763),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_16_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_16_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_16_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41057),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46060),
            .ce(N__41024),
            .sr(N__45551));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_16_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_16_14_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_16_14_0  (
            .in0(N__44459),
            .in1(N__36782),
            .in2(_gnd_net_),
            .in3(N__40928),
            .lcout(\current_shift_inst.control_input_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_16_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_16_14_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_16_14_1  (
            .in0(N__40929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.N_1572_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_16_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_16_14_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_16_14_2  (
            .in0(N__47256),
            .in1(N__36772),
            .in2(N__46800),
            .in3(N__36734),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_16_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_16_14_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_16_14_3  (
            .in0(N__40931),
            .in1(N__44630),
            .in2(_gnd_net_),
            .in3(N__37016),
            .lcout(\current_shift_inst.control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_14_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_14_4  (
            .in0(N__37007),
            .in1(N__44399),
            .in2(_gnd_net_),
            .in3(N__40930),
            .lcout(\current_shift_inst.control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_16_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_16_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37033),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_16_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_16_14_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_16_14_6  (
            .in0(N__47257),
            .in1(N__42394),
            .in2(N__46801),
            .in3(N__36985),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_16_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_16_14_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_16_14_7  (
            .in0(N__40932),
            .in1(N__44615),
            .in2(_gnd_net_),
            .in3(N__36950),
            .lcout(\current_shift_inst.control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_0_LC_16_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_0_LC_16_15_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_0_LC_16_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_0_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__36941),
            .in2(N__36934),
            .in3(N__36935),
            .lcout(\current_shift_inst.control_inputZ0Z_0 ),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\current_shift_inst.control_input_1_cry_0 ),
            .clk(N__46046),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_LC_16_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_1_LC_16_15_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_1_LC_16_15_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_1_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37292),
            .in3(N__36881),
            .lcout(\current_shift_inst.control_inputZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_0 ),
            .carryout(\current_shift_inst.control_input_1_cry_1 ),
            .clk(N__46046),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_2_LC_16_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_2_LC_16_15_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_2_LC_16_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_2_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__37253),
            .in2(_gnd_net_),
            .in3(N__36863),
            .lcout(\current_shift_inst.control_inputZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_1 ),
            .carryout(\current_shift_inst.control_input_1_cry_2 ),
            .clk(N__46046),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_3_LC_16_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_3_LC_16_15_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_3_LC_16_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_3_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(N__36860),
            .in2(_gnd_net_),
            .in3(N__37157),
            .lcout(\current_shift_inst.control_inputZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_2 ),
            .carryout(\current_shift_inst.control_input_1_cry_3 ),
            .clk(N__46046),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_4_LC_16_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_4_LC_16_15_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_4_LC_16_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_4_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__37154),
            .in2(_gnd_net_),
            .in3(N__37136),
            .lcout(\current_shift_inst.control_inputZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_3 ),
            .carryout(\current_shift_inst.control_input_1_cry_4 ),
            .clk(N__46046),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_5_LC_16_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_5_LC_16_15_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_5_LC_16_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_5_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(N__37133),
            .in2(_gnd_net_),
            .in3(N__37112),
            .lcout(\current_shift_inst.control_inputZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_4 ),
            .carryout(\current_shift_inst.control_input_1_cry_5 ),
            .clk(N__46046),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_6_LC_16_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_6_LC_16_15_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_6_LC_16_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_6_LC_16_15_6  (
            .in0(_gnd_net_),
            .in1(N__40979),
            .in2(_gnd_net_),
            .in3(N__37100),
            .lcout(\current_shift_inst.control_inputZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_5 ),
            .carryout(\current_shift_inst.control_input_1_cry_6 ),
            .clk(N__46046),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_7_LC_16_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_7_LC_16_15_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_7_LC_16_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_7_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__37277),
            .in2(_gnd_net_),
            .in3(N__37082),
            .lcout(\current_shift_inst.control_inputZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_6 ),
            .carryout(\current_shift_inst.control_input_1_cry_7 ),
            .clk(N__46046),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_8_LC_16_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_8_LC_16_16_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_8_LC_16_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_8_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(N__40958),
            .in2(_gnd_net_),
            .in3(N__37067),
            .lcout(\current_shift_inst.control_inputZ0Z_8 ),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(\current_shift_inst.control_input_1_cry_8 ),
            .clk(N__46040),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_9_LC_16_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_9_LC_16_16_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_9_LC_16_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_9_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(N__40877),
            .in2(_gnd_net_),
            .in3(N__37064),
            .lcout(\current_shift_inst.control_inputZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_8 ),
            .carryout(\current_shift_inst.control_input_1_cry_9 ),
            .clk(N__46040),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_10_LC_16_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_10_LC_16_16_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_10_LC_16_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_10_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(N__37265),
            .in2(_gnd_net_),
            .in3(N__37049),
            .lcout(\current_shift_inst.control_inputZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_9 ),
            .carryout(\current_shift_inst.control_input_1_cry_10 ),
            .clk(N__46040),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_11_LC_16_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_11_LC_16_16_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_11_LC_16_16_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.control_input_11_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(N__37046),
            .in2(_gnd_net_),
            .in3(N__37040),
            .lcout(\current_shift_inst.control_inputZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46040),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_16_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_16_16_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_16_16_4  (
            .in0(N__37298),
            .in1(N__44438),
            .in2(_gnd_net_),
            .in3(N__40933),
            .lcout(\current_shift_inst.control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_16_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_16_5  (
            .in0(N__40935),
            .in1(N__37283),
            .in2(_gnd_net_),
            .in3(N__44582),
            .lcout(\current_shift_inst.control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_16_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_16_16_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_16_16_6  (
            .in0(N__37271),
            .in1(N__44516),
            .in2(_gnd_net_),
            .in3(N__40936),
            .lcout(\current_shift_inst.control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_16_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_16_7  (
            .in0(N__40934),
            .in1(N__44411),
            .in2(_gnd_net_),
            .in3(N__37259),
            .lcout(\current_shift_inst.control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_16_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_16_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_16_17_0  (
            .in0(_gnd_net_),
            .in1(N__37240),
            .in2(N__37223),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_16_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_16_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(N__37817),
            .in2(N__37202),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_16_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_16_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(N__37190),
            .in2(N__37880),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_16_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_16_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(N__37821),
            .in2(N__37178),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_16_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_16_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(N__37373),
            .in2(N__37881),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_16_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_16_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(N__37825),
            .in2(N__37361),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_16_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_16_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(N__37346),
            .in2(N__37882),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_16_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_16_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(N__37829),
            .in2(N__37334),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_16_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_16_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_16_18_0  (
            .in0(_gnd_net_),
            .in1(N__37842),
            .in2(N__42056),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_16_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_16_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(N__37319),
            .in2(N__37886),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_16_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_16_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(N__37830),
            .in2(N__37313),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_16_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_16_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_16_18_3  (
            .in0(_gnd_net_),
            .in1(N__37304),
            .in2(N__37883),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_16_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_16_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(N__37834),
            .in2(N__42410),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_16_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_16_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_16_18_5  (
            .in0(_gnd_net_),
            .in1(N__37604),
            .in2(N__37884),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_16_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_16_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_16_18_6  (
            .in0(_gnd_net_),
            .in1(N__37838),
            .in2(N__37421),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_16_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_16_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(N__37412),
            .in2(N__37885),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_16_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_16_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__37887),
            .in2(N__37406),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_16_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_16_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__41276),
            .in2(N__37912),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_16_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_16_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__37891),
            .in2(N__37397),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_16_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_16_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__37388),
            .in2(N__37913),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_16_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_16_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__37895),
            .in2(N__37382),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_16_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_16_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(N__37897),
            .in2(N__41069),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_16_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_16_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(N__37896),
            .in2(N__42266),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_16_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_16_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_16_19_7  (
            .in0(_gnd_net_),
            .in1(N__37898),
            .in2(N__41270),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_16_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_16_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__37899),
            .in2(N__37595),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_20_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_16_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_16_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(N__37583),
            .in2(N__37914),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_16_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_16_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(N__37903),
            .in2(N__37466),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_16_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_16_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(N__37448),
            .in2(N__37915),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_16_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_16_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(N__37907),
            .in2(N__41150),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_16_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_16_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_16_20_5  (
            .in0(_gnd_net_),
            .in1(N__37433),
            .in2(N__37916),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_16_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_16_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(N__37911),
            .in2(N__37622),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_20_7  (
            .in0(_gnd_net_),
            .in1(N__47369),
            .in2(_gnd_net_),
            .in3(N__37607),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_21_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_21_0  (
            .in0(N__42255),
            .in1(N__45060),
            .in2(_gnd_net_),
            .in3(N__45037),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_21_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_21_1  (
            .in0(N__42256),
            .in1(N__44841),
            .in2(_gnd_net_),
            .in3(N__44818),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_21_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_21_2  (
            .in0(N__47368),
            .in1(N__44979),
            .in2(_gnd_net_),
            .in3(N__44953),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42311),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_16_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_16_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_16_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_16_22_0  (
            .in0(N__38909),
            .in1(N__37554),
            .in2(_gnd_net_),
            .in3(N__37535),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_16_22_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__46018),
            .ce(N__38750),
            .sr(N__45594));
    defparam \current_shift_inst.timer_s1.counter_1_LC_16_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_16_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_16_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_16_22_1  (
            .in0(N__38905),
            .in1(N__37518),
            .in2(_gnd_net_),
            .in3(N__37499),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__46018),
            .ce(N__38750),
            .sr(N__45594));
    defparam \current_shift_inst.timer_s1.counter_2_LC_16_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_16_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_16_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_16_22_2  (
            .in0(N__38910),
            .in1(N__37483),
            .in2(_gnd_net_),
            .in3(N__37469),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__46018),
            .ce(N__38750),
            .sr(N__45594));
    defparam \current_shift_inst.timer_s1.counter_3_LC_16_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_16_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_16_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_16_22_3  (
            .in0(N__38906),
            .in1(N__38112),
            .in2(_gnd_net_),
            .in3(N__38093),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__46018),
            .ce(N__38750),
            .sr(N__45594));
    defparam \current_shift_inst.timer_s1.counter_4_LC_16_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_16_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_16_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_16_22_4  (
            .in0(N__38911),
            .in1(N__38088),
            .in2(_gnd_net_),
            .in3(N__38072),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__46018),
            .ce(N__38750),
            .sr(N__45594));
    defparam \current_shift_inst.timer_s1.counter_5_LC_16_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_16_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_16_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_16_22_5  (
            .in0(N__38907),
            .in1(N__38064),
            .in2(_gnd_net_),
            .in3(N__38045),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__46018),
            .ce(N__38750),
            .sr(N__45594));
    defparam \current_shift_inst.timer_s1.counter_6_LC_16_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_16_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_16_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_16_22_6  (
            .in0(N__38912),
            .in1(N__38034),
            .in2(_gnd_net_),
            .in3(N__38018),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__46018),
            .ce(N__38750),
            .sr(N__45594));
    defparam \current_shift_inst.timer_s1.counter_7_LC_16_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_16_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_16_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_16_22_7  (
            .in0(N__38908),
            .in1(N__38013),
            .in2(_gnd_net_),
            .in3(N__37997),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__46018),
            .ce(N__38750),
            .sr(N__45594));
    defparam \current_shift_inst.timer_s1.counter_8_LC_16_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_16_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_16_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_16_23_0  (
            .in0(N__38900),
            .in1(N__37989),
            .in2(_gnd_net_),
            .in3(N__37970),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_16_23_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__46015),
            .ce(N__38767),
            .sr(N__45601));
    defparam \current_shift_inst.timer_s1.counter_9_LC_16_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_16_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_16_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_16_23_1  (
            .in0(N__38904),
            .in1(N__37959),
            .in2(_gnd_net_),
            .in3(N__37940),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__46015),
            .ce(N__38767),
            .sr(N__45601));
    defparam \current_shift_inst.timer_s1.counter_10_LC_16_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_16_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_16_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_16_23_2  (
            .in0(N__38897),
            .in1(N__37935),
            .in2(_gnd_net_),
            .in3(N__37919),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__46015),
            .ce(N__38767),
            .sr(N__45601));
    defparam \current_shift_inst.timer_s1.counter_11_LC_16_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_16_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_16_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_16_23_3  (
            .in0(N__38901),
            .in1(N__38346),
            .in2(_gnd_net_),
            .in3(N__38327),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__46015),
            .ce(N__38767),
            .sr(N__45601));
    defparam \current_shift_inst.timer_s1.counter_12_LC_16_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_16_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_16_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_16_23_4  (
            .in0(N__38898),
            .in1(N__38319),
            .in2(_gnd_net_),
            .in3(N__38300),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__46015),
            .ce(N__38767),
            .sr(N__45601));
    defparam \current_shift_inst.timer_s1.counter_13_LC_16_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_16_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_16_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_16_23_5  (
            .in0(N__38902),
            .in1(N__38292),
            .in2(_gnd_net_),
            .in3(N__38273),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__46015),
            .ce(N__38767),
            .sr(N__45601));
    defparam \current_shift_inst.timer_s1.counter_14_LC_16_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_16_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_16_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_16_23_6  (
            .in0(N__38899),
            .in1(N__38262),
            .in2(_gnd_net_),
            .in3(N__38246),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__46015),
            .ce(N__38767),
            .sr(N__45601));
    defparam \current_shift_inst.timer_s1.counter_15_LC_16_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_16_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_16_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_16_23_7  (
            .in0(N__38903),
            .in1(N__38241),
            .in2(_gnd_net_),
            .in3(N__38225),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__46015),
            .ce(N__38767),
            .sr(N__45601));
    defparam \current_shift_inst.timer_s1.counter_16_LC_16_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_16_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_16_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_16_24_0  (
            .in0(N__38869),
            .in1(N__38217),
            .in2(_gnd_net_),
            .in3(N__38198),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_16_24_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__46012),
            .ce(N__38768),
            .sr(N__45608));
    defparam \current_shift_inst.timer_s1.counter_17_LC_16_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_16_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_16_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_16_24_1  (
            .in0(N__38873),
            .in1(N__38184),
            .in2(_gnd_net_),
            .in3(N__38165),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__46012),
            .ce(N__38768),
            .sr(N__45608));
    defparam \current_shift_inst.timer_s1.counter_18_LC_16_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_16_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_16_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_16_24_2  (
            .in0(N__38870),
            .in1(N__38160),
            .in2(_gnd_net_),
            .in3(N__38144),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__46012),
            .ce(N__38768),
            .sr(N__45608));
    defparam \current_shift_inst.timer_s1.counter_19_LC_16_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_16_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_16_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_16_24_3  (
            .in0(N__38874),
            .in1(N__38136),
            .in2(_gnd_net_),
            .in3(N__38561),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__46012),
            .ce(N__38768),
            .sr(N__45608));
    defparam \current_shift_inst.timer_s1.counter_20_LC_16_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_16_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_16_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_16_24_4  (
            .in0(N__38871),
            .in1(N__38553),
            .in2(_gnd_net_),
            .in3(N__38534),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__46012),
            .ce(N__38768),
            .sr(N__45608));
    defparam \current_shift_inst.timer_s1.counter_21_LC_16_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_16_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_16_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_16_24_5  (
            .in0(N__38875),
            .in1(N__38526),
            .in2(_gnd_net_),
            .in3(N__38507),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__46012),
            .ce(N__38768),
            .sr(N__45608));
    defparam \current_shift_inst.timer_s1.counter_22_LC_16_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_16_24_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_16_24_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_16_24_6  (
            .in0(N__38872),
            .in1(N__38496),
            .in2(_gnd_net_),
            .in3(N__38480),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__46012),
            .ce(N__38768),
            .sr(N__45608));
    defparam \current_shift_inst.timer_s1.counter_23_LC_16_24_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_16_24_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_16_24_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_16_24_7  (
            .in0(N__38876),
            .in1(N__38475),
            .in2(_gnd_net_),
            .in3(N__38459),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__46012),
            .ce(N__38768),
            .sr(N__45608));
    defparam \current_shift_inst.timer_s1.counter_24_LC_16_25_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_16_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_16_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_16_25_0  (
            .in0(N__38865),
            .in1(N__38451),
            .in2(_gnd_net_),
            .in3(N__38432),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_16_25_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__46006),
            .ce(N__38766),
            .sr(N__45622));
    defparam \current_shift_inst.timer_s1.counter_25_LC_16_25_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_16_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_16_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_16_25_1  (
            .in0(N__38877),
            .in1(N__38421),
            .in2(_gnd_net_),
            .in3(N__38402),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__46006),
            .ce(N__38766),
            .sr(N__45622));
    defparam \current_shift_inst.timer_s1.counter_26_LC_16_25_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_16_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_16_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_16_25_2  (
            .in0(N__38866),
            .in1(N__38397),
            .in2(_gnd_net_),
            .in3(N__38381),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__46006),
            .ce(N__38766),
            .sr(N__45622));
    defparam \current_shift_inst.timer_s1.counter_27_LC_16_25_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_16_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_16_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_16_25_3  (
            .in0(N__38878),
            .in1(N__38373),
            .in2(_gnd_net_),
            .in3(N__38354),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__46006),
            .ce(N__38766),
            .sr(N__45622));
    defparam \current_shift_inst.timer_s1.counter_28_LC_16_25_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_16_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_16_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_16_25_4  (
            .in0(N__38867),
            .in1(N__38929),
            .in2(_gnd_net_),
            .in3(N__38915),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__46006),
            .ce(N__38766),
            .sr(N__45622));
    defparam \current_shift_inst.timer_s1.counter_29_LC_16_25_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_16_25_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_16_25_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_16_25_5  (
            .in0(N__38782),
            .in1(N__38868),
            .in2(_gnd_net_),
            .in3(N__38786),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46006),
            .ce(N__38766),
            .sr(N__45622));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_17_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_17_6_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_17_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_17_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38725),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46108),
            .ce(N__38695),
            .sr(N__45515));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_17_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_17_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_17_7_0  (
            .in0(N__38670),
            .in1(N__38619),
            .in2(N__38653),
            .in3(N__38635),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_17_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_17_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_17_7_1 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKL65B1_3_LC_17_7_1  (
            .in0(N__38590),
            .in1(N__43141),
            .in2(N__38624),
            .in3(N__39109),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_17_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_17_7_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRHL2M1_3_LC_17_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38606),
            .in3(N__42695),
            .lcout(elapsed_time_ns_1_RNIRHL2M1_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_17_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_17_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_17_7_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_16_LC_17_7_3  (
            .in0(N__42670),
            .in1(N__42614),
            .in2(N__42647),
            .in3(N__42632),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_381 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_381_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_17_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_17_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_17_7_4 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_17_7_4  (
            .in0(N__43427),
            .in1(N__43378),
            .in2(N__38564),
            .in3(N__42581),
            .lcout(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ),
            .ltout(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_17_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_17_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_17_7_5 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_17_7_5  (
            .in0(N__39398),
            .in1(N__39308),
            .in2(N__39152),
            .in3(N__42962),
            .lcout(elapsed_time_ns_1_RNIRAIF91_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_17_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_17_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_17_7_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILL1NA_6_LC_17_7_6  (
            .in0(N__45716),
            .in1(N__43377),
            .in2(_gnd_net_),
            .in3(N__42580),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_17_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_17_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_17_7_7 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAKOL_31_LC_17_7_7  (
            .in0(N__43428),
            .in1(N__45717),
            .in2(N__39149),
            .in3(N__39146),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_17_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_17_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_17_8_0  (
            .in0(N__38992),
            .in1(N__39317),
            .in2(N__39040),
            .in3(N__42810),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_17_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_17_8_1 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_17_8_1  (
            .in0(N__39064),
            .in1(N__39033),
            .in2(N__42596),
            .in3(N__38991),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_348_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_17_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_17_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_17_8_2 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_17_8_2  (
            .in0(_gnd_net_),
            .in1(N__39316),
            .in2(N__39020),
            .in3(N__39013),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_17_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_17_8_3 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_17_8_3  (
            .in0(N__43099),
            .in1(N__39331),
            .in2(N__39231),
            .in3(N__42957),
            .lcout(elapsed_time_ns_1_RNIR9HF91_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_17_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_17_8_4 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_17_8_4  (
            .in0(N__38993),
            .in1(N__43101),
            .in2(N__42983),
            .in3(N__38981),
            .lcout(elapsed_time_ns_1_RNIFJ2591_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_17_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_17_8_5 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_17_8_5  (
            .in0(N__43100),
            .in1(N__38939),
            .in2(N__39293),
            .in3(N__42958),
            .lcout(elapsed_time_ns_1_RNITCIF91_0_23),
            .ltout(elapsed_time_ns_1_RNITCIF91_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_17_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_17_8_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_17_8_6  (
            .in0(N__42529),
            .in1(N__43240),
            .in2(N__39401),
            .in3(N__39397),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_17_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_17_8_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_17_8_7  (
            .in0(N__43204),
            .in1(N__43463),
            .in2(N__39386),
            .in3(N__40091),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_17_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_17_9_0 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_17_9_0  (
            .in0(N__43107),
            .in1(N__39383),
            .in2(N__39363),
            .in3(N__42951),
            .lcout(elapsed_time_ns_1_RNIDH2591_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_17_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_17_9_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_17_9_1  (
            .in0(N__39274),
            .in1(N__43351),
            .in2(N__39332),
            .in3(N__40039),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_347 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_17_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_17_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_17_9_2  (
            .in0(N__39169),
            .in1(N__43453),
            .in2(N__43306),
            .in3(N__43189),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_9_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_9_3  (
            .in0(N__42544),
            .in1(N__39304),
            .in2(N__43267),
            .in3(N__39286),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_17_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_17_9_4 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_17_9_4  (
            .in0(N__43103),
            .in1(N__39252),
            .in2(N__42975),
            .in3(N__39275),
            .lcout(elapsed_time_ns_1_RNIQ8HF91_0_11),
            .ltout(elapsed_time_ns_1_RNIQ8HF91_0_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_17_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_17_9_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_17_9_5  (
            .in0(N__40017),
            .in1(N__43323),
            .in2(N__39239),
            .in3(N__39216),
            .lcout(\phase_controller_inst1.stoper_tr.N_244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_17_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_17_9_6 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_17_9_6  (
            .in0(N__39170),
            .in1(N__42950),
            .in2(N__43145),
            .in3(N__39158),
            .lcout(elapsed_time_ns_1_RNI3JIF91_0_29),
            .ltout(elapsed_time_ns_1_RNI3JIF91_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_17_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_17_9_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_17_9_7  (
            .in0(N__42853),
            .in1(_gnd_net_),
            .in2(N__40094),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_17_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_17_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_17_10_0 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_17_10_0  (
            .in0(N__39998),
            .in1(N__39899),
            .in2(N__40085),
            .in3(N__39716),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46087),
            .ce(N__39597),
            .sr(N__45534));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_17_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_17_10_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_17_10_3  (
            .in0(N__43137),
            .in1(N__40040),
            .in2(N__42992),
            .in3(N__40024),
            .lcout(elapsed_time_ns_1_RNISAHF91_0_13),
            .ltout(elapsed_time_ns_1_RNISAHF91_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_17_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_17_10_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_17_10_4  (
            .in0(N__39997),
            .in1(N__39898),
            .in2(N__39941),
            .in3(N__39715),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46087),
            .ce(N__39597),
            .sr(N__45534));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_17_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_17_10_6 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_17_10_6  (
            .in0(N__39926),
            .in1(N__39897),
            .in2(_gnd_net_),
            .in3(N__39714),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46087),
            .ce(N__39597),
            .sr(N__45534));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_1_c_inv_LC_17_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_1_c_inv_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_1_c_inv_LC_17_11_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_1_c_inv_LC_17_11_0  (
            .in0(N__44122),
            .in1(N__39467),
            .in2(N__39455),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_2_c_inv_LC_17_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_2_c_inv_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_2_c_inv_LC_17_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_2_c_inv_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__39443),
            .in2(N__39431),
            .in3(N__40490),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_3_c_inv_LC_17_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_3_c_inv_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_3_c_inv_LC_17_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_3_c_inv_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__39422),
            .in2(N__39410),
            .in3(N__40472),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_4_c_inv_LC_17_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_4_c_inv_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_4_c_inv_LC_17_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_4_c_inv_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(N__40265),
            .in2(N__40253),
            .in3(N__40454),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_5_c_inv_LC_17_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_5_c_inv_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_5_c_inv_LC_17_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_5_c_inv_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(N__40244),
            .in2(N__40232),
            .in3(N__40745),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_6_c_inv_LC_17_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_6_c_inv_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_6_c_inv_LC_17_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_6_c_inv_LC_17_11_5  (
            .in0(N__40727),
            .in1(N__40223),
            .in2(N__40211),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_7_c_inv_LC_17_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_7_c_inv_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_7_c_inv_LC_17_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_7_c_inv_LC_17_11_6  (
            .in0(_gnd_net_),
            .in1(N__40202),
            .in2(N__40190),
            .in3(N__40709),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_8_c_inv_LC_17_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_8_c_inv_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_8_c_inv_LC_17_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_8_c_inv_LC_17_11_7  (
            .in0(_gnd_net_),
            .in1(N__40181),
            .in2(N__40169),
            .in3(N__40691),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_9_c_inv_LC_17_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_9_c_inv_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_9_c_inv_LC_17_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_9_c_inv_LC_17_12_0  (
            .in0(_gnd_net_),
            .in1(N__40157),
            .in2(N__40145),
            .in3(N__40673),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_10_c_inv_LC_17_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_10_c_inv_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_10_c_inv_LC_17_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_10_c_inv_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__40136),
            .in2(N__40124),
            .in3(N__40655),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_11_c_inv_LC_17_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_11_c_inv_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_11_c_inv_LC_17_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_11_c_inv_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(N__40115),
            .in2(N__40103),
            .in3(N__40637),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_12_c_inv_LC_17_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_12_c_inv_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_12_c_inv_LC_17_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_12_c_inv_LC_17_12_3  (
            .in0(_gnd_net_),
            .in1(N__40436),
            .in2(N__40424),
            .in3(N__40619),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_13_c_inv_LC_17_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_13_c_inv_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_13_c_inv_LC_17_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_13_c_inv_LC_17_12_4  (
            .in0(_gnd_net_),
            .in1(N__40415),
            .in2(N__40403),
            .in3(N__40601),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_14_c_inv_LC_17_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_14_c_inv_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_14_c_inv_LC_17_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_14_c_inv_LC_17_12_5  (
            .in0(N__40868),
            .in1(N__40394),
            .in2(N__40382),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_15_c_inv_LC_17_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_15_c_inv_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_15_c_inv_LC_17_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_15_c_inv_LC_17_12_6  (
            .in0(_gnd_net_),
            .in1(N__40370),
            .in2(N__40358),
            .in3(N__40850),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_16_c_inv_LC_17_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_16_c_inv_LC_17_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_16_c_inv_LC_17_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_16_c_inv_LC_17_12_7  (
            .in0(_gnd_net_),
            .in1(N__40349),
            .in2(N__40337),
            .in3(N__40829),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_17_c_inv_LC_17_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_17_c_inv_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_17_c_inv_LC_17_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_17_c_inv_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(N__40328),
            .in2(N__40316),
            .in3(N__40811),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_18_c_inv_LC_17_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_18_c_inv_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_18_c_inv_LC_17_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_18_c_inv_LC_17_13_1  (
            .in0(_gnd_net_),
            .in1(N__40307),
            .in2(N__40295),
            .in3(N__40793),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_inv_LC_17_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_inv_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_inv_LC_17_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_inv_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(N__40286),
            .in2(N__40274),
            .in3(N__40772),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_17_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_17_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_LUT4_0_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40583),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_17_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_17_13_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_17_13_5  (
            .in0(N__43496),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44139),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNILGTP_LC_17_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNILGTP_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNILGTP_LC_17_13_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNILGTP_LC_17_13_6  (
            .in0(_gnd_net_),
            .in1(N__43565),
            .in2(_gnd_net_),
            .in3(N__43608),
            .lcout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_17_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_17_13_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a3_1_LC_17_13_7  (
            .in0(_gnd_net_),
            .in1(N__40551),
            .in2(_gnd_net_),
            .in3(N__43664),
            .lcout(state_ns_i_a3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(N__40496),
            .in2(N__44123),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_17_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_17_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_17_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_17_14_1  (
            .in0(N__44256),
            .in1(N__40489),
            .in2(_gnd_net_),
            .in3(N__40475),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__46061),
            .ce(),
            .sr(N__45552));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_17_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_17_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_17_14_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_17_14_2  (
            .in0(N__44271),
            .in1(N__40471),
            .in2(N__43592),
            .in3(N__40457),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__46061),
            .ce(),
            .sr(N__45552));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_17_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_17_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_17_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_17_14_3  (
            .in0(N__44257),
            .in1(N__40453),
            .in2(_gnd_net_),
            .in3(N__40439),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__46061),
            .ce(),
            .sr(N__45552));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_17_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_17_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_17_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_17_14_4  (
            .in0(N__44272),
            .in1(N__40744),
            .in2(_gnd_net_),
            .in3(N__40730),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__46061),
            .ce(),
            .sr(N__45552));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_17_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_17_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_17_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_17_14_5  (
            .in0(N__44258),
            .in1(N__40726),
            .in2(_gnd_net_),
            .in3(N__40712),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__46061),
            .ce(),
            .sr(N__45552));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_17_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_17_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_17_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_17_14_6  (
            .in0(N__44273),
            .in1(N__40708),
            .in2(_gnd_net_),
            .in3(N__40694),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__46061),
            .ce(),
            .sr(N__45552));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_17_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_17_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_17_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_17_14_7  (
            .in0(N__44259),
            .in1(N__40690),
            .in2(_gnd_net_),
            .in3(N__40676),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__46061),
            .ce(),
            .sr(N__45552));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_17_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_17_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_17_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_17_15_0  (
            .in0(N__44267),
            .in1(N__40672),
            .in2(_gnd_net_),
            .in3(N__40658),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__46053),
            .ce(),
            .sr(N__45556));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_17_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_17_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_17_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_17_15_1  (
            .in0(N__44260),
            .in1(N__40654),
            .in2(_gnd_net_),
            .in3(N__40640),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__46053),
            .ce(),
            .sr(N__45556));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_17_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_17_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_17_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_17_15_2  (
            .in0(N__44264),
            .in1(N__40636),
            .in2(_gnd_net_),
            .in3(N__40622),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__46053),
            .ce(),
            .sr(N__45556));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_17_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_17_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_17_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_17_15_3  (
            .in0(N__44261),
            .in1(N__40618),
            .in2(_gnd_net_),
            .in3(N__40604),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__46053),
            .ce(),
            .sr(N__45556));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_17_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_17_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_17_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_17_15_4  (
            .in0(N__44265),
            .in1(N__40600),
            .in2(_gnd_net_),
            .in3(N__40586),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__46053),
            .ce(),
            .sr(N__45556));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_17_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_17_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_17_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_17_15_5  (
            .in0(N__44262),
            .in1(N__40867),
            .in2(_gnd_net_),
            .in3(N__40853),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__46053),
            .ce(),
            .sr(N__45556));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_17_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_17_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_17_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_17_15_6  (
            .in0(N__44266),
            .in1(N__40846),
            .in2(_gnd_net_),
            .in3(N__40832),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__46053),
            .ce(),
            .sr(N__45556));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_17_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_17_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_17_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_17_15_7  (
            .in0(N__44263),
            .in1(N__40828),
            .in2(_gnd_net_),
            .in3(N__40814),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__46053),
            .ce(),
            .sr(N__45556));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_17_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_17_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_17_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_17_16_0  (
            .in0(N__44268),
            .in1(N__40810),
            .in2(_gnd_net_),
            .in3(N__40796),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__46047),
            .ce(),
            .sr(N__45560));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_17_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_17_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_17_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_17_16_1  (
            .in0(N__44270),
            .in1(N__40792),
            .in2(_gnd_net_),
            .in3(N__40778),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__46047),
            .ce(),
            .sr(N__45560));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_17_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_17_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_17_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_17_16_2  (
            .in0(N__44269),
            .in1(N__40771),
            .in2(_gnd_net_),
            .in3(N__40775),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46047),
            .ce(),
            .sr(N__45560));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_17_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_17_17_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_17_17_0  (
            .in0(N__47344),
            .in1(N__41197),
            .in2(N__46980),
            .in3(N__41167),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_17_1 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_17_1  (
            .in0(N__41198),
            .in1(N__47345),
            .in2(N__41171),
            .in3(N__46922),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_17_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_17_2  (
            .in0(N__47341),
            .in1(N__41196),
            .in2(_gnd_net_),
            .in3(N__41166),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_1_11_LC_17_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_1_11_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_1_11_LC_17_17_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_RNO_1_11_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__47346),
            .in2(_gnd_net_),
            .in3(N__46918),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_17_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_17_4  (
            .in0(N__47342),
            .in1(N__41116),
            .in2(N__46981),
            .in3(N__41086),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_17_5 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_17_5  (
            .in0(N__41117),
            .in1(N__47343),
            .in2(N__41090),
            .in3(N__46926),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_17_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_17_6  (
            .in0(N__42190),
            .in1(N__41115),
            .in2(_gnd_net_),
            .in3(N__41085),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41052),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46041),
            .ce(N__41023),
            .sr(N__45564));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_17_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_17_18_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_17_18_0  (
            .in0(N__44591),
            .in1(N__40991),
            .in2(_gnd_net_),
            .in3(N__40925),
            .lcout(\current_shift_inst.control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_17_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_17_18_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_17_18_1  (
            .in0(N__40926),
            .in1(N__44558),
            .in2(_gnd_net_),
            .in3(N__40970),
            .lcout(\current_shift_inst.control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_17_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_17_18_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_17_18_2  (
            .in0(N__40949),
            .in1(N__44549),
            .in2(_gnd_net_),
            .in3(N__40927),
            .lcout(\current_shift_inst.control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_17_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_17_18_4 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_17_18_4  (
            .in0(N__47339),
            .in1(N__41786),
            .in2(N__41750),
            .in3(N__46972),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_17_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_17_18_5 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI81DJ11_2_LC_17_18_5  (
            .in0(N__41717),
            .in1(N__41609),
            .in2(N__41579),
            .in3(N__41373),
            .lcout(elapsed_time_ns_1_RNI81DJ11_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_18_6 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_18_6  (
            .in0(N__47338),
            .in1(N__46971),
            .in2(N__42446),
            .in3(N__42488),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_18_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_18_7  (
            .in0(N__46970),
            .in1(N__47340),
            .in2(N__41354),
            .in3(N__41303),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_17_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_17_19_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_17_19_0  (
            .in0(N__46984),
            .in1(N__47354),
            .in2(N__42122),
            .in3(N__42083),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_19_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_19_1  (
            .in0(N__42218),
            .in1(N__41226),
            .in2(_gnd_net_),
            .in3(N__41253),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_19_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_19_2  (
            .in0(N__44775),
            .in1(N__42219),
            .in2(_gnd_net_),
            .in3(N__44734),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_17_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_17_19_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_17_19_3  (
            .in0(N__47355),
            .in1(N__46983),
            .in2(N__41260),
            .in3(N__41227),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_17_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_17_19_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_17_19_6  (
            .in0(N__46982),
            .in1(N__47356),
            .in2(N__42340),
            .in3(N__42291),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_20_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_20_2  (
            .in0(N__42217),
            .in1(N__42486),
            .in2(_gnd_net_),
            .in3(N__42441),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_17_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_17_20_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_17_20_3  (
            .in0(N__42386),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_20_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_20_5  (
            .in0(N__42220),
            .in1(N__42330),
            .in2(_gnd_net_),
            .in3(N__42293),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_20_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_20_6  (
            .in0(N__42216),
            .in1(N__42111),
            .in2(_gnd_net_),
            .in3(N__42082),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_17_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_17_20_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_17_20_7  (
            .in0(N__47353),
            .in1(N__42043),
            .in2(N__47005),
            .in3(N__42014),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.T01_LC_17_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.T01_LC_17_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T01_LC_17_21_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst2.T01_LC_17_21_1  (
            .in0(N__41899),
            .in1(N__41986),
            .in2(_gnd_net_),
            .in3(N__41857),
            .lcout(T01_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46026),
            .ce(),
            .sr(N__45583));
    defparam \phase_controller_inst2.state_1_LC_17_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_17_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_17_23_5 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst2.state_1_LC_17_23_5  (
            .in0(N__43748),
            .in1(N__41887),
            .in2(N__46221),
            .in3(N__41846),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46019),
            .ce(),
            .sr(N__45595));
    defparam \phase_controller_inst2.T12_LC_17_25_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.T12_LC_17_25_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T12_LC_17_25_1 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_inst2.T12_LC_17_25_1  (
            .in0(N__41797),
            .in1(N__46229),
            .in2(_gnd_net_),
            .in3(N__41858),
            .lcout(T12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46013),
            .ce(),
            .sr(N__45609));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_18_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_18_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_18_7_0 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_18_7_0  (
            .in0(N__42838),
            .in1(N__42823),
            .in2(N__42794),
            .in3(N__42755),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_363_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_18_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_18_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_18_7_1 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_18_7_1  (
            .in0(N__43426),
            .in1(N__42631),
            .in2(N__42749),
            .in3(N__42643),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_18_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_18_7_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_16_LC_18_7_2  (
            .in0(N__45714),
            .in1(N__42674),
            .in2(N__42659),
            .in3(N__42613),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_18_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_18_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_18_7_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIME943_20_LC_18_7_3  (
            .in0(N__42517),
            .in1(N__43228),
            .in2(N__42571),
            .in3(N__42656),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_18_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_18_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_18_7_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI56UV7_1_LC_18_7_4  (
            .in0(N__42630),
            .in1(N__42612),
            .in2(N__42599),
            .in3(N__42595),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_359_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_18_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_18_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_18_7_5 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_18_7_5  (
            .in0(N__43475),
            .in1(N__42956),
            .in2(N__42572),
            .in3(N__43140),
            .lcout(elapsed_time_ns_1_RNI0GIF91_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_18_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_18_8_0 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_18_8_0  (
            .in0(N__42942),
            .in1(N__42551),
            .in2(N__42533),
            .in3(N__43073),
            .lcout(elapsed_time_ns_1_RNIUDIF91_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_18_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_18_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_18_8_1 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_18_8_1  (
            .in0(N__42518),
            .in1(N__42494),
            .in2(N__43121),
            .in3(N__42940),
            .lcout(elapsed_time_ns_1_RNIVEIF91_0_25),
            .ltout(elapsed_time_ns_1_RNIVEIF91_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_18_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_18_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_18_8_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_18_8_2  (
            .in0(N__43438),
            .in1(N__43279),
            .in2(N__43478),
            .in3(N__43474),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_18_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_18_8_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_18_8_3  (
            .in0(N__43069),
            .in1(N__43457),
            .in2(N__42991),
            .in3(N__43439),
            .lcout(elapsed_time_ns_1_RNI2IIF91_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_18_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_18_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_18_8_4 .LUT_INIT=16'b1111111111001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_18_8_4  (
            .in0(N__43429),
            .in1(N__45715),
            .in2(N__43385),
            .in3(N__43361),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_18_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_18_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_18_8_5 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_18_8_5  (
            .in0(N__43070),
            .in1(N__43355),
            .in2(N__43340),
            .in3(N__43329),
            .lcout(elapsed_time_ns_1_RNIP7HF91_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_18_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_18_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_18_8_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_18_8_6  (
            .in0(N__42941),
            .in1(N__43071),
            .in2(N__43286),
            .in3(N__43307),
            .lcout(elapsed_time_ns_1_RNI1HIF91_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_18_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_18_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_18_8_7 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_18_8_7  (
            .in0(N__43072),
            .in1(N__43268),
            .in2(N__43244),
            .in3(N__42943),
            .lcout(elapsed_time_ns_1_RNISBIF91_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_18_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_18_9_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_18_9_0  (
            .in0(N__43139),
            .in1(N__43229),
            .in2(N__42982),
            .in3(N__43205),
            .lcout(elapsed_time_ns_1_RNIQ9IF91_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_18_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_18_9_1 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_18_9_1  (
            .in0(N__43193),
            .in1(N__43138),
            .in2(N__42857),
            .in3(N__42952),
            .lcout(elapsed_time_ns_1_RNIRBJF91_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_18_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_18_9_7 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_18_9_7  (
            .in0(N__43825),
            .in1(N__43763),
            .in2(_gnd_net_),
            .in3(N__43933),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_18_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_18_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_18_10_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_18_10_1  (
            .in0(_gnd_net_),
            .in1(N__43934),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46094),
            .ce(),
            .sr(N__45530));
    defparam \phase_controller_inst1.stoper_hc.running_LC_18_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_18_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_18_11_3 .LUT_INIT=16'b1010111000101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_18_11_3  (
            .in0(N__43762),
            .in1(N__43877),
            .in2(N__43835),
            .in3(N__43793),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46088),
            .ce(),
            .sr(N__45535));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_18_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_18_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_18_12_4  (
            .in0(_gnd_net_),
            .in1(N__46233),
            .in2(_gnd_net_),
            .in3(N__43741),
            .lcout(\phase_controller_inst2.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_LC_18_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_18_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_18_13_0 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_18_13_0  (
            .in0(N__43700),
            .in1(N__43694),
            .in2(N__43679),
            .in3(N__43524),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46073),
            .ce(),
            .sr(N__45544));
    defparam \phase_controller_inst2.stoper_tr.running_LC_18_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_18_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_18_13_2 .LUT_INIT=16'b1100111001001110;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_18_13_2  (
            .in0(N__43498),
            .in1(N__43538),
            .in2(N__43572),
            .in3(N__43612),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46073),
            .ce(),
            .sr(N__45544));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_18_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_18_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_18_13_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_18_13_3  (
            .in0(N__43525),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46073),
            .ce(),
            .sr(N__45544));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIUMLH1_LC_18_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIUMLH1_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIUMLH1_LC_18_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIUMLH1_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(N__43497),
            .in2(_gnd_net_),
            .in3(N__44140),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_19_c_RNIUMLHZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_18_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_18_13_6 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_18_13_6  (
            .in0(N__43561),
            .in1(N__43537),
            .in2(_gnd_net_),
            .in3(N__43523),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(\phase_controller_inst2.stoper_tr.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_18_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_18_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_18_13_7 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_18_13_7  (
            .in0(N__44243),
            .in1(N__44141),
            .in2(N__44126),
            .in3(N__44121),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46073),
            .ce(),
            .sr(N__45544));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_18_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_18_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(N__44099),
            .in2(N__44077),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_18_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_18_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(N__44044),
            .in2(N__44021),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_18_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_18_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(N__46651),
            .in2(N__44003),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_18_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_18_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__43988),
            .in2(N__46824),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_18_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_18_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(N__46655),
            .in2(N__43976),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_18_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_18_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(N__43961),
            .in2(N__46825),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_18_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_18_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__46659),
            .in2(N__43946),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_18_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_18_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(N__44384),
            .in2(N__46826),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_18_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_18_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__46827),
            .in2(N__44375),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_18_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_18_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_LC_18_15_1  (
            .in0(_gnd_net_),
            .in1(N__44360),
            .in2(N__46957),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_18_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_18_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(N__46831),
            .in2(N__44348),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_18_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_18_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(N__45089),
            .in2(N__46958),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_18_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_18_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(N__46835),
            .in2(N__44336),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_18_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_18_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(N__45005),
            .in2(N__46959),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_18_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_18_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(N__46839),
            .in2(N__44321),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_18_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_18_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(N__44306),
            .in2(N__46960),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_18_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_18_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(N__46843),
            .in2(N__45167),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_18_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_18_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(N__44486),
            .in2(N__46961),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_18_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_18_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(N__46847),
            .in2(N__44477),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_18_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_18_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(N__47411),
            .in2(N__46962),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_18_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_18_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(N__46851),
            .in2(N__44645),
            .in3(N__44447),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_18_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_18_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(N__44444),
            .in2(N__46963),
            .in3(N__44429),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_18_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_18_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(N__46855),
            .in2(N__44426),
            .in3(N__44402),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_18_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_18_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_18_16_7  (
            .in0(_gnd_net_),
            .in1(N__44714),
            .in2(N__46964),
            .in3(N__44387),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_18_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_18_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__46859),
            .in2(N__44792),
            .in3(N__44618),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_18_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_18_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__44927),
            .in2(N__46965),
            .in3(N__44603),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_18_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_18_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(N__46863),
            .in2(N__44600),
            .in3(N__44585),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_18_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_18_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(N__46364),
            .in2(N__46966),
            .in3(N__44570),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_18_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_18_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__46867),
            .in2(N__44567),
            .in3(N__44552),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_18_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_18_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__44864),
            .in2(N__46967),
            .in3(N__44543),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_18_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_18_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(N__46871),
            .in2(N__44540),
            .in3(N__44504),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_2_11_LC_18_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_2_11_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_2_11_LC_18_17_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.control_input_RNO_2_11_LC_18_17_7  (
            .in0(N__46872),
            .in1(N__47367),
            .in2(_gnd_net_),
            .in3(N__44501),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_18_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_18_18_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_18_18_1  (
            .in0(N__46877),
            .in1(N__47364),
            .in2(N__45238),
            .in3(N__45191),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_18_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_18_18_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_18_18_2  (
            .in0(N__47362),
            .in1(N__46875),
            .in2(N__45155),
            .in3(N__45113),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_18_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_18_18_3 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_18_18_3  (
            .in0(N__46876),
            .in1(N__45079),
            .in2(N__45041),
            .in3(N__47363),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_18_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_18_18_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_18_18_6  (
            .in0(N__47365),
            .in1(N__46874),
            .in2(N__44996),
            .in3(N__44957),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_18_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_18_18_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_18_18_7  (
            .in0(N__46873),
            .in1(N__47366),
            .in2(N__44921),
            .in3(N__44885),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_18_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_18_19_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_18_19_1  (
            .in0(N__46987),
            .in1(N__47360),
            .in2(N__44858),
            .in3(N__44819),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_19_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_19_3  (
            .in0(N__46985),
            .in1(N__47359),
            .in2(N__44780),
            .in3(N__44735),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_18_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_18_19_6 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_18_19_6  (
            .in0(N__47358),
            .in1(N__46986),
            .in2(N__44705),
            .in3(N__44681),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_18_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_18_19_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_18_19_7  (
            .in0(N__46988),
            .in1(N__47357),
            .in2(N__47474),
            .in3(N__47449),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_18_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_18_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47399),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_18_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_18_20_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_18_20_2  (
            .in0(N__47361),
            .in1(N__47047),
            .in2(N__47006),
            .in3(N__46393),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_18_26_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_18_26_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_18_26_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_18_26_1  (
            .in0(N__46273),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46256),
            .ce(),
            .sr(N__45610));
    defparam \delay_measurement_inst.start_timer_tr_LC_18_26_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_18_26_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_18_26_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_18_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46272),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46256),
            .ce(),
            .sr(N__45610));
    defparam \phase_controller_inst2.T23_LC_18_27_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.T23_LC_18_27_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.T23_LC_18_27_5 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst2.T23_LC_18_27_5  (
            .in0(N__46129),
            .in1(N__46228),
            .in2(_gnd_net_),
            .in3(N__46175),
            .lcout(T23_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46007),
            .ce(),
            .sr(N__45623));
endmodule // MAIN
